magic
tech sky130A
magscale 1 2
timestamp 1607540551
<< locali >>
rect 299765 666587 299799 684437
rect 364349 666587 364383 676141
rect 429485 666587 429519 684437
rect 494069 666587 494103 676141
rect 559205 666587 559239 684437
rect 299765 656999 299799 659685
rect 299581 648227 299615 656829
rect 429301 648023 429335 656829
rect 559021 647887 559055 656829
rect 79609 643127 79643 643365
rect 117237 643263 117271 643637
rect 125793 641767 125827 643705
rect 60657 42619 60691 42721
rect 60599 42585 60691 42619
rect 59829 41939 59863 42517
rect 59921 41463 59955 42585
rect 60013 42075 60047 42449
rect 60105 42347 60139 42449
rect 64613 41531 64647 41905
rect 66821 41803 66855 42585
rect 67557 42007 67591 42721
rect 68201 41599 68235 41973
rect 69489 41803 69523 41905
rect 74365 41803 74399 42721
rect 74457 42619 74491 42789
rect 129565 42789 129749 42823
rect 129565 42687 129599 42789
rect 117053 42143 117087 42381
rect 120457 42279 120491 42449
rect 75377 41871 75411 41973
rect 69581 41463 69615 41769
rect 80253 41531 80287 41633
rect 108957 38675 108991 41973
rect 113189 41803 113223 42109
rect 122481 42075 122515 42449
rect 125333 42347 125367 42653
rect 122699 42245 122791 42279
rect 122757 41803 122791 42245
rect 123861 41871 123895 42313
rect 125367 42109 125609 42143
rect 136189 41871 136223 42585
rect 123953 41599 123987 41837
rect 124045 41599 124079 41769
rect 127633 41667 127667 41837
rect 31677 29019 31711 38573
rect 53297 29019 53331 38573
rect 73537 29019 73571 38573
rect 75745 27659 75779 37213
rect 108957 29019 108991 38505
rect 175013 29019 175047 35853
rect 244381 27659 244415 37213
rect 245945 29019 245979 38573
rect 433441 27659 433475 37213
rect 75469 9707 75503 20961
rect 117697 9707 117731 27557
rect 120457 12427 120491 27557
rect 244289 9707 244323 22729
rect 246037 9707 246071 19261
rect 404461 9707 404495 19261
rect 31493 595 31527 9605
rect 40601 3519 40635 3621
rect 56425 595 56459 3621
rect 75193 3587 75227 4097
rect 82553 3587 82587 3825
rect 82461 3315 82495 3553
rect 57621 595 57655 2805
rect 100493 595 100527 9605
rect 108773 595 108807 9605
rect 433441 8415 433475 17901
rect 115949 3723 115983 4369
rect 395905 3383 395939 3961
rect 401425 3383 401459 3961
rect 422861 3179 422895 3893
rect 422953 3791 422987 3893
rect 423045 3791 423079 3961
rect 431693 3791 431727 3893
rect 431233 3383 431267 3757
rect 432429 3315 432463 3961
rect 432613 3179 432647 3893
rect 431785 2703 431819 2941
rect 432705 2907 432739 3145
rect 431877 2873 432739 2907
rect 431877 2839 431911 2873
rect 433533 595 433567 8245
rect 437431 5321 437489 5355
rect 443009 5219 443043 5321
rect 445585 5219 445619 5321
rect 454049 4947 454083 5321
rect 462329 4947 462363 5253
rect 437489 3791 437523 4165
rect 434487 3145 434579 3179
rect 434545 2975 434579 3145
rect 434729 3111 434763 3349
rect 434821 3111 434855 3281
rect 438593 3247 438627 3961
rect 434453 2771 434487 2941
rect 434729 2295 434763 2941
rect 440065 2907 440099 4029
rect 445493 3859 445527 4165
rect 449633 3723 449667 3893
rect 451841 3791 451875 3893
rect 451841 3757 452669 3791
rect 453773 3723 453807 3893
rect 442181 3247 442215 3281
rect 442181 3213 442457 3247
rect 441537 2771 441571 3009
rect 451749 2839 451783 3689
rect 451933 3451 451967 3621
rect 457361 3451 457395 3893
rect 506155 3757 506305 3791
rect 514033 3655 514067 3893
rect 511089 3451 511123 3553
rect 469229 2975 469263 3417
rect 518173 2839 518207 3689
rect 534641 3043 534675 3281
rect 539517 3247 539551 3349
rect 541541 3145 541909 3179
rect 538781 2975 538815 3077
rect 541541 2975 541575 3145
rect 542921 3009 543105 3043
rect 542829 2771 542863 2941
rect 542921 2907 542955 3009
<< viali >>
rect 299765 684437 299799 684471
rect 429485 684437 429519 684471
rect 299765 666553 299799 666587
rect 364349 676141 364383 676175
rect 364349 666553 364383 666587
rect 559205 684437 559239 684471
rect 429485 666553 429519 666587
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 559205 666553 559239 666587
rect 299765 659685 299799 659719
rect 299765 656965 299799 656999
rect 299581 656829 299615 656863
rect 299581 648193 299615 648227
rect 429301 656829 429335 656863
rect 429301 647989 429335 648023
rect 559021 656829 559055 656863
rect 559021 647853 559055 647887
rect 125793 643705 125827 643739
rect 117237 643637 117271 643671
rect 79609 643365 79643 643399
rect 117237 643229 117271 643263
rect 79609 643093 79643 643127
rect 125793 641733 125827 641767
rect 74457 42789 74491 42823
rect 60657 42721 60691 42755
rect 67557 42721 67591 42755
rect 59921 42585 59955 42619
rect 60565 42585 60599 42619
rect 66821 42585 66855 42619
rect 59829 42517 59863 42551
rect 59829 41905 59863 41939
rect 60013 42449 60047 42483
rect 60105 42449 60139 42483
rect 60105 42313 60139 42347
rect 60013 42041 60047 42075
rect 64613 41905 64647 41939
rect 74365 42721 74399 42755
rect 67557 41973 67591 42007
rect 68201 41973 68235 42007
rect 66821 41769 66855 41803
rect 69489 41905 69523 41939
rect 129749 42789 129783 42823
rect 74457 42585 74491 42619
rect 125333 42653 125367 42687
rect 129565 42653 129599 42687
rect 120457 42449 120491 42483
rect 117053 42381 117087 42415
rect 120457 42245 120491 42279
rect 122481 42449 122515 42483
rect 113189 42109 113223 42143
rect 117053 42109 117087 42143
rect 75377 41973 75411 42007
rect 75377 41837 75411 41871
rect 108957 41973 108991 42007
rect 69489 41769 69523 41803
rect 69581 41769 69615 41803
rect 74365 41769 74399 41803
rect 68201 41565 68235 41599
rect 64613 41497 64647 41531
rect 59921 41429 59955 41463
rect 80253 41633 80287 41667
rect 80253 41497 80287 41531
rect 69581 41429 69615 41463
rect 123861 42313 123895 42347
rect 125333 42313 125367 42347
rect 136189 42585 136223 42619
rect 122665 42245 122699 42279
rect 122481 42041 122515 42075
rect 113189 41769 113223 41803
rect 125333 42109 125367 42143
rect 125609 42109 125643 42143
rect 123861 41837 123895 41871
rect 123953 41837 123987 41871
rect 122757 41769 122791 41803
rect 127633 41837 127667 41871
rect 136189 41837 136223 41871
rect 123953 41565 123987 41599
rect 124045 41769 124079 41803
rect 127633 41633 127667 41667
rect 124045 41565 124079 41599
rect 108957 38641 108991 38675
rect 31677 38573 31711 38607
rect 31677 28985 31711 29019
rect 53297 38573 53331 38607
rect 53297 28985 53331 29019
rect 73537 38573 73571 38607
rect 245945 38573 245979 38607
rect 108957 38505 108991 38539
rect 73537 28985 73571 29019
rect 75745 37213 75779 37247
rect 244381 37213 244415 37247
rect 108957 28985 108991 29019
rect 175013 35853 175047 35887
rect 175013 28985 175047 29019
rect 75745 27625 75779 27659
rect 245945 28985 245979 29019
rect 433441 37213 433475 37247
rect 244381 27625 244415 27659
rect 433441 27625 433475 27659
rect 117697 27557 117731 27591
rect 75469 20961 75503 20995
rect 75469 9673 75503 9707
rect 120457 27557 120491 27591
rect 120457 12393 120491 12427
rect 244289 22729 244323 22763
rect 117697 9673 117731 9707
rect 244289 9673 244323 9707
rect 246037 19261 246071 19295
rect 246037 9673 246071 9707
rect 404461 19261 404495 19295
rect 404461 9673 404495 9707
rect 433441 17901 433475 17935
rect 31493 9605 31527 9639
rect 100493 9605 100527 9639
rect 75193 4097 75227 4131
rect 40601 3621 40635 3655
rect 40601 3485 40635 3519
rect 56425 3621 56459 3655
rect 31493 561 31527 595
rect 82553 3825 82587 3859
rect 75193 3553 75227 3587
rect 82461 3553 82495 3587
rect 82553 3553 82587 3587
rect 82461 3281 82495 3315
rect 56425 561 56459 595
rect 57621 2805 57655 2839
rect 57621 561 57655 595
rect 100493 561 100527 595
rect 108773 9605 108807 9639
rect 433441 8381 433475 8415
rect 433533 8245 433567 8279
rect 115949 4369 115983 4403
rect 115949 3689 115983 3723
rect 395905 3961 395939 3995
rect 395905 3349 395939 3383
rect 401425 3961 401459 3995
rect 423045 3961 423079 3995
rect 401425 3349 401459 3383
rect 422861 3893 422895 3927
rect 422953 3893 422987 3927
rect 422953 3757 422987 3791
rect 432429 3961 432463 3995
rect 431693 3893 431727 3927
rect 423045 3757 423079 3791
rect 431233 3757 431267 3791
rect 431693 3757 431727 3791
rect 431233 3349 431267 3383
rect 432429 3281 432463 3315
rect 432613 3893 432647 3927
rect 422861 3145 422895 3179
rect 432613 3145 432647 3179
rect 432705 3145 432739 3179
rect 431785 2941 431819 2975
rect 431877 2805 431911 2839
rect 431785 2669 431819 2703
rect 108773 561 108807 595
rect 437397 5321 437431 5355
rect 437489 5321 437523 5355
rect 443009 5321 443043 5355
rect 443009 5185 443043 5219
rect 445585 5321 445619 5355
rect 445585 5185 445619 5219
rect 454049 5321 454083 5355
rect 454049 4913 454083 4947
rect 462329 5253 462363 5287
rect 462329 4913 462363 4947
rect 437489 4165 437523 4199
rect 445493 4165 445527 4199
rect 440065 4029 440099 4063
rect 437489 3757 437523 3791
rect 438593 3961 438627 3995
rect 434729 3349 434763 3383
rect 434453 3145 434487 3179
rect 434729 3077 434763 3111
rect 434821 3281 434855 3315
rect 438593 3213 438627 3247
rect 434821 3077 434855 3111
rect 434453 2941 434487 2975
rect 434545 2941 434579 2975
rect 434729 2941 434763 2975
rect 434453 2737 434487 2771
rect 445493 3825 445527 3859
rect 449633 3893 449667 3927
rect 451841 3893 451875 3927
rect 453773 3893 453807 3927
rect 452669 3757 452703 3791
rect 449633 3689 449667 3723
rect 451749 3689 451783 3723
rect 453773 3689 453807 3723
rect 457361 3893 457395 3927
rect 442181 3281 442215 3315
rect 442457 3213 442491 3247
rect 440065 2873 440099 2907
rect 441537 3009 441571 3043
rect 451933 3621 451967 3655
rect 451933 3417 451967 3451
rect 514033 3893 514067 3927
rect 506121 3757 506155 3791
rect 506305 3757 506339 3791
rect 514033 3621 514067 3655
rect 518173 3689 518207 3723
rect 511089 3553 511123 3587
rect 457361 3417 457395 3451
rect 469229 3417 469263 3451
rect 511089 3417 511123 3451
rect 469229 2941 469263 2975
rect 451749 2805 451783 2839
rect 539517 3349 539551 3383
rect 534641 3281 534675 3315
rect 539517 3213 539551 3247
rect 541909 3145 541943 3179
rect 534641 3009 534675 3043
rect 538781 3077 538815 3111
rect 538781 2941 538815 2975
rect 543105 3009 543139 3043
rect 541541 2941 541575 2975
rect 542829 2941 542863 2975
rect 518173 2805 518207 2839
rect 441537 2737 441571 2771
rect 542921 2873 542955 2907
rect 542829 2737 542863 2771
rect 434729 2261 434763 2295
rect 433533 561 433567 595
<< metal1 >>
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 318794 700992 318800 701004
rect 154172 700964 318800 700992
rect 154172 700952 154178 700964
rect 318794 700952 318800 700964
rect 318852 700952 318858 701004
rect 137830 700884 137836 700936
rect 137888 700924 137894 700936
rect 314654 700924 314660 700936
rect 137888 700896 314660 700924
rect 137888 700884 137894 700896
rect 314654 700884 314660 700896
rect 314712 700884 314718 700936
rect 252462 700816 252468 700868
rect 252520 700856 252526 700868
rect 462314 700856 462320 700868
rect 252520 700828 462320 700856
rect 252520 700816 252526 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 105446 700748 105452 700800
rect 105504 700788 105510 700800
rect 322934 700788 322940 700800
rect 105504 700760 322940 700788
rect 105504 700748 105510 700760
rect 322934 700748 322940 700760
rect 322992 700748 322998 700800
rect 256602 700680 256608 700732
rect 256660 700720 256666 700732
rect 478506 700720 478512 700732
rect 256660 700692 478512 700720
rect 256660 700680 256666 700692
rect 478506 700680 478512 700692
rect 478564 700680 478570 700732
rect 89162 700612 89168 700664
rect 89220 700652 89226 700664
rect 331214 700652 331220 700664
rect 89220 700624 331220 700652
rect 89220 700612 89226 700624
rect 331214 700612 331220 700624
rect 331272 700612 331278 700664
rect 72970 700544 72976 700596
rect 73028 700584 73034 700596
rect 327074 700584 327080 700596
rect 73028 700556 327080 700584
rect 73028 700544 73034 700556
rect 327074 700544 327080 700556
rect 327132 700544 327138 700596
rect 240042 700476 240048 700528
rect 240100 700516 240106 700528
rect 527174 700516 527180 700528
rect 240100 700488 527180 700516
rect 240100 700476 240106 700488
rect 527174 700476 527180 700488
rect 527232 700476 527238 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 335354 700448 335360 700460
rect 40552 700420 335360 700448
rect 40552 700408 40558 700420
rect 335354 700408 335360 700420
rect 335412 700408 335418 700460
rect 244182 700340 244188 700392
rect 244240 700380 244246 700392
rect 543458 700380 543464 700392
rect 244240 700352 543464 700380
rect 244240 700340 244246 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 343634 700312 343640 700324
rect 24360 700284 343640 700312
rect 24360 700272 24366 700284
rect 343634 700272 343640 700284
rect 343692 700272 343698 700324
rect 269022 700204 269028 700256
rect 269080 700244 269086 700256
rect 413646 700244 413652 700256
rect 269080 700216 413652 700244
rect 269080 700204 269086 700216
rect 413646 700204 413652 700216
rect 413704 700204 413710 700256
rect 170306 700136 170312 700188
rect 170364 700176 170370 700188
rect 310514 700176 310520 700188
rect 170364 700148 310520 700176
rect 170364 700136 170370 700148
rect 310514 700136 310520 700148
rect 310572 700136 310578 700188
rect 264882 700068 264888 700120
rect 264940 700108 264946 700120
rect 397454 700108 397460 700120
rect 264940 700080 397460 700108
rect 264940 700068 264946 700080
rect 397454 700068 397460 700080
rect 397512 700068 397518 700120
rect 202782 700000 202788 700052
rect 202840 700040 202846 700052
rect 302234 700040 302240 700052
rect 202840 700012 302240 700040
rect 202840 700000 202846 700012
rect 302234 700000 302240 700012
rect 302292 700000 302298 700052
rect 218974 699932 218980 699984
rect 219032 699972 219038 699984
rect 306374 699972 306380 699984
rect 219032 699944 306380 699972
rect 219032 699932 219038 699944
rect 306374 699932 306380 699944
rect 306432 699932 306438 699984
rect 281442 699864 281448 699916
rect 281500 699904 281506 699916
rect 348786 699904 348792 699916
rect 281500 699876 348792 699904
rect 281500 699864 281506 699876
rect 348786 699864 348792 699876
rect 348844 699864 348850 699916
rect 277302 699796 277308 699848
rect 277360 699836 277366 699848
rect 332502 699836 332508 699848
rect 277360 699808 332508 699836
rect 277360 699796 277366 699808
rect 332502 699796 332508 699808
rect 332560 699796 332566 699848
rect 267642 699728 267648 699780
rect 267700 699768 267706 699780
rect 288434 699768 288440 699780
rect 267700 699740 288440 699768
rect 267700 699728 267706 699740
rect 288434 699728 288440 699740
rect 288492 699728 288498 699780
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 283834 699660 283840 699712
rect 283892 699700 283898 699712
rect 293954 699700 293960 699712
rect 283892 699672 293960 699700
rect 283892 699660 283898 699672
rect 293954 699660 293960 699672
rect 294012 699660 294018 699712
rect 227622 696940 227628 696992
rect 227680 696980 227686 696992
rect 580166 696980 580172 696992
rect 227680 696952 580172 696980
rect 227680 696940 227686 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 299658 688576 299664 688628
rect 299716 688616 299722 688628
rect 300118 688616 300124 688628
rect 299716 688588 300124 688616
rect 299716 688576 299722 688588
rect 300118 688576 300124 688588
rect 300176 688576 300182 688628
rect 429378 688576 429384 688628
rect 429436 688616 429442 688628
rect 429838 688616 429844 688628
rect 429436 688588 429844 688616
rect 429436 688576 429442 688588
rect 429838 688576 429844 688588
rect 429896 688576 429902 688628
rect 559098 688576 559104 688628
rect 559156 688616 559162 688628
rect 559650 688616 559656 688628
rect 559156 688588 559656 688616
rect 559156 688576 559162 688588
rect 559650 688576 559656 688588
rect 559708 688576 559714 688628
rect 299492 685936 301268 685964
rect 231762 685856 231768 685908
rect 231820 685896 231826 685908
rect 299492 685896 299520 685936
rect 231820 685868 299520 685896
rect 301240 685896 301268 685936
rect 429212 685936 429976 685964
rect 429212 685896 429240 685936
rect 301240 685868 429240 685896
rect 429948 685896 429976 685936
rect 552584 685936 559788 685964
rect 552584 685896 552612 685936
rect 429948 685868 552612 685896
rect 559760 685896 559788 685936
rect 580166 685896 580172 685908
rect 559760 685868 580172 685896
rect 231820 685856 231826 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 299566 684428 299572 684480
rect 299624 684468 299630 684480
rect 299753 684471 299811 684477
rect 299753 684468 299765 684471
rect 299624 684440 299765 684468
rect 299624 684428 299630 684440
rect 299753 684437 299765 684440
rect 299799 684437 299811 684471
rect 299753 684431 299811 684437
rect 429286 684428 429292 684480
rect 429344 684468 429350 684480
rect 429473 684471 429531 684477
rect 429473 684468 429485 684471
rect 429344 684440 429485 684468
rect 429344 684428 429350 684440
rect 429473 684437 429485 684440
rect 429519 684437 429531 684471
rect 429473 684431 429531 684437
rect 559006 684428 559012 684480
rect 559064 684468 559070 684480
rect 559193 684471 559251 684477
rect 559193 684468 559205 684471
rect 559064 684440 559205 684468
rect 559064 684428 559070 684440
rect 559193 684437 559205 684440
rect 559239 684437 559251 684471
rect 559193 684431 559251 684437
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 347774 681748 347780 681760
rect 3568 681720 347780 681748
rect 3568 681708 3574 681720
rect 347774 681708 347780 681720
rect 347832 681708 347838 681760
rect 364334 676172 364340 676184
rect 364295 676144 364340 676172
rect 364334 676132 364340 676144
rect 364392 676132 364398 676184
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 223482 673480 223488 673532
rect 223540 673520 223546 673532
rect 580166 673520 580172 673532
rect 223540 673492 580172 673520
rect 223540 673480 223546 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 356054 667944 356060 667956
rect 3476 667916 356060 667944
rect 3476 667904 3482 667916
rect 356054 667904 356060 667916
rect 356112 667904 356118 667956
rect 299750 666584 299756 666596
rect 299711 666556 299756 666584
rect 299750 666544 299756 666556
rect 299808 666544 299814 666596
rect 364337 666587 364395 666593
rect 364337 666553 364349 666587
rect 364383 666584 364395 666587
rect 364426 666584 364432 666596
rect 364383 666556 364432 666584
rect 364383 666553 364395 666556
rect 364337 666547 364395 666553
rect 364426 666544 364432 666556
rect 364484 666544 364490 666596
rect 429470 666584 429476 666596
rect 429431 666556 429476 666584
rect 429470 666544 429476 666556
rect 429528 666544 429534 666596
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 559190 666584 559196 666596
rect 559151 666556 559196 666584
rect 559190 666544 559196 666556
rect 559248 666544 559254 666596
rect 299750 659716 299756 659728
rect 299711 659688 299756 659716
rect 299750 659676 299756 659688
rect 299808 659676 299814 659728
rect 299658 656956 299664 657008
rect 299716 656996 299722 657008
rect 299753 656999 299811 657005
rect 299753 656996 299765 656999
rect 299716 656968 299765 656996
rect 299716 656956 299722 656968
rect 299753 656965 299765 656968
rect 299799 656965 299811 656999
rect 299753 656959 299811 656965
rect 299566 656860 299572 656872
rect 299527 656832 299572 656860
rect 299566 656820 299572 656832
rect 299624 656820 299630 656872
rect 429286 656860 429292 656872
rect 429247 656832 429292 656860
rect 429286 656820 429292 656832
rect 429344 656820 429350 656872
rect 559006 656860 559012 656872
rect 558967 656832 559012 656860
rect 559006 656820 559012 656832
rect 559064 656820 559070 656872
rect 364334 654100 364340 654152
rect 364392 654140 364398 654152
rect 364518 654140 364524 654152
rect 364392 654112 364524 654140
rect 364392 654100 364398 654112
rect 364518 654100 364524 654112
rect 364576 654100 364582 654152
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 351914 652780 351920 652792
rect 3108 652752 351920 652780
rect 3108 652740 3114 652752
rect 351914 652740 351920 652752
rect 351972 652740 351978 652792
rect 215202 650020 215208 650072
rect 215260 650060 215266 650072
rect 580166 650060 580172 650072
rect 215260 650032 580172 650060
rect 215260 650020 215266 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 285490 648184 285496 648236
rect 285548 648224 285554 648236
rect 299569 648227 299627 648233
rect 299569 648224 299581 648227
rect 285548 648196 299581 648224
rect 285548 648184 285554 648196
rect 299569 648193 299581 648196
rect 299615 648193 299627 648227
rect 299569 648187 299627 648193
rect 235902 648116 235908 648168
rect 235960 648156 235966 648168
rect 298094 648156 298100 648168
rect 235960 648128 298100 648156
rect 235960 648116 235966 648128
rect 298094 648116 298100 648128
rect 298152 648116 298158 648168
rect 272886 648048 272892 648100
rect 272944 648088 272950 648100
rect 364334 648088 364340 648100
rect 272944 648060 364340 648088
rect 272944 648048 272950 648060
rect 364334 648048 364340 648060
rect 364392 648048 364398 648100
rect 260190 647980 260196 648032
rect 260248 648020 260254 648032
rect 429289 648023 429347 648029
rect 429289 648020 429301 648023
rect 260248 647992 429301 648020
rect 260248 647980 260254 647992
rect 429289 647989 429301 647992
rect 429335 647989 429347 648023
rect 429289 647983 429347 647989
rect 247586 647912 247592 647964
rect 247644 647952 247650 647964
rect 494054 647952 494060 647964
rect 247644 647924 494060 647952
rect 247644 647912 247650 647924
rect 494054 647912 494060 647924
rect 494112 647912 494118 647964
rect 234982 647844 234988 647896
rect 235040 647884 235046 647896
rect 559009 647887 559067 647893
rect 559009 647884 559021 647887
rect 235040 647856 559021 647884
rect 235040 647844 235046 647856
rect 559009 647853 559021 647856
rect 559055 647853 559067 647887
rect 559009 647847 559067 647853
rect 180242 647164 180248 647216
rect 180300 647204 180306 647216
rect 386598 647204 386604 647216
rect 180300 647176 386604 647204
rect 180300 647164 180306 647176
rect 386598 647164 386604 647176
rect 386656 647164 386662 647216
rect 125502 647096 125508 647148
rect 125560 647136 125566 647148
rect 168190 647136 168196 647148
rect 125560 647108 168196 647136
rect 125560 647096 125566 647108
rect 168190 647096 168196 647108
rect 168248 647096 168254 647148
rect 191834 647096 191840 647148
rect 191892 647136 191898 647148
rect 407574 647136 407580 647148
rect 191892 647108 407580 647136
rect 191892 647096 191898 647108
rect 407574 647096 407580 647108
rect 407632 647096 407638 647148
rect 167638 647028 167644 647080
rect 167696 647068 167702 647080
rect 522666 647068 522672 647080
rect 167696 647040 522672 647068
rect 167696 647028 167702 647040
rect 522666 647028 522672 647040
rect 522724 647028 522730 647080
rect 3970 646960 3976 647012
rect 4028 647000 4034 647012
rect 365530 647000 365536 647012
rect 4028 646972 365536 647000
rect 4028 646960 4034 646972
rect 365530 646960 365536 646972
rect 365588 646960 365594 647012
rect 150802 646892 150808 646944
rect 150860 646932 150866 646944
rect 525518 646932 525524 646944
rect 150860 646904 525524 646932
rect 150860 646892 150866 646904
rect 525518 646892 525524 646904
rect 525576 646892 525582 646944
rect 5074 646824 5080 646876
rect 5132 646864 5138 646876
rect 382366 646864 382372 646876
rect 5132 646836 382372 646864
rect 5132 646824 5138 646836
rect 382366 646824 382372 646836
rect 382424 646824 382430 646876
rect 154942 646756 154948 646808
rect 155000 646796 155006 646808
rect 537478 646796 537484 646808
rect 155000 646768 537484 646796
rect 155000 646756 155006 646768
rect 537478 646756 537484 646768
rect 537536 646756 537542 646808
rect 104434 646688 104440 646740
rect 104492 646728 104498 646740
rect 140038 646728 140044 646740
rect 104492 646700 140044 646728
rect 104492 646688 104498 646700
rect 140038 646688 140044 646700
rect 140096 646688 140102 646740
rect 142338 646688 142344 646740
rect 142396 646728 142402 646740
rect 525334 646728 525340 646740
rect 142396 646700 525340 646728
rect 142396 646688 142402 646700
rect 525334 646688 525340 646700
rect 525392 646688 525398 646740
rect 138106 646620 138112 646672
rect 138164 646660 138170 646672
rect 525426 646660 525432 646672
rect 138164 646632 525432 646660
rect 138164 646620 138170 646632
rect 525426 646620 525432 646632
rect 525484 646620 525490 646672
rect 129734 646552 129740 646604
rect 129792 646592 129798 646604
rect 525242 646592 525248 646604
rect 129792 646564 525248 646592
rect 129792 646552 129798 646564
rect 525242 646552 525248 646564
rect 525300 646552 525306 646604
rect 3602 646484 3608 646536
rect 3660 646524 3666 646536
rect 432874 646524 432880 646536
rect 3660 646496 432880 646524
rect 3660 646484 3666 646496
rect 432874 646484 432880 646496
rect 432932 646484 432938 646536
rect 4982 646416 4988 646468
rect 5040 646456 5046 646468
rect 441246 646456 441252 646468
rect 5040 646428 441252 646456
rect 5040 646416 5046 646428
rect 441246 646416 441252 646428
rect 441304 646416 441310 646468
rect 6454 646348 6460 646400
rect 6512 646388 6518 646400
rect 445478 646388 445484 646400
rect 6512 646360 445484 646388
rect 6512 646348 6518 646360
rect 445478 646348 445484 646360
rect 445536 646348 445542 646400
rect 6270 646280 6276 646332
rect 6328 646320 6334 646332
rect 458082 646320 458088 646332
rect 6328 646292 458088 646320
rect 6328 646280 6334 646292
rect 458082 646280 458088 646292
rect 458140 646280 458146 646332
rect 4890 646212 4896 646264
rect 4948 646252 4954 646264
rect 466546 646252 466552 646264
rect 4948 646224 466552 646252
rect 4948 646212 4954 646224
rect 466546 646212 466552 646224
rect 466604 646212 466610 646264
rect 6178 646144 6184 646196
rect 6236 646184 6242 646196
rect 470778 646184 470784 646196
rect 6236 646156 470784 646184
rect 6236 646144 6242 646156
rect 470778 646144 470784 646156
rect 470836 646144 470842 646196
rect 10318 646076 10324 646128
rect 10376 646116 10382 646128
rect 483382 646116 483388 646128
rect 10376 646088 483388 646116
rect 10376 646076 10382 646088
rect 483382 646076 483388 646088
rect 483440 646076 483446 646128
rect 13078 646008 13084 646060
rect 13136 646048 13142 646060
rect 495986 646048 495992 646060
rect 13136 646020 495992 646048
rect 13136 646008 13142 646020
rect 495986 646008 495992 646020
rect 496044 646008 496050 646060
rect 4798 645940 4804 645992
rect 4856 645980 4862 645992
rect 491754 645980 491760 645992
rect 4856 645952 491760 645980
rect 4856 645940 4862 645952
rect 491754 645940 491760 645952
rect 491812 645940 491818 645992
rect 14458 645872 14464 645924
rect 14516 645912 14522 645924
rect 508590 645912 508596 645924
rect 14516 645884 508596 645912
rect 14516 645872 14522 645884
rect 508590 645872 508596 645884
rect 508648 645872 508654 645924
rect 25590 645668 25596 645720
rect 25648 645708 25654 645720
rect 378134 645708 378140 645720
rect 25648 645680 378140 645708
rect 25648 645668 25654 645680
rect 378134 645668 378140 645680
rect 378192 645668 378198 645720
rect 159174 645600 159180 645652
rect 159232 645640 159238 645652
rect 525610 645640 525616 645652
rect 159232 645612 525616 645640
rect 159232 645600 159238 645612
rect 525610 645600 525616 645612
rect 525668 645600 525674 645652
rect 40678 645532 40684 645584
rect 40736 645572 40742 645584
rect 416038 645572 416044 645584
rect 40736 645544 416044 645572
rect 40736 645532 40742 645544
rect 416038 645532 416044 645544
rect 416096 645532 416102 645584
rect 7926 645464 7932 645516
rect 7984 645504 7990 645516
rect 386506 645504 386512 645516
rect 7984 645476 386512 645504
rect 7984 645464 7990 645476
rect 386506 645464 386512 645476
rect 386564 645464 386570 645516
rect 386598 645464 386604 645516
rect 386656 645504 386662 645516
rect 580810 645504 580816 645516
rect 386656 645476 580816 645504
rect 386656 645464 386662 645476
rect 580810 645464 580816 645476
rect 580868 645464 580874 645516
rect 133966 645396 133972 645448
rect 134024 645436 134030 645448
rect 524138 645436 524144 645448
rect 134024 645408 524144 645436
rect 134024 645396 134030 645408
rect 524138 645396 524144 645408
rect 524196 645396 524202 645448
rect 7834 645328 7840 645380
rect 7892 645368 7898 645380
rect 399202 645368 399208 645380
rect 7892 645340 399208 645368
rect 7892 645328 7898 645340
rect 399202 645328 399208 645340
rect 399260 645328 399266 645380
rect 7742 645260 7748 645312
rect 7800 645300 7806 645312
rect 411806 645300 411812 645312
rect 7800 645272 411812 645300
rect 7800 645260 7806 645272
rect 411806 645260 411812 645272
rect 411864 645260 411870 645312
rect 168190 645192 168196 645244
rect 168248 645232 168254 645244
rect 580718 645232 580724 645244
rect 168248 645204 580724 645232
rect 168248 645192 168254 645204
rect 580718 645192 580724 645204
rect 580776 645192 580782 645244
rect 7650 645124 7656 645176
rect 7708 645164 7714 645176
rect 424410 645164 424416 645176
rect 7708 645136 424416 645164
rect 7708 645124 7714 645136
rect 424410 645124 424416 645136
rect 424468 645124 424474 645176
rect 108666 645056 108672 645108
rect 108724 645096 108730 645108
rect 523954 645096 523960 645108
rect 108724 645068 523960 645096
rect 108724 645056 108730 645068
rect 523954 645056 523960 645068
rect 524012 645056 524018 645108
rect 9214 644988 9220 645040
rect 9272 645028 9278 645040
rect 437014 645028 437020 645040
rect 9272 645000 437020 645028
rect 9272 644988 9278 645000
rect 437014 644988 437020 645000
rect 437072 644988 437078 645040
rect 83366 644920 83372 644972
rect 83424 644960 83430 644972
rect 522574 644960 522580 644972
rect 83424 644932 522580 644960
rect 83424 644920 83430 644932
rect 522574 644920 522580 644932
rect 522632 644920 522638 644972
rect 6362 644852 6368 644904
rect 6420 644892 6426 644904
rect 449710 644892 449716 644904
rect 6420 644864 449716 644892
rect 6420 644852 6426 644864
rect 449710 644852 449716 644864
rect 449768 644852 449774 644904
rect 70762 644784 70768 644836
rect 70820 644824 70826 644836
rect 522482 644824 522488 644836
rect 70820 644796 522488 644824
rect 70820 644784 70826 644796
rect 522482 644784 522488 644796
rect 522540 644784 522546 644836
rect 7558 644716 7564 644768
rect 7616 644756 7622 644768
rect 462314 644756 462320 644768
rect 7616 644728 462320 644756
rect 7616 644716 7622 644728
rect 462314 644716 462320 644728
rect 462372 644716 462378 644768
rect 9122 644648 9128 644700
rect 9180 644688 9186 644700
rect 474918 644688 474924 644700
rect 9180 644660 474924 644688
rect 9180 644648 9186 644660
rect 474918 644648 474924 644660
rect 474976 644648 474982 644700
rect 9030 644580 9036 644632
rect 9088 644620 9094 644632
rect 487614 644620 487620 644632
rect 9088 644592 487620 644620
rect 9088 644580 9094 644592
rect 487614 644580 487620 644592
rect 487672 644580 487678 644632
rect 25498 644512 25504 644564
rect 25556 644552 25562 644564
rect 512822 644552 512828 644564
rect 25556 644524 512828 644552
rect 25556 644512 25562 644524
rect 512822 644512 512828 644524
rect 512880 644512 512886 644564
rect 8938 644444 8944 644496
rect 8996 644484 9002 644496
rect 500218 644484 500224 644496
rect 8996 644456 500224 644484
rect 8996 644444 9002 644456
rect 500218 644444 500224 644456
rect 500276 644444 500282 644496
rect 209682 644376 209688 644428
rect 209740 644416 209746 644428
rect 523402 644416 523408 644428
rect 209740 644388 523408 644416
rect 209740 644376 209746 644388
rect 523402 644376 523408 644388
rect 523460 644376 523466 644428
rect 3878 644308 3884 644360
rect 3936 644348 3942 644360
rect 191834 644348 191840 644360
rect 3936 644320 191840 644348
rect 3936 644308 3942 644320
rect 191834 644308 191840 644320
rect 191892 644308 191898 644360
rect 197078 644308 197084 644360
rect 197136 644348 197142 644360
rect 523494 644348 523500 644360
rect 197136 644320 523500 644348
rect 197136 644308 197142 644320
rect 523494 644308 523500 644320
rect 523552 644308 523558 644360
rect 184474 644240 184480 644292
rect 184532 644280 184538 644292
rect 523586 644280 523592 644292
rect 184532 644252 523592 644280
rect 184532 644240 184538 644252
rect 523586 644240 523592 644252
rect 523644 644240 523650 644292
rect 192846 644172 192852 644224
rect 192904 644212 192910 644224
rect 531958 644212 531964 644224
rect 192904 644184 531964 644212
rect 192904 644172 192910 644184
rect 531958 644172 531964 644184
rect 532016 644172 532022 644224
rect 176010 644104 176016 644156
rect 176068 644144 176074 644156
rect 524322 644144 524328 644156
rect 176068 644116 524328 644144
rect 176068 644104 176074 644116
rect 524322 644104 524328 644116
rect 524380 644104 524386 644156
rect 8110 644036 8116 644088
rect 8168 644076 8174 644088
rect 361298 644076 361304 644088
rect 8168 644048 361304 644076
rect 8168 644036 8174 644048
rect 361298 644036 361304 644048
rect 361356 644036 361362 644088
rect 8018 643968 8024 644020
rect 8076 644008 8082 644020
rect 373534 644008 373540 644020
rect 8076 643980 373540 644008
rect 8076 643968 8082 643980
rect 373534 643968 373540 643980
rect 373592 643968 373598 644020
rect 140038 643900 140044 643952
rect 140096 643940 140102 643952
rect 580534 643940 580540 643952
rect 140096 643912 580540 643940
rect 140096 643900 140102 643912
rect 580534 643900 580540 643912
rect 580592 643900 580598 643952
rect 146938 643832 146944 643884
rect 146996 643872 147002 643884
rect 524230 643872 524236 643884
rect 146996 643844 524236 643872
rect 146996 643832 147002 643844
rect 524230 643832 524236 643844
rect 524288 643832 524294 643884
rect 9398 643764 9404 643816
rect 9456 643804 9462 643816
rect 402974 643804 402980 643816
rect 9456 643776 402980 643804
rect 9456 643764 9462 643776
rect 402974 643764 402980 643776
rect 403032 643764 403038 643816
rect 125778 643736 125784 643748
rect 125739 643708 125784 643736
rect 125778 643696 125784 643708
rect 125836 643696 125842 643748
rect 172146 643696 172152 643748
rect 172204 643736 172210 643748
rect 567838 643736 567844 643748
rect 172204 643708 567844 643736
rect 172204 643696 172210 643708
rect 567838 643696 567844 643708
rect 567896 643696 567902 643748
rect 117222 643668 117228 643680
rect 117183 643640 117228 643668
rect 117222 643628 117228 643640
rect 117280 643628 117286 643680
rect 121362 643628 121368 643680
rect 121420 643668 121426 643680
rect 524046 643668 524052 643680
rect 121420 643640 524052 643668
rect 121420 643628 121426 643640
rect 524046 643628 524052 643640
rect 524104 643628 524110 643680
rect 3786 643560 3792 643612
rect 3844 643600 3850 643612
rect 419902 643600 419908 643612
rect 3844 643572 419908 643600
rect 3844 643560 3850 643572
rect 419902 643560 419908 643572
rect 419960 643560 419966 643612
rect 96338 643492 96344 643544
rect 96396 643532 96402 643544
rect 523862 643532 523868 643544
rect 96396 643504 523868 643532
rect 96396 643492 96402 643504
rect 523862 643492 523868 643504
rect 523920 643492 523926 643544
rect 92106 643424 92112 643476
rect 92164 643464 92170 643476
rect 525058 643464 525064 643476
rect 92164 643436 525064 643464
rect 92164 643424 92170 643436
rect 525058 643424 525064 643436
rect 525116 643424 525122 643476
rect 79594 643396 79600 643408
rect 79555 643368 79600 643396
rect 79594 643356 79600 643368
rect 79652 643356 79658 643408
rect 87874 643356 87880 643408
rect 87932 643396 87938 643408
rect 523770 643396 523776 643408
rect 87932 643368 523776 643396
rect 87932 643356 87938 643368
rect 523770 643356 523776 643368
rect 523828 643356 523834 643408
rect 45830 643288 45836 643340
rect 45888 643288 45894 643340
rect 58434 643288 58440 643340
rect 58492 643328 58498 643340
rect 522390 643328 522396 643340
rect 58492 643300 522396 643328
rect 58492 643288 58498 643300
rect 522390 643288 522396 643300
rect 522448 643288 522454 643340
rect 45848 643192 45876 643288
rect 117225 643263 117283 643269
rect 117225 643229 117237 643263
rect 117271 643260 117283 643263
rect 580626 643260 580632 643272
rect 117271 643232 580632 643260
rect 117271 643229 117283 643232
rect 117225 643223 117283 643229
rect 580626 643220 580632 643232
rect 580684 643220 580690 643272
rect 522298 643192 522304 643204
rect 45848 643164 522304 643192
rect 522298 643152 522304 643164
rect 522356 643152 522362 643204
rect 79597 643127 79655 643133
rect 79597 643093 79609 643127
rect 79643 643124 79655 643127
rect 580442 643124 580448 643136
rect 79643 643096 580448 643124
rect 79643 643093 79655 643096
rect 79597 643087 79655 643093
rect 580442 643084 580448 643096
rect 580500 643084 580506 643136
rect 125781 641767 125839 641773
rect 125781 641733 125793 641767
rect 125827 641764 125839 641767
rect 580350 641764 580356 641776
rect 125827 641736 580356 641764
rect 125827 641733 125839 641736
rect 125781 641727 125839 641733
rect 580350 641724 580356 641736
rect 580408 641724 580414 641776
rect 571978 640228 571984 640280
rect 572036 640268 572042 640280
rect 580166 640268 580172 640280
rect 572036 640240 580172 640268
rect 572036 640228 572042 640240
rect 580166 640228 580172 640240
rect 580224 640228 580230 640280
rect 523402 627852 523408 627904
rect 523460 627892 523466 627904
rect 579798 627892 579804 627904
rect 523460 627864 579804 627892
rect 523460 627852 523466 627864
rect 579798 627852 579804 627864
rect 579856 627852 579862 627904
rect 3326 624860 3332 624912
rect 3384 624900 3390 624912
rect 8110 624900 8116 624912
rect 3384 624872 8116 624900
rect 3384 624860 3390 624872
rect 8110 624860 8116 624872
rect 8168 624860 8174 624912
rect 3326 611260 3332 611312
rect 3384 611300 3390 611312
rect 10410 611300 10416 611312
rect 3384 611272 10416 611300
rect 3384 611260 3390 611272
rect 10410 611260 10416 611272
rect 10468 611260 10474 611312
rect 544378 593308 544384 593360
rect 544436 593348 544442 593360
rect 579982 593348 579988 593360
rect 544436 593320 579988 593348
rect 544436 593308 544442 593320
rect 579982 593308 579988 593320
rect 580040 593308 580046 593360
rect 523494 580932 523500 580984
rect 523552 580972 523558 580984
rect 579798 580972 579804 580984
rect 523552 580944 579804 580972
rect 523552 580932 523558 580944
rect 579798 580932 579804 580944
rect 579856 580932 579862 580984
rect 3234 568080 3240 568132
rect 3292 568120 3298 568132
rect 8018 568120 8024 568132
rect 3292 568092 8024 568120
rect 3292 568080 3298 568092
rect 8018 568080 8024 568092
rect 8076 568080 8082 568132
rect 2774 553052 2780 553104
rect 2832 553092 2838 553104
rect 5074 553092 5080 553104
rect 2832 553064 5080 553092
rect 2832 553052 2838 553064
rect 5074 553052 5080 553064
rect 5132 553052 5138 553104
rect 531958 546388 531964 546440
rect 532016 546428 532022 546440
rect 579982 546428 579988 546440
rect 532016 546400 579988 546428
rect 532016 546388 532022 546400
rect 579982 546388 579988 546400
rect 580040 546388 580046 546440
rect 3050 539520 3056 539572
rect 3108 539560 3114 539572
rect 25590 539560 25596 539572
rect 3108 539532 25596 539560
rect 3108 539520 3114 539532
rect 25590 539520 25596 539532
rect 25648 539520 25654 539572
rect 523586 534012 523592 534064
rect 523644 534052 523650 534064
rect 579798 534052 579804 534064
rect 523644 534024 579804 534052
rect 523644 534012 523650 534024
rect 579798 534012 579804 534024
rect 579856 534012 579862 534064
rect 524322 510552 524328 510604
rect 524380 510592 524386 510604
rect 580166 510592 580172 510604
rect 524380 510564 580172 510592
rect 524380 510552 524386 510564
rect 580166 510552 580172 510564
rect 580224 510552 580230 510604
rect 3326 509940 3332 509992
rect 3384 509980 3390 509992
rect 7926 509980 7932 509992
rect 3384 509952 7932 509980
rect 3384 509940 3390 509952
rect 7926 509940 7932 509952
rect 7984 509940 7990 509992
rect 3326 495524 3332 495576
rect 3384 495564 3390 495576
rect 8846 495564 8852 495576
rect 3384 495536 8852 495564
rect 3384 495524 3390 495536
rect 8846 495524 8852 495536
rect 8904 495524 8910 495576
rect 567838 487092 567844 487144
rect 567896 487132 567902 487144
rect 579614 487132 579620 487144
rect 567896 487104 579620 487132
rect 567896 487092 567902 487104
rect 579614 487092 579620 487104
rect 579672 487092 579678 487144
rect 3326 481108 3332 481160
rect 3384 481148 3390 481160
rect 9490 481148 9496 481160
rect 3384 481120 9496 481148
rect 3384 481108 3390 481120
rect 9490 481108 9496 481120
rect 9548 481108 9554 481160
rect 553302 462476 553308 462528
rect 553360 462516 553366 462528
rect 560202 462516 560208 462528
rect 553360 462488 560208 462516
rect 553360 462476 553366 462488
rect 560202 462476 560208 462488
rect 560260 462476 560266 462528
rect 522666 452548 522672 452600
rect 522724 452588 522730 452600
rect 579982 452588 579988 452600
rect 522724 452560 579988 452588
rect 522724 452548 522730 452560
rect 579982 452548 579988 452560
rect 580040 452548 580046 452600
rect 3326 452480 3332 452532
rect 3384 452520 3390 452532
rect 7834 452520 7840 452532
rect 3384 452492 7840 452520
rect 3384 452480 3390 452492
rect 7834 452480 7840 452492
rect 7892 452480 7898 452532
rect 525610 440172 525616 440224
rect 525668 440212 525674 440224
rect 579614 440212 579620 440224
rect 525668 440184 579620 440212
rect 525668 440172 525674 440184
rect 579614 440172 579620 440184
rect 579672 440172 579678 440224
rect 3326 424056 3332 424108
rect 3384 424096 3390 424108
rect 9398 424096 9404 424108
rect 3384 424068 9404 424096
rect 3384 424056 3390 424068
rect 9398 424056 9404 424068
rect 9456 424056 9462 424108
rect 525518 416712 525524 416764
rect 525576 416752 525582 416764
rect 580166 416752 580172 416764
rect 525576 416724 580172 416752
rect 525576 416712 525582 416724
rect 580166 416712 580172 416724
rect 580224 416712 580230 416764
rect 537478 405628 537484 405680
rect 537536 405668 537542 405680
rect 579982 405668 579988 405680
rect 537536 405640 579988 405668
rect 537536 405628 537542 405640
rect 579982 405628 579988 405640
rect 580040 405628 580046 405680
rect 3050 395224 3056 395276
rect 3108 395264 3114 395276
rect 7742 395264 7748 395276
rect 3108 395236 7748 395264
rect 3108 395224 3114 395236
rect 7742 395224 7748 395236
rect 7800 395224 7806 395276
rect 524230 393252 524236 393304
rect 524288 393292 524294 393304
rect 579614 393292 579620 393304
rect 524288 393264 579620 393292
rect 524288 393252 524294 393264
rect 579614 393252 579620 393264
rect 579672 393252 579678 393304
rect 525426 369792 525432 369844
rect 525484 369832 525490 369844
rect 580166 369832 580172 369844
rect 525484 369804 580172 369832
rect 525484 369792 525490 369804
rect 580166 369792 580172 369804
rect 580224 369792 580230 369844
rect 3142 367004 3148 367056
rect 3200 367044 3206 367056
rect 40678 367044 40684 367056
rect 3200 367016 40684 367044
rect 3200 367004 3206 367016
rect 40678 367004 40684 367016
rect 40736 367004 40742 367056
rect 525334 358708 525340 358760
rect 525392 358748 525398 358760
rect 579982 358748 579988 358760
rect 525392 358720 579988 358748
rect 525392 358708 525398 358720
rect 579982 358708 579988 358720
rect 580040 358708 580046 358760
rect 524138 346332 524144 346384
rect 524196 346372 524202 346384
rect 579614 346372 579620 346384
rect 524196 346344 579620 346372
rect 524196 346332 524202 346344
rect 579614 346332 579620 346344
rect 579672 346332 579678 346384
rect 3142 337764 3148 337816
rect 3200 337804 3206 337816
rect 7650 337804 7656 337816
rect 3200 337776 7656 337804
rect 3200 337764 3206 337776
rect 7650 337764 7656 337776
rect 7708 337764 7714 337816
rect 525242 311788 525248 311840
rect 525300 311828 525306 311840
rect 580166 311828 580172 311840
rect 525300 311800 580172 311828
rect 525300 311788 525306 311800
rect 580166 311788 580172 311800
rect 580224 311788 580230 311840
rect 3326 308796 3332 308848
rect 3384 308836 3390 308848
rect 9306 308836 9312 308848
rect 3384 308808 9312 308836
rect 3384 308796 3390 308808
rect 9306 308796 9312 308808
rect 9364 308796 9370 308848
rect 524046 299412 524052 299464
rect 524104 299452 524110 299464
rect 580166 299452 580172 299464
rect 524104 299424 580172 299452
rect 524104 299412 524110 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 3602 294924 3608 294976
rect 3660 294964 3666 294976
rect 9214 294964 9220 294976
rect 3660 294936 9220 294964
rect 3660 294924 3666 294936
rect 9214 294924 9220 294936
rect 9272 294924 9278 294976
rect 3234 280100 3240 280152
rect 3292 280140 3298 280152
rect 6454 280140 6460 280152
rect 3292 280112 6460 280140
rect 3292 280100 3298 280112
rect 6454 280100 6460 280112
rect 6512 280100 6518 280152
rect 553302 274796 553308 274848
rect 553360 274836 553366 274848
rect 560202 274836 560208 274848
rect 553360 274808 560208 274836
rect 553360 274796 553366 274808
rect 560202 274796 560208 274808
rect 560260 274796 560266 274848
rect 2774 266160 2780 266212
rect 2832 266200 2838 266212
rect 4982 266200 4988 266212
rect 2832 266172 4988 266200
rect 2832 266160 2838 266172
rect 4982 266160 4988 266172
rect 5040 266160 5046 266212
rect 523954 252492 523960 252544
rect 524012 252532 524018 252544
rect 579706 252532 579712 252544
rect 524012 252504 579712 252532
rect 524012 252492 524018 252504
rect 579706 252492 579712 252504
rect 579764 252492 579770 252544
rect 3142 251268 3148 251320
rect 3200 251308 3206 251320
rect 6362 251308 6368 251320
rect 3200 251280 6368 251308
rect 3200 251268 3206 251280
rect 6362 251268 6368 251280
rect 6420 251268 6426 251320
rect 3142 237056 3148 237108
rect 3200 237096 3206 237108
rect 6270 237096 6276 237108
rect 3200 237068 6276 237096
rect 3200 237056 3206 237068
rect 6270 237056 6276 237068
rect 6328 237056 6334 237108
rect 525150 229032 525156 229084
rect 525208 229072 525214 229084
rect 580166 229072 580172 229084
rect 525208 229044 580172 229072
rect 525208 229032 525214 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 3326 208156 3332 208208
rect 3384 208196 3390 208208
rect 7558 208196 7564 208208
rect 3384 208168 7564 208196
rect 3384 208156 3390 208168
rect 7558 208156 7564 208168
rect 7616 208156 7622 208208
rect 523862 205572 523868 205624
rect 523920 205612 523926 205624
rect 580166 205612 580172 205624
rect 523920 205584 580172 205612
rect 523920 205572 523926 205584
rect 580166 205572 580172 205584
rect 580224 205572 580230 205624
rect 3050 193944 3056 193996
rect 3108 193984 3114 193996
rect 6178 193984 6184 193996
rect 3108 193956 6184 193984
rect 3108 193944 3114 193956
rect 6178 193944 6184 193956
rect 6236 193944 6242 193996
rect 523770 182112 523776 182164
rect 523828 182152 523834 182164
rect 580166 182152 580172 182164
rect 523828 182124 580172 182152
rect 523828 182112 523834 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 2774 179460 2780 179512
rect 2832 179500 2838 179512
rect 4890 179500 4896 179512
rect 2832 179472 4896 179500
rect 2832 179460 2838 179472
rect 4890 179460 4896 179472
rect 4948 179460 4954 179512
rect 525058 171028 525064 171080
rect 525116 171068 525122 171080
rect 580166 171068 580172 171080
rect 525116 171040 580172 171068
rect 525116 171028 525122 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 3142 165180 3148 165232
rect 3200 165220 3206 165232
rect 9122 165220 9128 165232
rect 3200 165192 9128 165220
rect 3200 165180 3206 165192
rect 9122 165180 9128 165192
rect 9180 165180 9186 165232
rect 522574 158652 522580 158704
rect 522632 158692 522638 158704
rect 580166 158692 580172 158704
rect 522632 158664 580172 158692
rect 522632 158652 522638 158664
rect 580166 158652 580172 158664
rect 580224 158652 580230 158704
rect 3326 151716 3332 151768
rect 3384 151756 3390 151768
rect 10318 151756 10324 151768
rect 3384 151728 10324 151756
rect 3384 151716 3390 151728
rect 10318 151716 10324 151728
rect 10376 151716 10382 151768
rect 523678 135192 523684 135244
rect 523736 135232 523742 135244
rect 580166 135232 580172 135244
rect 523736 135204 580172 135232
rect 523736 135192 523742 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 2958 122748 2964 122800
rect 3016 122788 3022 122800
rect 9030 122788 9036 122800
rect 3016 122760 9036 122788
rect 3016 122748 3022 122760
rect 9030 122748 9036 122760
rect 9088 122748 9094 122800
rect 522482 111732 522488 111784
rect 522540 111772 522546 111784
rect 579614 111772 579620 111784
rect 522540 111744 579620 111772
rect 522540 111732 522546 111744
rect 579614 111732 579620 111744
rect 579672 111732 579678 111784
rect 3234 108944 3240 108996
rect 3292 108984 3298 108996
rect 13078 108984 13084 108996
rect 3292 108956 13084 108984
rect 3292 108944 3298 108956
rect 13078 108944 13084 108956
rect 13136 108944 13142 108996
rect 2774 93236 2780 93288
rect 2832 93276 2838 93288
rect 4798 93276 4804 93288
rect 2832 93248 4804 93276
rect 2832 93236 2838 93248
rect 4798 93236 4804 93248
rect 4856 93236 4862 93288
rect 553302 87116 553308 87168
rect 553360 87156 553366 87168
rect 560202 87156 560208 87168
rect 553360 87128 560208 87156
rect 553360 87116 553366 87128
rect 560202 87116 560208 87128
rect 560260 87116 560266 87168
rect 3050 79840 3056 79892
rect 3108 79880 3114 79892
rect 8938 79880 8944 79892
rect 3108 79852 8944 79880
rect 3108 79840 3114 79852
rect 8938 79840 8944 79852
rect 8996 79840 9002 79892
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 14458 64852 14464 64864
rect 3384 64824 14464 64852
rect 3384 64812 3390 64824
rect 14458 64812 14464 64824
rect 14516 64812 14522 64864
rect 522482 64812 522488 64864
rect 522540 64852 522546 64864
rect 580166 64852 580172 64864
rect 522540 64824 580172 64852
rect 522540 64812 522546 64824
rect 580166 64812 580172 64824
rect 580224 64812 580230 64864
rect 129384 42860 129688 42888
rect 69014 42820 69020 42832
rect 68848 42792 69020 42820
rect 21910 42712 21916 42764
rect 21968 42752 21974 42764
rect 60550 42752 60556 42764
rect 21968 42724 60556 42752
rect 21968 42712 21974 42724
rect 60550 42712 60556 42724
rect 60608 42712 60614 42764
rect 60645 42755 60703 42761
rect 60645 42721 60657 42755
rect 60691 42752 60703 42755
rect 67450 42752 67456 42764
rect 60691 42724 67456 42752
rect 60691 42721 60703 42724
rect 60645 42715 60703 42721
rect 67450 42712 67456 42724
rect 67508 42712 67514 42764
rect 67545 42755 67603 42761
rect 67545 42721 67557 42755
rect 67591 42752 67603 42755
rect 68848 42752 68876 42792
rect 69014 42780 69020 42792
rect 69072 42780 69078 42832
rect 74445 42823 74503 42829
rect 74445 42820 74457 42823
rect 74276 42792 74457 42820
rect 67591 42724 68876 42752
rect 67591 42721 67603 42724
rect 67545 42715 67603 42721
rect 68922 42712 68928 42764
rect 68980 42752 68986 42764
rect 74276 42752 74304 42792
rect 74445 42789 74457 42792
rect 74491 42789 74503 42823
rect 74445 42783 74503 42789
rect 68980 42724 74304 42752
rect 74353 42755 74411 42761
rect 68980 42712 68986 42724
rect 74353 42721 74365 42755
rect 74399 42752 74411 42755
rect 98822 42752 98828 42764
rect 74399 42724 98828 42752
rect 74399 42721 74411 42724
rect 74353 42715 74411 42721
rect 98822 42712 98828 42724
rect 98880 42712 98886 42764
rect 107562 42712 107568 42764
rect 107620 42752 107626 42764
rect 129384 42752 129412 42860
rect 107620 42724 129412 42752
rect 129660 42752 129688 42860
rect 129737 42823 129795 42829
rect 129737 42789 129749 42823
rect 129783 42820 129795 42823
rect 129783 42792 131436 42820
rect 129783 42789 129795 42792
rect 129737 42783 129795 42789
rect 131206 42752 131212 42764
rect 129660 42724 131212 42752
rect 107620 42712 107626 42724
rect 131206 42712 131212 42724
rect 131264 42712 131270 42764
rect 23382 42644 23388 42696
rect 23440 42684 23446 42696
rect 62574 42684 62580 42696
rect 23440 42656 62580 42684
rect 23440 42644 23446 42656
rect 62574 42644 62580 42656
rect 62632 42644 62638 42696
rect 64782 42644 64788 42696
rect 64840 42684 64846 42696
rect 95878 42684 95884 42696
rect 64840 42656 73568 42684
rect 64840 42644 64846 42656
rect 19242 42576 19248 42628
rect 19300 42616 19306 42628
rect 58618 42616 58624 42628
rect 19300 42588 58624 42616
rect 19300 42576 19306 42588
rect 58618 42576 58624 42588
rect 58676 42576 58682 42628
rect 59909 42619 59967 42625
rect 59909 42585 59921 42619
rect 59955 42616 59967 42619
rect 60553 42619 60611 42625
rect 60553 42616 60565 42619
rect 59955 42588 60565 42616
rect 59955 42585 59967 42588
rect 59909 42579 59967 42585
rect 60553 42585 60565 42588
rect 60599 42585 60611 42619
rect 60553 42579 60611 42585
rect 60642 42576 60648 42628
rect 60700 42616 60706 42628
rect 66809 42619 66867 42625
rect 60700 42588 66300 42616
rect 60700 42576 60706 42588
rect 20622 42508 20628 42560
rect 20680 42548 20686 42560
rect 59630 42548 59636 42560
rect 20680 42520 59636 42548
rect 20680 42508 20686 42520
rect 59630 42508 59636 42520
rect 59688 42508 59694 42560
rect 59817 42551 59875 42557
rect 59817 42517 59829 42551
rect 59863 42548 59875 42551
rect 66162 42548 66168 42560
rect 59863 42520 66168 42548
rect 59863 42517 59875 42520
rect 59817 42511 59875 42517
rect 66162 42508 66168 42520
rect 66220 42508 66226 42560
rect 66272 42548 66300 42588
rect 66809 42585 66821 42619
rect 66855 42616 66867 42619
rect 72326 42616 72332 42628
rect 66855 42588 72332 42616
rect 66855 42585 66867 42588
rect 66809 42579 66867 42585
rect 72326 42576 72332 42588
rect 72384 42576 72390 42628
rect 73540 42616 73568 42656
rect 74368 42656 95884 42684
rect 74368 42616 74396 42656
rect 95878 42644 95884 42656
rect 95936 42644 95942 42696
rect 99282 42644 99288 42696
rect 99340 42684 99346 42696
rect 125226 42684 125232 42696
rect 99340 42656 125232 42684
rect 99340 42644 99346 42656
rect 125226 42644 125232 42656
rect 125284 42644 125290 42696
rect 125321 42687 125379 42693
rect 125321 42653 125333 42687
rect 125367 42684 125379 42687
rect 129553 42687 129611 42693
rect 129553 42684 129565 42687
rect 125367 42656 129565 42684
rect 125367 42653 125379 42656
rect 125321 42647 125379 42653
rect 129553 42653 129565 42656
rect 129599 42653 129611 42687
rect 129553 42647 129611 42653
rect 129642 42644 129648 42696
rect 129700 42684 129706 42696
rect 131408 42684 131436 42792
rect 135088 42792 136128 42820
rect 133782 42712 133788 42764
rect 133840 42752 133846 42764
rect 135088 42752 135116 42792
rect 133840 42724 135116 42752
rect 136100 42752 136128 42792
rect 153654 42752 153660 42764
rect 136100 42724 153660 42752
rect 133840 42712 133846 42724
rect 153654 42712 153660 42724
rect 153712 42712 153718 42764
rect 154482 42712 154488 42764
rect 154540 42752 154546 42764
rect 170306 42752 170312 42764
rect 154540 42724 170312 42752
rect 154540 42712 154546 42724
rect 170306 42712 170312 42724
rect 170364 42712 170370 42764
rect 173802 42712 173808 42764
rect 173860 42752 173866 42764
rect 185946 42752 185952 42764
rect 173860 42724 185952 42752
rect 173860 42712 173866 42724
rect 185946 42712 185952 42724
rect 186004 42712 186010 42764
rect 190362 42712 190368 42764
rect 190420 42752 190426 42764
rect 199654 42752 199660 42764
rect 190420 42724 199660 42752
rect 190420 42712 190426 42724
rect 199654 42712 199660 42724
rect 199712 42712 199718 42764
rect 237282 42712 237288 42764
rect 237340 42752 237346 42764
rect 238846 42752 238852 42764
rect 237340 42724 238852 42752
rect 237340 42712 237346 42724
rect 238846 42712 238852 42724
rect 238904 42712 238910 42764
rect 240042 42712 240048 42764
rect 240100 42752 240106 42764
rect 240870 42752 240876 42764
rect 240100 42724 240876 42752
rect 240100 42712 240106 42724
rect 240870 42712 240876 42724
rect 240928 42712 240934 42764
rect 251634 42712 251640 42764
rect 251692 42752 251698 42764
rect 252462 42752 252468 42764
rect 251692 42724 252468 42752
rect 251692 42712 251698 42724
rect 252462 42712 252468 42724
rect 252520 42712 252526 42764
rect 382826 42712 382832 42764
rect 382884 42752 382890 42764
rect 411438 42752 411444 42764
rect 382884 42724 411444 42752
rect 382884 42712 382890 42724
rect 411438 42712 411444 42724
rect 411496 42712 411502 42764
rect 414198 42712 414204 42764
rect 414256 42752 414262 42764
rect 422938 42752 422944 42764
rect 414256 42724 422944 42752
rect 414256 42712 414262 42724
rect 422938 42712 422944 42724
rect 422996 42712 423002 42764
rect 455322 42712 455328 42764
rect 455380 42752 455386 42764
rect 499666 42752 499672 42764
rect 455380 42724 499672 42752
rect 455380 42712 455386 42724
rect 499666 42712 499672 42724
rect 499724 42712 499730 42764
rect 502334 42712 502340 42764
rect 502392 42752 502398 42764
rect 542998 42752 543004 42764
rect 502392 42724 543004 42752
rect 502392 42712 502398 42724
rect 542998 42712 543004 42724
rect 543056 42712 543062 42764
rect 134058 42684 134064 42696
rect 129700 42656 131252 42684
rect 131408 42656 134064 42684
rect 129700 42644 129706 42656
rect 73540 42588 74396 42616
rect 74445 42619 74503 42625
rect 74445 42585 74457 42619
rect 74491 42616 74503 42619
rect 99742 42616 99748 42628
rect 74491 42588 99748 42616
rect 74491 42585 74503 42588
rect 74445 42579 74503 42585
rect 99742 42576 99748 42588
rect 99800 42576 99806 42628
rect 107470 42576 107476 42628
rect 107528 42616 107534 42628
rect 131114 42616 131120 42628
rect 107528 42588 131120 42616
rect 107528 42576 107534 42588
rect 131114 42576 131120 42588
rect 131172 42576 131178 42628
rect 131224 42616 131252 42656
rect 134058 42644 134064 42656
rect 134116 42644 134122 42696
rect 149698 42684 149704 42696
rect 135916 42656 149704 42684
rect 135916 42616 135944 42656
rect 149698 42644 149704 42656
rect 149756 42644 149762 42696
rect 151630 42644 151636 42696
rect 151688 42684 151694 42696
rect 167362 42684 167368 42696
rect 151688 42656 167368 42684
rect 151688 42644 151694 42656
rect 167362 42644 167368 42656
rect 167420 42644 167426 42696
rect 169662 42644 169668 42696
rect 169720 42684 169726 42696
rect 183002 42684 183008 42696
rect 169720 42656 183008 42684
rect 169720 42644 169726 42656
rect 183002 42644 183008 42656
rect 183060 42644 183066 42696
rect 183462 42644 183468 42696
rect 183520 42684 183526 42696
rect 193766 42684 193772 42696
rect 183520 42656 193772 42684
rect 183520 42644 183526 42656
rect 193766 42644 193772 42656
rect 193824 42644 193830 42696
rect 399478 42644 399484 42696
rect 399536 42684 399542 42696
rect 402238 42684 402244 42696
rect 399536 42656 402244 42684
rect 399536 42644 399542 42656
rect 402238 42644 402244 42656
rect 402296 42644 402302 42696
rect 403434 42644 403440 42696
rect 403492 42684 403498 42696
rect 404262 42684 404268 42696
rect 403492 42656 404268 42684
rect 403492 42644 403498 42656
rect 404262 42644 404268 42656
rect 404320 42644 404326 42696
rect 404446 42644 404452 42696
rect 404504 42684 404510 42696
rect 405642 42684 405648 42696
rect 404504 42656 405648 42684
rect 404504 42644 404510 42656
rect 405642 42644 405648 42656
rect 405700 42644 405706 42696
rect 417418 42684 417424 42696
rect 406948 42656 417424 42684
rect 131224 42588 135944 42616
rect 136177 42619 136235 42625
rect 136177 42585 136189 42619
rect 136223 42616 136235 42619
rect 154666 42616 154672 42628
rect 136223 42588 154672 42616
rect 136223 42585 136235 42588
rect 136177 42579 136235 42585
rect 154666 42576 154672 42588
rect 154724 42576 154730 42628
rect 155862 42576 155868 42628
rect 155920 42616 155926 42628
rect 171318 42616 171324 42628
rect 155920 42588 171324 42616
rect 155920 42576 155926 42588
rect 171318 42576 171324 42588
rect 171376 42576 171382 42628
rect 172422 42576 172428 42628
rect 172480 42616 172486 42628
rect 185026 42616 185032 42628
rect 172480 42588 185032 42616
rect 172480 42576 172486 42588
rect 185026 42576 185032 42588
rect 185084 42576 185090 42628
rect 186222 42576 186228 42628
rect 186280 42616 186286 42628
rect 196710 42616 196716 42628
rect 186280 42588 196716 42616
rect 186280 42576 186286 42588
rect 196710 42576 196716 42588
rect 196768 42576 196774 42628
rect 197262 42576 197268 42628
rect 197320 42616 197326 42628
rect 205542 42616 205548 42628
rect 197320 42588 205548 42616
rect 197320 42576 197326 42588
rect 205542 42576 205548 42588
rect 205600 42576 205606 42628
rect 365254 42576 365260 42628
rect 365312 42616 365318 42628
rect 390646 42616 390652 42628
rect 365312 42588 390652 42616
rect 365312 42576 365318 42588
rect 390646 42576 390652 42588
rect 390704 42576 390710 42628
rect 405366 42576 405372 42628
rect 405424 42616 405430 42628
rect 406948 42616 406976 42656
rect 417418 42644 417424 42656
rect 417476 42644 417482 42696
rect 461210 42644 461216 42696
rect 461268 42684 461274 42696
rect 506474 42684 506480 42696
rect 461268 42656 506480 42684
rect 461268 42644 461274 42656
rect 506474 42644 506480 42656
rect 506532 42644 506538 42696
rect 508222 42644 508228 42696
rect 508280 42684 508286 42696
rect 544378 42684 544384 42696
rect 508280 42656 544384 42684
rect 508280 42644 508286 42656
rect 544378 42644 544384 42656
rect 544436 42644 544442 42696
rect 433978 42616 433984 42628
rect 405424 42588 406976 42616
rect 408420 42588 433984 42616
rect 405424 42576 405430 42588
rect 92934 42548 92940 42560
rect 66272 42520 92940 42548
rect 92934 42508 92940 42520
rect 92992 42508 92998 42560
rect 96522 42508 96528 42560
rect 96580 42548 96586 42560
rect 122282 42548 122288 42560
rect 96580 42520 122288 42548
rect 96580 42508 96586 42520
rect 122282 42508 122288 42520
rect 122340 42508 122346 42560
rect 142890 42548 142896 42560
rect 122392 42520 142896 42548
rect 9582 42440 9588 42492
rect 9640 42480 9646 42492
rect 50798 42480 50804 42492
rect 9640 42452 50804 42480
rect 9640 42440 9646 42452
rect 50798 42440 50804 42452
rect 50856 42440 50862 42492
rect 50982 42440 50988 42492
rect 51040 42480 51046 42492
rect 60001 42483 60059 42489
rect 60001 42480 60013 42483
rect 51040 42452 60013 42480
rect 51040 42440 51046 42452
rect 60001 42449 60013 42452
rect 60047 42449 60059 42483
rect 60001 42443 60059 42449
rect 60093 42483 60151 42489
rect 60093 42449 60105 42483
rect 60139 42480 60151 42483
rect 91002 42480 91008 42492
rect 60139 42452 91008 42480
rect 60139 42449 60151 42452
rect 60093 42443 60151 42449
rect 91002 42440 91008 42452
rect 91060 42440 91066 42492
rect 92382 42440 92388 42492
rect 92440 42480 92446 42492
rect 119338 42480 119344 42492
rect 92440 42452 119344 42480
rect 92440 42440 92446 42452
rect 119338 42440 119344 42452
rect 119396 42440 119402 42492
rect 120445 42483 120503 42489
rect 120445 42480 120457 42483
rect 119448 42452 120457 42480
rect 13630 42372 13636 42424
rect 13688 42412 13694 42424
rect 54754 42412 54760 42424
rect 13688 42384 54760 42412
rect 13688 42372 13694 42384
rect 54754 42372 54760 42384
rect 54812 42372 54818 42424
rect 55122 42372 55128 42424
rect 55180 42412 55186 42424
rect 88058 42412 88064 42424
rect 55180 42384 88064 42412
rect 55180 42372 55186 42384
rect 88058 42372 88064 42384
rect 88116 42372 88122 42424
rect 89622 42372 89628 42424
rect 89680 42412 89686 42424
rect 116394 42412 116400 42424
rect 89680 42384 116400 42412
rect 89680 42372 89686 42384
rect 116394 42372 116400 42384
rect 116452 42372 116458 42424
rect 117041 42415 117099 42421
rect 117041 42381 117053 42415
rect 117087 42412 117099 42415
rect 119448 42412 119476 42452
rect 120445 42449 120457 42452
rect 120491 42449 120503 42483
rect 120445 42443 120503 42449
rect 121362 42440 121368 42492
rect 121420 42480 121426 42492
rect 122392 42480 122420 42520
rect 142890 42508 142896 42520
rect 142948 42508 142954 42560
rect 144638 42508 144644 42560
rect 144696 42548 144702 42560
rect 162486 42548 162492 42560
rect 144696 42520 162492 42548
rect 144696 42508 144702 42520
rect 162486 42508 162492 42520
rect 162544 42508 162550 42560
rect 168282 42508 168288 42560
rect 168340 42548 168346 42560
rect 181070 42548 181076 42560
rect 168340 42520 181076 42548
rect 168340 42508 168346 42520
rect 181070 42508 181076 42520
rect 181128 42508 181134 42560
rect 182174 42508 182180 42560
rect 182232 42548 182238 42560
rect 192846 42548 192852 42560
rect 182232 42520 192852 42548
rect 182232 42508 182238 42520
rect 192846 42508 192852 42520
rect 192904 42508 192910 42560
rect 347590 42508 347596 42560
rect 347648 42548 347654 42560
rect 368566 42548 368572 42560
rect 347648 42520 368572 42548
rect 347648 42508 347654 42520
rect 368566 42508 368572 42520
rect 368624 42508 368630 42560
rect 374086 42508 374092 42560
rect 374144 42548 374150 42560
rect 400398 42548 400404 42560
rect 374144 42520 400404 42548
rect 374144 42508 374150 42520
rect 400398 42508 400404 42520
rect 400456 42508 400462 42560
rect 121420 42452 122420 42480
rect 122469 42483 122527 42489
rect 121420 42440 121426 42452
rect 122469 42449 122481 42483
rect 122515 42480 122527 42483
rect 138934 42480 138940 42492
rect 122515 42452 138940 42480
rect 122515 42449 122527 42452
rect 122469 42443 122527 42449
rect 138934 42440 138940 42452
rect 138992 42440 138998 42492
rect 139302 42440 139308 42492
rect 139360 42480 139366 42492
rect 157610 42480 157616 42492
rect 139360 42452 157616 42480
rect 139360 42440 139366 42452
rect 157610 42440 157616 42452
rect 157668 42440 157674 42492
rect 158622 42440 158628 42492
rect 158680 42480 158686 42492
rect 173250 42480 173256 42492
rect 158680 42452 173256 42480
rect 158680 42440 158686 42452
rect 173250 42440 173256 42452
rect 173308 42440 173314 42492
rect 175182 42440 175188 42492
rect 175240 42480 175246 42492
rect 186958 42480 186964 42492
rect 175240 42452 186964 42480
rect 175240 42440 175246 42452
rect 186958 42440 186964 42452
rect 187016 42440 187022 42492
rect 187602 42440 187608 42492
rect 187660 42480 187666 42492
rect 197722 42480 197728 42492
rect 187660 42452 197728 42480
rect 187660 42440 187666 42452
rect 197722 42440 197728 42452
rect 197780 42440 197786 42492
rect 198642 42440 198648 42492
rect 198700 42480 198706 42492
rect 206554 42480 206560 42492
rect 198700 42452 206560 42480
rect 198700 42440 198706 42452
rect 206554 42440 206560 42452
rect 206612 42440 206618 42492
rect 359366 42440 359372 42492
rect 359424 42480 359430 42492
rect 382458 42480 382464 42492
rect 359424 42452 382464 42480
rect 359424 42440 359430 42452
rect 382458 42440 382464 42452
rect 382516 42440 382522 42492
rect 402422 42440 402428 42492
rect 402480 42480 402486 42492
rect 408420 42480 408448 42588
rect 433978 42576 433984 42588
rect 434036 42576 434042 42628
rect 452378 42576 452384 42628
rect 452436 42616 452442 42628
rect 494698 42616 494704 42628
rect 452436 42588 494704 42616
rect 452436 42576 452442 42588
rect 494698 42576 494704 42588
rect 494756 42576 494762 42628
rect 496446 42576 496452 42628
rect 496504 42616 496510 42628
rect 541618 42616 541624 42628
rect 496504 42588 541624 42616
rect 496504 42576 496510 42588
rect 541618 42576 541624 42588
rect 541676 42576 541682 42628
rect 411254 42508 411260 42560
rect 411312 42548 411318 42560
rect 445754 42548 445760 42560
rect 411312 42520 445760 42548
rect 411312 42508 411318 42520
rect 445754 42508 445760 42520
rect 445812 42508 445818 42560
rect 471974 42508 471980 42560
rect 472032 42548 472038 42560
rect 483658 42548 483664 42560
rect 472032 42520 483664 42548
rect 472032 42508 472038 42520
rect 483658 42508 483664 42520
rect 483716 42508 483722 42560
rect 486694 42508 486700 42560
rect 486752 42548 486758 42560
rect 531958 42548 531964 42560
rect 486752 42520 531964 42548
rect 486752 42508 486758 42520
rect 531958 42508 531964 42520
rect 532016 42508 532022 42560
rect 402480 42452 408448 42480
rect 402480 42440 402486 42452
rect 417142 42440 417148 42492
rect 417200 42480 417206 42492
rect 451918 42480 451924 42492
rect 417200 42452 451924 42480
rect 417200 42440 417206 42452
rect 451918 42440 451924 42452
rect 451976 42440 451982 42492
rect 467098 42440 467104 42492
rect 467156 42480 467162 42492
rect 512638 42480 512644 42492
rect 467156 42452 512644 42480
rect 467156 42440 467162 42452
rect 512638 42440 512644 42452
rect 512696 42440 512702 42492
rect 514110 42440 514116 42492
rect 514168 42480 514174 42492
rect 545758 42480 545764 42492
rect 514168 42452 545764 42480
rect 514168 42440 514174 42452
rect 545758 42440 545764 42452
rect 545816 42440 545822 42492
rect 117087 42384 119476 42412
rect 117087 42381 117099 42384
rect 117041 42375 117099 42381
rect 119982 42372 119988 42424
rect 120040 42412 120046 42424
rect 141878 42412 141884 42424
rect 120040 42384 141884 42412
rect 120040 42372 120046 42384
rect 141878 42372 141884 42384
rect 141936 42372 141942 42424
rect 141970 42372 141976 42424
rect 142028 42412 142034 42424
rect 159542 42412 159548 42424
rect 142028 42384 159548 42412
rect 142028 42372 142034 42384
rect 159542 42372 159548 42384
rect 159600 42372 159606 42424
rect 159910 42372 159916 42424
rect 159968 42412 159974 42424
rect 174262 42412 174268 42424
rect 159968 42384 174268 42412
rect 159968 42372 159974 42384
rect 174262 42372 174268 42384
rect 174320 42372 174326 42424
rect 176470 42372 176476 42424
rect 176528 42412 176534 42424
rect 187970 42412 187976 42424
rect 176528 42384 187976 42412
rect 176528 42372 176534 42384
rect 187970 42372 187976 42384
rect 188028 42372 188034 42424
rect 191742 42372 191748 42424
rect 191800 42412 191806 42424
rect 200666 42412 200672 42424
rect 191800 42384 200672 42412
rect 191800 42372 191806 42384
rect 200666 42372 200672 42384
rect 200724 42372 200730 42424
rect 219342 42372 219348 42424
rect 219400 42412 219406 42424
rect 223206 42412 223212 42424
rect 219400 42384 223212 42412
rect 219400 42372 219406 42384
rect 223206 42372 223212 42384
rect 223264 42372 223270 42424
rect 353478 42372 353484 42424
rect 353536 42412 353542 42424
rect 375466 42412 375472 42424
rect 353536 42384 375472 42412
rect 353536 42372 353542 42384
rect 375466 42372 375472 42384
rect 375524 42372 375530 42424
rect 379882 42372 379888 42424
rect 379940 42412 379946 42424
rect 408586 42412 408592 42424
rect 379940 42384 408592 42412
rect 379940 42372 379946 42384
rect 408586 42372 408592 42384
rect 408644 42372 408650 42424
rect 418154 42372 418160 42424
rect 418212 42412 418218 42424
rect 454126 42412 454132 42424
rect 418212 42384 454132 42412
rect 418212 42372 418218 42384
rect 454126 42372 454132 42384
rect 454184 42372 454190 42424
rect 483750 42372 483756 42424
rect 483808 42412 483814 42424
rect 530578 42412 530584 42424
rect 483808 42384 530584 42412
rect 483808 42372 483814 42384
rect 530578 42372 530584 42384
rect 530636 42372 530642 42424
rect 16482 42304 16488 42356
rect 16540 42344 16546 42356
rect 56686 42344 56692 42356
rect 16540 42316 56692 42344
rect 16540 42304 16546 42316
rect 56686 42304 56692 42316
rect 56744 42304 56750 42356
rect 57882 42304 57888 42356
rect 57940 42344 57946 42356
rect 60093 42347 60151 42353
rect 60093 42344 60105 42347
rect 57940 42316 60105 42344
rect 57940 42304 57946 42316
rect 60093 42313 60105 42316
rect 60139 42313 60151 42347
rect 60093 42307 60151 42313
rect 62022 42304 62028 42356
rect 62080 42344 62086 42356
rect 93854 42344 93860 42356
rect 62080 42316 93860 42344
rect 62080 42304 62086 42316
rect 93854 42304 93860 42316
rect 93912 42304 93918 42356
rect 97902 42304 97908 42356
rect 97960 42344 97966 42356
rect 123294 42344 123300 42356
rect 97960 42316 123300 42344
rect 97960 42304 97966 42316
rect 123294 42304 123300 42316
rect 123352 42304 123358 42356
rect 123849 42347 123907 42353
rect 123849 42313 123861 42347
rect 123895 42344 123907 42347
rect 125321 42347 125379 42353
rect 125321 42344 125333 42347
rect 123895 42316 125333 42344
rect 123895 42313 123907 42316
rect 123849 42307 123907 42313
rect 125321 42313 125333 42316
rect 125367 42313 125379 42347
rect 125321 42307 125379 42313
rect 125410 42304 125416 42356
rect 125468 42344 125474 42356
rect 145834 42344 145840 42356
rect 125468 42316 145840 42344
rect 125468 42304 125474 42316
rect 145834 42304 145840 42316
rect 145892 42304 145898 42356
rect 151722 42304 151728 42356
rect 151780 42344 151786 42356
rect 168374 42344 168380 42356
rect 151780 42316 168380 42344
rect 151780 42304 151786 42316
rect 168374 42304 168380 42316
rect 168432 42304 168438 42356
rect 171042 42304 171048 42356
rect 171100 42344 171106 42356
rect 184014 42344 184020 42356
rect 171100 42316 184020 42344
rect 171100 42304 171106 42316
rect 184014 42304 184020 42316
rect 184072 42304 184078 42356
rect 188982 42304 188988 42356
rect 189040 42344 189046 42356
rect 198734 42344 198740 42356
rect 189040 42316 198740 42344
rect 189040 42304 189046 42316
rect 198734 42304 198740 42316
rect 198792 42304 198798 42356
rect 200022 42304 200028 42356
rect 200080 42344 200086 42356
rect 207566 42344 207572 42356
rect 200080 42316 207572 42344
rect 200080 42304 200086 42316
rect 207566 42304 207572 42316
rect 207624 42304 207630 42356
rect 208302 42304 208308 42356
rect 208360 42344 208366 42356
rect 214374 42344 214380 42356
rect 208360 42316 214380 42344
rect 208360 42304 208366 42316
rect 214374 42304 214380 42316
rect 214432 42304 214438 42356
rect 356422 42304 356428 42356
rect 356480 42344 356486 42356
rect 379514 42344 379520 42356
rect 356480 42316 379520 42344
rect 356480 42304 356486 42316
rect 379514 42304 379520 42316
rect 379572 42304 379578 42356
rect 385770 42304 385776 42356
rect 385828 42344 385834 42356
rect 415486 42344 415492 42356
rect 385828 42316 415492 42344
rect 385828 42304 385834 42316
rect 415486 42304 415492 42316
rect 415544 42304 415550 42356
rect 428918 42304 428924 42356
rect 428976 42344 428982 42356
rect 464338 42344 464344 42356
rect 428976 42316 464344 42344
rect 428976 42304 428982 42316
rect 464338 42304 464344 42316
rect 464396 42304 464402 42356
rect 472986 42304 472992 42356
rect 473044 42344 473050 42356
rect 520458 42344 520464 42356
rect 473044 42316 520464 42344
rect 473044 42304 473050 42316
rect 520458 42304 520464 42316
rect 520516 42304 520522 42356
rect 522942 42304 522948 42356
rect 523000 42344 523006 42356
rect 547230 42344 547236 42356
rect 523000 42316 547236 42344
rect 523000 42304 523006 42316
rect 547230 42304 547236 42316
rect 547288 42304 547294 42356
rect 12342 42236 12348 42288
rect 12400 42276 12406 42288
rect 52730 42276 52736 42288
rect 12400 42248 52736 42276
rect 12400 42236 12406 42248
rect 52730 42236 52736 42248
rect 52788 42236 52794 42288
rect 56502 42236 56508 42288
rect 56560 42276 56566 42288
rect 89990 42276 89996 42288
rect 56560 42248 89996 42276
rect 56560 42236 56566 42248
rect 89990 42236 89996 42248
rect 90048 42236 90054 42288
rect 93762 42236 93768 42288
rect 93820 42276 93826 42288
rect 120350 42276 120356 42288
rect 93820 42248 120356 42276
rect 93820 42236 93826 42248
rect 120350 42236 120356 42248
rect 120408 42236 120414 42288
rect 120445 42279 120503 42285
rect 120445 42245 120457 42279
rect 120491 42276 120503 42279
rect 122653 42279 122711 42285
rect 122653 42276 122665 42279
rect 120491 42248 122665 42276
rect 120491 42245 120503 42248
rect 120445 42239 120503 42245
rect 122653 42245 122665 42248
rect 122699 42245 122711 42279
rect 122653 42239 122711 42245
rect 122742 42236 122748 42288
rect 122800 42276 122806 42288
rect 143810 42276 143816 42288
rect 122800 42248 143816 42276
rect 122800 42236 122806 42248
rect 143810 42236 143816 42248
rect 143868 42236 143874 42288
rect 146202 42236 146208 42288
rect 146260 42276 146266 42288
rect 163406 42276 163412 42288
rect 146260 42248 163412 42276
rect 146260 42236 146266 42248
rect 163406 42236 163412 42248
rect 163464 42236 163470 42288
rect 165522 42236 165528 42288
rect 165580 42276 165586 42288
rect 179138 42276 179144 42288
rect 165580 42248 179144 42276
rect 165580 42236 165586 42248
rect 179138 42236 179144 42248
rect 179196 42236 179202 42288
rect 180702 42236 180708 42288
rect 180760 42276 180766 42288
rect 191834 42276 191840 42288
rect 180760 42248 191840 42276
rect 180760 42236 180766 42248
rect 191834 42236 191840 42248
rect 191892 42236 191898 42288
rect 209682 42236 209688 42288
rect 209740 42276 209746 42288
rect 215386 42276 215392 42288
rect 209740 42248 215392 42276
rect 209740 42236 209746 42248
rect 215386 42236 215392 42248
rect 215444 42236 215450 42288
rect 362310 42236 362316 42288
rect 362368 42276 362374 42288
rect 386506 42276 386512 42288
rect 362368 42248 386512 42276
rect 362368 42236 362374 42248
rect 386506 42236 386512 42248
rect 386564 42236 386570 42288
rect 388714 42236 388720 42288
rect 388772 42276 388778 42288
rect 418246 42276 418252 42288
rect 388772 42248 418252 42276
rect 388772 42236 388778 42248
rect 418246 42236 418252 42248
rect 418304 42236 418310 42288
rect 423030 42236 423036 42288
rect 423088 42276 423094 42288
rect 459646 42276 459652 42288
rect 423088 42248 459652 42276
rect 423088 42236 423094 42248
rect 459646 42236 459652 42248
rect 459704 42236 459710 42288
rect 469030 42236 469036 42288
rect 469088 42276 469094 42288
rect 478138 42276 478144 42288
rect 469088 42248 478144 42276
rect 469088 42236 469094 42248
rect 478138 42236 478144 42248
rect 478196 42236 478202 42288
rect 478874 42236 478880 42288
rect 478932 42276 478938 42288
rect 528554 42276 528560 42288
rect 478932 42248 528560 42276
rect 478932 42236 478938 42248
rect 528554 42236 528560 42248
rect 528612 42236 528618 42288
rect 10962 42168 10968 42220
rect 11020 42208 11026 42220
rect 51810 42208 51816 42220
rect 11020 42180 51816 42208
rect 11020 42168 11026 42180
rect 51810 42168 51816 42180
rect 51868 42168 51874 42220
rect 53742 42168 53748 42220
rect 53800 42208 53806 42220
rect 87046 42208 87052 42220
rect 53800 42180 87052 42208
rect 53800 42168 53806 42180
rect 87046 42168 87052 42180
rect 87104 42168 87110 42220
rect 91002 42168 91008 42220
rect 91060 42208 91066 42220
rect 117406 42208 117412 42220
rect 91060 42180 117412 42208
rect 91060 42168 91066 42180
rect 117406 42168 117412 42180
rect 117464 42168 117470 42220
rect 117516 42180 125548 42208
rect 4062 42100 4068 42152
rect 4120 42140 4126 42152
rect 46842 42140 46848 42152
rect 4120 42112 46848 42140
rect 4120 42100 4126 42112
rect 46842 42100 46848 42112
rect 46900 42100 46906 42152
rect 46934 42100 46940 42152
rect 46992 42140 46998 42152
rect 81158 42140 81164 42152
rect 46992 42112 81164 42140
rect 46992 42100 46998 42112
rect 81158 42100 81164 42112
rect 81216 42100 81222 42152
rect 82722 42100 82728 42152
rect 82780 42140 82786 42152
rect 110506 42140 110512 42152
rect 82780 42112 110512 42140
rect 82780 42100 82786 42112
rect 110506 42100 110512 42112
rect 110564 42100 110570 42152
rect 113177 42143 113235 42149
rect 113177 42109 113189 42143
rect 113223 42140 113235 42143
rect 117041 42143 117099 42149
rect 117041 42140 117053 42143
rect 113223 42112 117053 42140
rect 113223 42109 113235 42112
rect 113177 42103 113235 42109
rect 117041 42109 117053 42112
rect 117087 42109 117099 42143
rect 117041 42103 117099 42109
rect 117130 42100 117136 42152
rect 117188 42140 117194 42152
rect 117516 42140 117544 42180
rect 117188 42112 117544 42140
rect 117188 42100 117194 42112
rect 118602 42100 118608 42152
rect 118660 42140 118666 42152
rect 125321 42143 125379 42149
rect 125321 42140 125333 42143
rect 118660 42112 125333 42140
rect 118660 42100 118666 42112
rect 125321 42109 125333 42112
rect 125367 42109 125379 42143
rect 125321 42103 125379 42109
rect 5442 42032 5448 42084
rect 5500 42072 5506 42084
rect 47854 42072 47860 42084
rect 5500 42044 47860 42072
rect 5500 42032 5506 42044
rect 47854 42032 47860 42044
rect 47912 42032 47918 42084
rect 49602 42032 49608 42084
rect 49660 42072 49666 42084
rect 59906 42072 59912 42084
rect 49660 42044 59912 42072
rect 49660 42032 49666 42044
rect 59906 42032 59912 42044
rect 59964 42032 59970 42084
rect 60001 42075 60059 42081
rect 60001 42041 60013 42075
rect 60047 42072 60059 42075
rect 85114 42072 85120 42084
rect 60047 42044 85120 42072
rect 60047 42041 60059 42044
rect 60001 42035 60059 42041
rect 85114 42032 85120 42044
rect 85172 42032 85178 42084
rect 85482 42032 85488 42084
rect 85540 42072 85546 42084
rect 113450 42072 113456 42084
rect 85540 42044 113456 42072
rect 85540 42032 85546 42044
rect 113450 42032 113456 42044
rect 113508 42032 113514 42084
rect 117222 42032 117228 42084
rect 117280 42072 117286 42084
rect 122469 42075 122527 42081
rect 122469 42072 122481 42075
rect 117280 42044 122481 42072
rect 117280 42032 117286 42044
rect 122469 42041 122481 42044
rect 122515 42041 122527 42075
rect 125520 42072 125548 42180
rect 125686 42168 125692 42220
rect 125744 42208 125750 42220
rect 146754 42208 146760 42220
rect 125744 42180 146760 42208
rect 125744 42168 125750 42180
rect 146754 42168 146760 42180
rect 146812 42168 146818 42220
rect 147582 42168 147588 42220
rect 147640 42208 147646 42220
rect 164418 42208 164424 42220
rect 147640 42180 164424 42208
rect 147640 42168 147646 42180
rect 164418 42168 164424 42180
rect 164476 42168 164482 42220
rect 168190 42168 168196 42220
rect 168248 42208 168254 42220
rect 182082 42208 182088 42220
rect 168248 42180 182088 42208
rect 168248 42168 168254 42180
rect 182082 42168 182088 42180
rect 182140 42168 182146 42220
rect 184750 42168 184756 42220
rect 184808 42208 184814 42220
rect 195790 42208 195796 42220
rect 184808 42180 195796 42208
rect 184808 42168 184814 42180
rect 195790 42168 195796 42180
rect 195848 42168 195854 42220
rect 195882 42168 195888 42220
rect 195940 42208 195946 42220
rect 204622 42208 204628 42220
rect 195940 42180 204628 42208
rect 195940 42168 195946 42180
rect 204622 42168 204628 42180
rect 204680 42168 204686 42220
rect 206922 42168 206928 42220
rect 206980 42208 206986 42220
rect 213362 42208 213368 42220
rect 206980 42180 213368 42208
rect 206980 42168 206986 42180
rect 213362 42168 213368 42180
rect 213420 42168 213426 42220
rect 213822 42168 213828 42220
rect 213880 42208 213886 42220
rect 219250 42208 219256 42220
rect 213880 42180 219256 42208
rect 213880 42168 213886 42180
rect 219250 42168 219256 42180
rect 219308 42168 219314 42220
rect 368198 42168 368204 42220
rect 368256 42208 368262 42220
rect 393498 42208 393504 42220
rect 368256 42180 393504 42208
rect 368256 42168 368262 42180
rect 393498 42168 393504 42180
rect 393556 42168 393562 42220
rect 407390 42168 407396 42220
rect 407448 42208 407454 42220
rect 408402 42208 408408 42220
rect 407448 42180 408408 42208
rect 407448 42168 407454 42180
rect 408402 42168 408408 42180
rect 408460 42168 408466 42220
rect 425974 42168 425980 42220
rect 426032 42208 426038 42220
rect 462958 42208 462964 42220
rect 426032 42180 462964 42208
rect 426032 42168 426038 42180
rect 462958 42168 462964 42180
rect 463016 42168 463022 42220
rect 477862 42168 477868 42220
rect 477920 42208 477926 42220
rect 527174 42208 527180 42220
rect 477920 42180 527180 42208
rect 477920 42168 477926 42180
rect 527174 42168 527180 42180
rect 527232 42168 527238 42220
rect 125597 42143 125655 42149
rect 125597 42109 125609 42143
rect 125643 42140 125655 42143
rect 140958 42140 140964 42152
rect 125643 42112 140964 42140
rect 125643 42109 125655 42112
rect 125597 42103 125655 42109
rect 140958 42100 140964 42112
rect 141016 42100 141022 42152
rect 143442 42100 143448 42152
rect 143500 42140 143506 42152
rect 161474 42140 161480 42152
rect 143500 42112 161480 42140
rect 143500 42100 143506 42112
rect 161474 42100 161480 42112
rect 161532 42100 161538 42152
rect 164142 42100 164148 42152
rect 164200 42140 164206 42152
rect 178126 42140 178132 42152
rect 164200 42112 178132 42140
rect 164200 42100 164206 42112
rect 178126 42100 178132 42112
rect 178184 42100 178190 42152
rect 179322 42100 179328 42152
rect 179380 42140 179386 42152
rect 190914 42140 190920 42152
rect 179380 42112 190920 42140
rect 179380 42100 179386 42112
rect 190914 42100 190920 42112
rect 190972 42100 190978 42152
rect 193122 42100 193128 42152
rect 193180 42140 193186 42152
rect 201678 42140 201684 42152
rect 193180 42112 201684 42140
rect 193180 42100 193186 42112
rect 201678 42100 201684 42112
rect 201736 42100 201742 42152
rect 202782 42100 202788 42152
rect 202840 42140 202846 42152
rect 210418 42140 210424 42152
rect 202840 42112 210424 42140
rect 202840 42100 202846 42112
rect 210418 42100 210424 42112
rect 210476 42100 210482 42152
rect 217962 42100 217968 42152
rect 218020 42140 218026 42152
rect 222194 42140 222200 42152
rect 218020 42112 222200 42140
rect 218020 42100 218026 42112
rect 222194 42100 222200 42112
rect 222252 42100 222258 42152
rect 344646 42100 344652 42152
rect 344704 42140 344710 42152
rect 365806 42140 365812 42152
rect 344704 42112 365812 42140
rect 344704 42100 344710 42112
rect 365806 42100 365812 42112
rect 365864 42100 365870 42152
rect 371142 42100 371148 42152
rect 371200 42140 371206 42152
rect 397638 42140 397644 42152
rect 371200 42112 397644 42140
rect 371200 42100 371206 42112
rect 397638 42100 397644 42112
rect 397696 42100 397702 42152
rect 400490 42100 400496 42152
rect 400548 42140 400554 42152
rect 433426 42140 433432 42152
rect 400548 42112 433432 42140
rect 400548 42100 400554 42112
rect 433426 42100 433432 42112
rect 433484 42100 433490 42152
rect 443546 42100 443552 42152
rect 443604 42140 443610 42152
rect 485774 42140 485780 42152
rect 443604 42112 485780 42140
rect 443604 42100 443610 42112
rect 485774 42100 485780 42112
rect 485832 42100 485838 42152
rect 490650 42100 490656 42152
rect 490708 42140 490714 42152
rect 540238 42140 540244 42152
rect 490708 42112 540244 42140
rect 490708 42100 490714 42112
rect 540238 42100 540244 42112
rect 540296 42100 540302 42152
rect 139946 42072 139952 42084
rect 125520 42044 139952 42072
rect 122469 42035 122527 42041
rect 139946 42032 139952 42044
rect 140004 42032 140010 42084
rect 142062 42032 142068 42084
rect 142120 42072 142126 42084
rect 160462 42072 160468 42084
rect 142120 42044 160468 42072
rect 142120 42032 142126 42044
rect 160462 42032 160468 42044
rect 160520 42032 160526 42084
rect 162762 42032 162768 42084
rect 162820 42072 162826 42084
rect 177114 42072 177120 42084
rect 162820 42044 177120 42072
rect 162820 42032 162826 42044
rect 177114 42032 177120 42044
rect 177172 42032 177178 42084
rect 177942 42032 177948 42084
rect 178000 42072 178006 42084
rect 189902 42072 189908 42084
rect 178000 42044 189908 42072
rect 178000 42032 178006 42044
rect 189902 42032 189908 42044
rect 189960 42032 189966 42084
rect 194410 42032 194416 42084
rect 194468 42072 194474 42084
rect 203610 42072 203616 42084
rect 194468 42044 203616 42072
rect 194468 42032 194474 42044
rect 203610 42032 203616 42044
rect 203668 42032 203674 42084
rect 219250 42032 219256 42084
rect 219308 42072 219314 42084
rect 224218 42072 224224 42084
rect 219308 42044 224224 42072
rect 219308 42032 219314 42044
rect 224218 42032 224224 42044
rect 224276 42032 224282 42084
rect 229002 42032 229008 42084
rect 229060 42072 229066 42084
rect 232038 42072 232044 42084
rect 229060 42044 232044 42072
rect 229060 42032 229066 42044
rect 232038 42032 232044 42044
rect 232096 42032 232102 42084
rect 350534 42032 350540 42084
rect 350592 42072 350598 42084
rect 372706 42072 372712 42084
rect 350592 42044 372712 42072
rect 350592 42032 350598 42044
rect 372706 42032 372712 42044
rect 372764 42032 372770 42084
rect 376938 42032 376944 42084
rect 376996 42072 377002 42084
rect 404538 42072 404544 42084
rect 376996 42044 404544 42072
rect 376996 42032 377002 42044
rect 404538 42032 404544 42044
rect 404596 42032 404602 42084
rect 408310 42032 408316 42084
rect 408368 42072 408374 42084
rect 442994 42072 443000 42084
rect 408368 42044 443000 42072
rect 408368 42032 408374 42044
rect 442994 42032 443000 42044
rect 443052 42032 443058 42084
rect 445570 42032 445576 42084
rect 445628 42072 445634 42084
rect 483750 42072 483756 42084
rect 445628 42044 483756 42072
rect 445628 42032 445634 42044
rect 483750 42032 483756 42044
rect 483808 42032 483814 42084
rect 484762 42032 484768 42084
rect 484820 42072 484826 42084
rect 535454 42072 535460 42084
rect 484820 42044 535460 42072
rect 484820 42032 484826 42044
rect 535454 42032 535460 42044
rect 535512 42032 535518 42084
rect 31662 41964 31668 42016
rect 31720 42004 31726 42016
rect 67545 42007 67603 42013
rect 67545 42004 67557 42007
rect 31720 41976 67557 42004
rect 31720 41964 31726 41976
rect 67545 41973 67557 41976
rect 67591 41973 67603 42007
rect 67545 41967 67603 41973
rect 68189 42007 68247 42013
rect 68189 41973 68201 42007
rect 68235 42004 68247 42007
rect 75365 42007 75423 42013
rect 75365 42004 75377 42007
rect 68235 41976 75377 42004
rect 68235 41973 68247 41976
rect 68189 41967 68247 41973
rect 75365 41973 75377 41976
rect 75411 41973 75423 42007
rect 75365 41967 75423 41973
rect 75822 41964 75828 42016
rect 75880 42004 75886 42016
rect 105630 42004 105636 42016
rect 75880 41976 105636 42004
rect 75880 41964 75886 41976
rect 105630 41964 105636 41976
rect 105688 41964 105694 42016
rect 108945 42007 109003 42013
rect 108945 41973 108957 42007
rect 108991 42004 109003 42007
rect 133046 42004 133052 42016
rect 108991 41976 133052 42004
rect 108991 41973 109003 41976
rect 108945 41967 109003 41973
rect 133046 41964 133052 41976
rect 133104 41964 133110 42016
rect 133690 41964 133696 42016
rect 133748 42004 133754 42016
rect 152642 42004 152648 42016
rect 133748 41976 152648 42004
rect 133748 41964 133754 41976
rect 152642 41964 152648 41976
rect 152700 41964 152706 42016
rect 153102 41964 153108 42016
rect 153160 42004 153166 42016
rect 169294 42004 169300 42016
rect 153160 41976 169300 42004
rect 153160 41964 153166 41976
rect 169294 41964 169300 41976
rect 169352 41964 169358 42016
rect 176562 41964 176568 42016
rect 176620 42004 176626 42016
rect 188890 42004 188896 42016
rect 176620 41976 188896 42004
rect 176620 41964 176626 41976
rect 188890 41964 188896 41976
rect 188948 41964 188954 42016
rect 394602 41964 394608 42016
rect 394660 42004 394666 42016
rect 425238 42004 425244 42016
rect 394660 41976 425244 42004
rect 394660 41964 394666 41976
rect 425238 41964 425244 41976
rect 425296 41964 425302 42016
rect 464154 41964 464160 42016
rect 464212 42004 464218 42016
rect 508498 42004 508504 42016
rect 464212 41976 508504 42004
rect 464212 41964 464218 41976
rect 508498 41964 508504 41976
rect 508556 41964 508562 42016
rect 519998 41964 520004 42016
rect 520056 42004 520062 42016
rect 547138 42004 547144 42016
rect 520056 41976 547144 42004
rect 520056 41964 520062 41976
rect 547138 41964 547144 41976
rect 547196 41964 547202 42016
rect 28902 41896 28908 41948
rect 28960 41936 28966 41948
rect 59817 41939 59875 41945
rect 59817 41936 59829 41939
rect 28960 41908 59829 41936
rect 28960 41896 28966 41908
rect 59817 41905 59829 41908
rect 59863 41905 59875 41939
rect 59817 41899 59875 41905
rect 59906 41896 59912 41948
rect 59964 41936 59970 41948
rect 64601 41939 64659 41945
rect 64601 41936 64613 41939
rect 59964 41908 64613 41936
rect 59964 41896 59970 41908
rect 64601 41905 64613 41908
rect 64647 41905 64659 41939
rect 64601 41899 64659 41905
rect 69477 41939 69535 41945
rect 69477 41905 69489 41939
rect 69523 41936 69535 41939
rect 96798 41936 96804 41948
rect 69523 41908 96804 41936
rect 69523 41905 69535 41908
rect 69477 41899 69535 41905
rect 96798 41896 96804 41908
rect 96856 41896 96862 41948
rect 104802 41896 104808 41948
rect 104860 41936 104866 41948
rect 129182 41936 129188 41948
rect 104860 41908 129188 41936
rect 104860 41896 104866 41908
rect 129182 41896 129188 41908
rect 129240 41896 129246 41948
rect 131022 41896 131028 41948
rect 131080 41936 131086 41948
rect 150710 41936 150716 41948
rect 131080 41908 150716 41936
rect 131080 41896 131086 41908
rect 150710 41896 150716 41908
rect 150768 41896 150774 41948
rect 160002 41896 160008 41948
rect 160060 41936 160066 41948
rect 174814 41936 174820 41948
rect 160060 41908 174820 41936
rect 160060 41896 160066 41908
rect 174814 41896 174820 41908
rect 174872 41896 174878 41948
rect 184842 41896 184848 41948
rect 184900 41936 184906 41948
rect 194778 41936 194784 41948
rect 184900 41908 194784 41936
rect 184900 41896 184906 41908
rect 194778 41896 194784 41908
rect 194836 41896 194842 41948
rect 458266 41896 458272 41948
rect 458324 41936 458330 41948
rect 502426 41936 502432 41948
rect 458324 41908 502432 41936
rect 458324 41896 458330 41908
rect 502426 41896 502432 41908
rect 502484 41896 502490 41948
rect 507302 41896 507308 41948
rect 507360 41936 507366 41948
rect 537478 41936 537484 41948
rect 507360 41908 537484 41936
rect 507360 41896 507366 41908
rect 537478 41896 537484 41908
rect 537536 41896 537542 41948
rect 38470 41828 38476 41880
rect 38528 41868 38534 41880
rect 75270 41868 75276 41880
rect 38528 41840 75276 41868
rect 38528 41828 38534 41840
rect 75270 41828 75276 41840
rect 75328 41828 75334 41880
rect 75365 41871 75423 41877
rect 75365 41837 75377 41871
rect 75411 41868 75423 41871
rect 77202 41868 77208 41880
rect 75411 41840 77208 41868
rect 75411 41837 75423 41840
rect 75365 41831 75423 41837
rect 77202 41828 77208 41840
rect 77260 41828 77266 41880
rect 78582 41828 78588 41880
rect 78640 41868 78646 41880
rect 107654 41868 107660 41880
rect 78640 41840 107660 41868
rect 78640 41828 78646 41840
rect 107654 41828 107660 41840
rect 107712 41828 107718 41880
rect 110322 41828 110328 41880
rect 110380 41868 110386 41880
rect 123849 41871 123907 41877
rect 123849 41868 123861 41871
rect 110380 41840 123861 41868
rect 110380 41828 110386 41840
rect 123849 41837 123861 41840
rect 123895 41837 123907 41871
rect 123849 41831 123907 41837
rect 123941 41871 123999 41877
rect 123941 41837 123953 41871
rect 123987 41868 123999 41871
rect 127526 41868 127532 41880
rect 123987 41840 127532 41868
rect 123987 41837 123999 41840
rect 123941 41831 123999 41837
rect 127526 41828 127532 41840
rect 127584 41828 127590 41880
rect 127621 41871 127679 41877
rect 127621 41837 127633 41871
rect 127667 41868 127679 41871
rect 135070 41868 135076 41880
rect 127667 41840 135076 41868
rect 127667 41837 127679 41840
rect 127621 41831 127679 41837
rect 135070 41828 135076 41840
rect 135128 41828 135134 41880
rect 135162 41828 135168 41880
rect 135220 41868 135226 41880
rect 136177 41871 136235 41877
rect 136177 41868 136189 41871
rect 135220 41840 136189 41868
rect 135220 41828 135226 41840
rect 136177 41837 136189 41840
rect 136223 41837 136235 41871
rect 136177 41831 136235 41837
rect 137922 41828 137928 41880
rect 137980 41868 137986 41880
rect 156598 41868 156604 41880
rect 137980 41840 156604 41868
rect 137980 41828 137986 41840
rect 156598 41828 156604 41840
rect 156656 41828 156662 41880
rect 157242 41828 157248 41880
rect 157300 41868 157306 41880
rect 172238 41868 172244 41880
rect 157300 41840 172244 41868
rect 157300 41828 157306 41840
rect 172238 41828 172244 41840
rect 172296 41828 172302 41880
rect 446490 41828 446496 41880
rect 446548 41868 446554 41880
rect 486418 41868 486424 41880
rect 446548 41840 486424 41868
rect 446548 41828 446554 41840
rect 486418 41828 486424 41840
rect 486476 41828 486482 41880
rect 495526 41828 495532 41880
rect 495584 41868 495590 41880
rect 533338 41868 533344 41880
rect 495584 41840 533344 41868
rect 495584 41828 495590 41840
rect 533338 41828 533344 41840
rect 533396 41828 533402 41880
rect 35802 41760 35808 41812
rect 35860 41800 35866 41812
rect 66809 41803 66867 41809
rect 66809 41800 66821 41803
rect 35860 41772 66821 41800
rect 35860 41760 35866 41772
rect 66809 41769 66821 41772
rect 66855 41769 66867 41803
rect 66809 41763 66867 41769
rect 66898 41760 66904 41812
rect 66956 41800 66962 41812
rect 69477 41803 69535 41809
rect 69477 41800 69489 41803
rect 66956 41772 69489 41800
rect 66956 41760 66962 41772
rect 69477 41769 69489 41772
rect 69523 41769 69535 41803
rect 69477 41763 69535 41769
rect 69569 41803 69627 41809
rect 69569 41769 69581 41803
rect 69615 41800 69627 41803
rect 74353 41803 74411 41809
rect 74353 41800 74365 41803
rect 69615 41772 74365 41800
rect 69615 41769 69627 41772
rect 69569 41763 69627 41769
rect 74353 41769 74365 41772
rect 74399 41769 74411 41803
rect 74353 41763 74411 41769
rect 74442 41760 74448 41812
rect 74500 41800 74506 41812
rect 104710 41800 104716 41812
rect 74500 41772 104716 41800
rect 74500 41760 74506 41772
rect 104710 41760 104716 41772
rect 104768 41760 104774 41812
rect 106182 41760 106188 41812
rect 106240 41800 106246 41812
rect 113177 41803 113235 41809
rect 113177 41800 113189 41803
rect 106240 41772 113189 41800
rect 106240 41760 106246 41772
rect 113177 41769 113189 41772
rect 113223 41769 113235 41803
rect 113177 41763 113235 41769
rect 122745 41803 122803 41809
rect 122745 41769 122757 41803
rect 122791 41800 122803 41803
rect 124033 41803 124091 41809
rect 124033 41800 124045 41803
rect 122791 41772 124045 41800
rect 122791 41769 122803 41772
rect 122745 41763 122803 41769
rect 124033 41769 124045 41772
rect 124079 41769 124091 41803
rect 124033 41763 124091 41769
rect 124122 41760 124128 41812
rect 124180 41800 124186 41812
rect 144822 41800 144828 41812
rect 124180 41772 144828 41800
rect 124180 41760 124186 41772
rect 144822 41760 144828 41772
rect 144880 41760 144886 41812
rect 148962 41760 148968 41812
rect 149020 41800 149026 41812
rect 165430 41800 165436 41812
rect 149020 41772 165436 41800
rect 149020 41760 149026 41772
rect 165430 41760 165436 41772
rect 165488 41760 165494 41812
rect 166902 41760 166908 41812
rect 166960 41800 166966 41812
rect 180058 41800 180064 41812
rect 166960 41772 180064 41800
rect 166960 41760 166966 41772
rect 180058 41760 180064 41772
rect 180116 41760 180122 41812
rect 463142 41760 463148 41812
rect 463200 41800 463206 41812
rect 501598 41800 501604 41812
rect 463200 41772 501604 41800
rect 463200 41760 463206 41772
rect 501598 41760 501604 41772
rect 501656 41760 501662 41812
rect 513098 41760 513104 41812
rect 513156 41800 513162 41812
rect 537570 41800 537576 41812
rect 513156 41772 537576 41800
rect 513156 41760 513162 41772
rect 537570 41760 537576 41772
rect 537628 41760 537634 41812
rect 42702 41692 42708 41744
rect 42760 41732 42766 41744
rect 78214 41732 78220 41744
rect 42760 41704 78220 41732
rect 42760 41692 42766 41704
rect 78214 41692 78220 41704
rect 78272 41692 78278 41744
rect 79962 41692 79968 41744
rect 80020 41732 80026 41744
rect 108574 41732 108580 41744
rect 80020 41704 108580 41732
rect 80020 41692 80026 41704
rect 108574 41692 108580 41704
rect 108632 41692 108638 41744
rect 115842 41692 115848 41744
rect 115900 41732 115906 41744
rect 138014 41732 138020 41744
rect 115900 41704 138020 41732
rect 115900 41692 115906 41704
rect 138014 41692 138020 41704
rect 138072 41692 138078 41744
rect 140682 41692 140688 41744
rect 140740 41732 140746 41744
rect 158530 41732 158536 41744
rect 140740 41704 158536 41732
rect 140740 41692 140746 41704
rect 158530 41692 158536 41704
rect 158588 41692 158594 41744
rect 161382 41692 161388 41744
rect 161440 41732 161446 41744
rect 176194 41732 176200 41744
rect 161440 41704 176200 41732
rect 161440 41692 161446 41704
rect 176194 41692 176200 41704
rect 176252 41692 176258 41744
rect 211062 41692 211068 41744
rect 211120 41732 211126 41744
rect 217318 41732 217324 41744
rect 211120 41704 217324 41732
rect 211120 41692 211126 41704
rect 217318 41692 217324 41704
rect 217376 41692 217382 41744
rect 434806 41692 434812 41744
rect 434864 41732 434870 41744
rect 467098 41732 467104 41744
rect 434864 41704 467104 41732
rect 434864 41692 434870 41704
rect 467098 41692 467104 41704
rect 467156 41692 467162 41744
rect 475930 41692 475936 41744
rect 475988 41732 475994 41744
rect 496078 41732 496084 41744
rect 475988 41704 496084 41732
rect 475988 41692 475994 41704
rect 496078 41692 496084 41704
rect 496136 41692 496142 41744
rect 501414 41692 501420 41744
rect 501472 41732 501478 41744
rect 534718 41732 534724 41744
rect 501472 41704 534724 41732
rect 501472 41692 501478 41704
rect 534718 41692 534724 41704
rect 534776 41692 534782 41744
rect 45462 41624 45468 41676
rect 45520 41664 45526 41676
rect 80146 41664 80152 41676
rect 45520 41636 80152 41664
rect 45520 41624 45526 41636
rect 80146 41624 80152 41636
rect 80204 41624 80210 41676
rect 80241 41667 80299 41673
rect 80241 41633 80253 41667
rect 80287 41664 80299 41667
rect 83366 41664 83372 41676
rect 80287 41636 83372 41664
rect 80287 41633 80299 41636
rect 80241 41627 80299 41633
rect 83366 41624 83372 41636
rect 83424 41624 83430 41676
rect 83458 41624 83464 41676
rect 83516 41664 83522 41676
rect 111518 41664 111524 41676
rect 83516 41636 111524 41664
rect 83516 41624 83522 41636
rect 111518 41624 111524 41636
rect 111576 41624 111582 41676
rect 111702 41624 111708 41676
rect 111760 41664 111766 41676
rect 127621 41667 127679 41673
rect 127621 41664 127633 41667
rect 111760 41636 127633 41664
rect 111760 41624 111766 41636
rect 127621 41633 127633 41636
rect 127667 41633 127679 41667
rect 130102 41664 130108 41676
rect 127621 41627 127679 41633
rect 127728 41636 130108 41664
rect 41322 41556 41328 41608
rect 41380 41596 41386 41608
rect 68189 41599 68247 41605
rect 68189 41596 68201 41599
rect 41380 41568 68201 41596
rect 41380 41556 41386 41568
rect 68189 41565 68201 41568
rect 68235 41565 68247 41599
rect 68189 41559 68247 41565
rect 68278 41556 68284 41608
rect 68336 41596 68342 41608
rect 73338 41596 73344 41608
rect 68336 41568 73344 41596
rect 68336 41556 68342 41568
rect 73338 41556 73344 41568
rect 73396 41556 73402 41608
rect 73798 41556 73804 41608
rect 73856 41596 73862 41608
rect 102686 41596 102692 41608
rect 73856 41568 102692 41596
rect 73856 41556 73862 41568
rect 102686 41556 102692 41568
rect 102744 41556 102750 41608
rect 103422 41556 103428 41608
rect 103480 41596 103486 41608
rect 123941 41599 123999 41605
rect 123941 41596 123953 41599
rect 103480 41568 123953 41596
rect 103480 41556 103486 41568
rect 123941 41565 123953 41568
rect 123987 41565 123999 41599
rect 123941 41559 123999 41565
rect 124033 41599 124091 41605
rect 124033 41565 124045 41599
rect 124079 41596 124091 41599
rect 127728 41596 127756 41636
rect 130102 41624 130108 41636
rect 130160 41624 130166 41676
rect 132402 41624 132408 41676
rect 132460 41664 132466 41676
rect 151446 41664 151452 41676
rect 132460 41636 151452 41664
rect 132460 41624 132466 41636
rect 151446 41624 151452 41636
rect 151504 41624 151510 41676
rect 201402 41624 201408 41676
rect 201460 41664 201466 41676
rect 208486 41664 208492 41676
rect 201460 41636 208492 41664
rect 201460 41624 201466 41636
rect 208486 41624 208492 41636
rect 208544 41624 208550 41676
rect 212534 41624 212540 41676
rect 212592 41664 212598 41676
rect 218330 41664 218336 41676
rect 212592 41636 218336 41664
rect 212592 41624 212598 41636
rect 218330 41624 218336 41636
rect 218388 41624 218394 41676
rect 220722 41624 220728 41676
rect 220780 41664 220786 41676
rect 225138 41664 225144 41676
rect 220780 41636 225144 41664
rect 220780 41624 220786 41636
rect 225138 41624 225144 41636
rect 225196 41624 225202 41676
rect 440694 41624 440700 41676
rect 440752 41664 440758 41676
rect 468478 41664 468484 41676
rect 440752 41636 468484 41664
rect 440752 41624 440758 41636
rect 468478 41624 468484 41636
rect 468536 41624 468542 41676
rect 518986 41624 518992 41676
rect 519044 41664 519050 41676
rect 538858 41664 538864 41676
rect 519044 41636 538864 41664
rect 519044 41624 519050 41636
rect 538858 41624 538864 41636
rect 538916 41624 538922 41676
rect 124079 41568 127756 41596
rect 124079 41565 124091 41568
rect 124033 41559 124091 41565
rect 128262 41556 128268 41608
rect 128320 41596 128326 41608
rect 148778 41596 148784 41608
rect 128320 41568 148784 41596
rect 128320 41556 128326 41568
rect 148778 41556 148784 41568
rect 148836 41556 148842 41608
rect 150342 41556 150348 41608
rect 150400 41596 150406 41608
rect 166350 41596 166356 41608
rect 150400 41568 166356 41596
rect 150400 41556 150406 41568
rect 166350 41556 166356 41568
rect 166408 41556 166414 41608
rect 202690 41556 202696 41608
rect 202748 41596 202754 41608
rect 209498 41596 209504 41608
rect 202748 41568 209504 41596
rect 202748 41556 202754 41568
rect 209498 41556 209504 41568
rect 209556 41556 209562 41608
rect 210970 41556 210976 41608
rect 211028 41596 211034 41608
rect 216306 41596 216312 41608
rect 211028 41568 216312 41596
rect 211028 41556 211034 41568
rect 216306 41556 216312 41568
rect 216364 41556 216370 41608
rect 224862 41556 224868 41608
rect 224920 41596 224926 41608
rect 228082 41596 228088 41608
rect 224920 41568 228088 41596
rect 224920 41556 224926 41568
rect 228082 41556 228088 41568
rect 228140 41556 228146 41608
rect 521010 41556 521016 41608
rect 521068 41596 521074 41608
rect 529198 41596 529204 41608
rect 521068 41568 529204 41596
rect 521068 41556 521074 41568
rect 529198 41556 529204 41568
rect 529256 41556 529262 41608
rect 46198 41488 46204 41540
rect 46256 41528 46262 41540
rect 48866 41528 48872 41540
rect 46256 41500 48872 41528
rect 46256 41488 46262 41500
rect 48866 41488 48872 41500
rect 48924 41488 48930 41540
rect 50338 41488 50344 41540
rect 50396 41528 50402 41540
rect 55674 41528 55680 41540
rect 50396 41500 55680 41528
rect 50396 41488 50402 41500
rect 55674 41488 55680 41500
rect 55732 41488 55738 41540
rect 57238 41488 57244 41540
rect 57296 41528 57302 41540
rect 64506 41528 64512 41540
rect 57296 41500 64512 41528
rect 57296 41488 57302 41500
rect 64506 41488 64512 41500
rect 64564 41488 64570 41540
rect 64601 41531 64659 41537
rect 64601 41497 64613 41531
rect 64647 41528 64659 41531
rect 80241 41531 80299 41537
rect 80241 41528 80253 41531
rect 64647 41500 80253 41528
rect 64647 41497 64659 41500
rect 64601 41491 64659 41497
rect 80241 41497 80253 41500
rect 80287 41497 80299 41531
rect 80241 41491 80299 41497
rect 80698 41488 80704 41540
rect 80756 41528 80762 41540
rect 82170 41528 82176 41540
rect 80756 41500 82176 41528
rect 80756 41488 80762 41500
rect 82170 41488 82176 41500
rect 82228 41488 82234 41540
rect 86862 41488 86868 41540
rect 86920 41528 86926 41540
rect 114094 41528 114100 41540
rect 86920 41500 114100 41528
rect 86920 41488 86926 41500
rect 114094 41488 114100 41500
rect 114152 41488 114158 41540
rect 114462 41488 114468 41540
rect 114520 41528 114526 41540
rect 137002 41528 137008 41540
rect 114520 41500 137008 41528
rect 114520 41488 114526 41500
rect 137002 41488 137008 41500
rect 137060 41488 137066 41540
rect 204162 41488 204168 41540
rect 204220 41528 204226 41540
rect 211430 41528 211436 41540
rect 204220 41500 211436 41528
rect 204220 41488 204226 41500
rect 211430 41488 211436 41500
rect 211488 41488 211494 41540
rect 215202 41488 215208 41540
rect 215260 41528 215266 41540
rect 220262 41528 220268 41540
rect 215260 41500 220268 41528
rect 215260 41488 215266 41500
rect 220262 41488 220268 41500
rect 220320 41488 220326 41540
rect 222102 41488 222108 41540
rect 222160 41528 222166 41540
rect 226150 41528 226156 41540
rect 222160 41500 226156 41528
rect 222160 41488 222166 41500
rect 226150 41488 226156 41500
rect 226208 41488 226214 41540
rect 226242 41488 226248 41540
rect 226300 41528 226306 41540
rect 229094 41528 229100 41540
rect 226300 41500 229100 41528
rect 226300 41488 226306 41500
rect 229094 41488 229100 41500
rect 229152 41488 229158 41540
rect 230382 41488 230388 41540
rect 230440 41528 230446 41540
rect 232958 41528 232964 41540
rect 230440 41500 232964 41528
rect 230440 41488 230446 41500
rect 232958 41488 232964 41500
rect 233016 41488 233022 41540
rect 233142 41488 233148 41540
rect 233200 41528 233206 41540
rect 234982 41528 234988 41540
rect 233200 41500 234988 41528
rect 233200 41488 233206 41500
rect 234982 41488 234988 41500
rect 235040 41488 235046 41540
rect 257522 41488 257528 41540
rect 257580 41528 257586 41540
rect 258718 41528 258724 41540
rect 257580 41500 258724 41528
rect 257580 41488 257586 41500
rect 258718 41488 258724 41500
rect 258776 41488 258782 41540
rect 264330 41488 264336 41540
rect 264388 41528 264394 41540
rect 266998 41528 267004 41540
rect 264388 41500 267004 41528
rect 264388 41488 264394 41500
rect 266998 41488 267004 41500
rect 267056 41488 267062 41540
rect 271230 41488 271236 41540
rect 271288 41528 271294 41540
rect 272518 41528 272524 41540
rect 271288 41500 272524 41528
rect 271288 41488 271294 41500
rect 272518 41488 272524 41500
rect 272576 41488 272582 41540
rect 396534 41488 396540 41540
rect 396592 41528 396598 41540
rect 396592 41500 399432 41528
rect 396592 41488 396598 41500
rect 39298 41420 39304 41472
rect 39356 41460 39362 41472
rect 59909 41463 59967 41469
rect 59909 41460 59921 41463
rect 39356 41432 59921 41460
rect 39356 41420 39362 41432
rect 59909 41429 59921 41432
rect 59955 41429 59967 41463
rect 59909 41423 59967 41429
rect 59998 41420 60004 41472
rect 60056 41460 60062 41472
rect 63494 41460 63500 41472
rect 60056 41432 63500 41460
rect 60056 41420 60062 41432
rect 63494 41420 63500 41432
rect 63552 41420 63558 41472
rect 67542 41420 67548 41472
rect 67600 41460 67606 41472
rect 69569 41463 69627 41469
rect 69569 41460 69581 41463
rect 67600 41432 69581 41460
rect 67600 41420 67606 41432
rect 69569 41429 69581 41432
rect 69615 41429 69627 41463
rect 69569 41423 69627 41429
rect 71682 41420 71688 41472
rect 71740 41460 71746 41472
rect 101766 41460 101772 41472
rect 71740 41432 101772 41460
rect 71740 41420 71746 41432
rect 101766 41420 101772 41432
rect 101824 41420 101830 41472
rect 113082 41420 113088 41472
rect 113140 41460 113146 41472
rect 135990 41460 135996 41472
rect 113140 41432 135996 41460
rect 113140 41420 113146 41432
rect 135990 41420 135996 41432
rect 136048 41420 136054 41472
rect 136542 41420 136548 41472
rect 136600 41460 136606 41472
rect 155586 41460 155592 41472
rect 136600 41432 155592 41460
rect 136600 41420 136606 41432
rect 155586 41420 155592 41432
rect 155644 41420 155650 41472
rect 194502 41420 194508 41472
rect 194560 41460 194566 41472
rect 202598 41460 202604 41472
rect 194560 41432 202604 41460
rect 194560 41420 194566 41432
rect 202598 41420 202604 41432
rect 202656 41420 202662 41472
rect 205542 41420 205548 41472
rect 205600 41460 205606 41472
rect 212442 41460 212448 41472
rect 205600 41432 212448 41460
rect 205600 41420 205606 41432
rect 212442 41420 212448 41432
rect 212500 41420 212506 41472
rect 216582 41420 216588 41472
rect 216640 41460 216646 41472
rect 221274 41460 221280 41472
rect 216640 41432 221280 41460
rect 216640 41420 216646 41432
rect 221274 41420 221280 41432
rect 221332 41420 221338 41472
rect 223482 41420 223488 41472
rect 223540 41460 223546 41472
rect 227070 41460 227076 41472
rect 223540 41432 227076 41460
rect 223540 41420 223546 41432
rect 227070 41420 227076 41432
rect 227128 41420 227134 41472
rect 227622 41420 227628 41472
rect 227680 41460 227686 41472
rect 230014 41460 230020 41472
rect 227680 41432 230020 41460
rect 227680 41420 227686 41432
rect 230014 41420 230020 41432
rect 230072 41420 230078 41472
rect 231762 41420 231768 41472
rect 231820 41460 231826 41472
rect 233970 41460 233976 41472
rect 231820 41432 233976 41460
rect 231820 41420 231826 41432
rect 233970 41420 233976 41432
rect 234028 41420 234034 41472
rect 234522 41420 234528 41472
rect 234580 41460 234586 41472
rect 235902 41460 235908 41472
rect 234580 41432 235908 41460
rect 234580 41420 234586 41432
rect 235902 41420 235908 41432
rect 235960 41420 235966 41472
rect 255498 41420 255504 41472
rect 255556 41460 255562 41472
rect 256694 41460 256700 41472
rect 255556 41432 256700 41460
rect 255556 41420 255562 41432
rect 256694 41420 256700 41432
rect 256752 41420 256758 41472
rect 258442 41420 258448 41472
rect 258500 41460 258506 41472
rect 259362 41460 259368 41472
rect 258500 41432 259368 41460
rect 258500 41420 258506 41432
rect 259362 41420 259368 41432
rect 259420 41420 259426 41472
rect 259454 41420 259460 41472
rect 259512 41460 259518 41472
rect 261478 41460 261484 41472
rect 259512 41432 261484 41460
rect 259512 41420 259518 41432
rect 261478 41420 261484 41432
rect 261536 41420 261542 41472
rect 262398 41420 262404 41472
rect 262456 41460 262462 41472
rect 263410 41460 263416 41472
rect 262456 41432 263416 41460
rect 262456 41420 262462 41432
rect 263410 41420 263416 41432
rect 263468 41420 263474 41472
rect 265342 41420 265348 41472
rect 265400 41460 265406 41472
rect 266170 41460 266176 41472
rect 265400 41432 266176 41460
rect 265400 41420 265406 41432
rect 266170 41420 266176 41432
rect 266228 41420 266234 41472
rect 268286 41420 268292 41472
rect 268344 41460 268350 41472
rect 269022 41460 269028 41472
rect 268344 41432 269028 41460
rect 268344 41420 268350 41432
rect 269022 41420 269028 41432
rect 269080 41420 269086 41472
rect 269206 41420 269212 41472
rect 269264 41460 269270 41472
rect 270402 41460 270408 41472
rect 269264 41432 270408 41460
rect 269264 41420 269270 41432
rect 270402 41420 270408 41432
rect 270460 41420 270466 41472
rect 272150 41420 272156 41472
rect 272208 41460 272214 41472
rect 273070 41460 273076 41472
rect 272208 41432 273076 41460
rect 272208 41420 272214 41432
rect 273070 41420 273076 41432
rect 273128 41420 273134 41472
rect 275094 41420 275100 41472
rect 275152 41460 275158 41472
rect 275922 41460 275928 41472
rect 275152 41432 275928 41460
rect 275152 41420 275158 41432
rect 275922 41420 275928 41432
rect 275980 41420 275986 41472
rect 276106 41420 276112 41472
rect 276164 41460 276170 41472
rect 277302 41460 277308 41472
rect 276164 41432 277308 41460
rect 276164 41420 276170 41432
rect 277302 41420 277308 41432
rect 277360 41420 277366 41472
rect 279050 41420 279056 41472
rect 279108 41460 279114 41472
rect 280062 41460 280068 41472
rect 279108 41432 280068 41460
rect 279108 41420 279114 41432
rect 280062 41420 280068 41432
rect 280120 41420 280126 41472
rect 281994 41420 282000 41472
rect 282052 41460 282058 41472
rect 282822 41460 282828 41472
rect 282052 41432 282828 41460
rect 282052 41420 282058 41432
rect 282822 41420 282828 41432
rect 282880 41420 282886 41472
rect 282914 41420 282920 41472
rect 282972 41460 282978 41472
rect 284110 41460 284116 41472
rect 282972 41432 284116 41460
rect 282972 41420 282978 41432
rect 284110 41420 284116 41432
rect 284168 41420 284174 41472
rect 285858 41420 285864 41472
rect 285916 41460 285922 41472
rect 286870 41460 286876 41472
rect 285916 41432 286876 41460
rect 285916 41420 285922 41432
rect 286870 41420 286876 41432
rect 286928 41420 286934 41472
rect 288802 41420 288808 41472
rect 288860 41460 288866 41472
rect 289722 41460 289728 41472
rect 288860 41432 289728 41460
rect 288860 41420 288866 41432
rect 289722 41420 289728 41432
rect 289780 41420 289786 41472
rect 289814 41420 289820 41472
rect 289872 41460 289878 41472
rect 291102 41460 291108 41472
rect 289872 41432 291108 41460
rect 289872 41420 289878 41432
rect 291102 41420 291108 41432
rect 291160 41420 291166 41472
rect 292758 41420 292764 41472
rect 292816 41460 292822 41472
rect 293770 41460 293776 41472
rect 292816 41432 293776 41460
rect 292816 41420 292822 41432
rect 293770 41420 293776 41432
rect 293828 41420 293834 41472
rect 295702 41420 295708 41472
rect 295760 41460 295766 41472
rect 296530 41460 296536 41472
rect 295760 41432 296536 41460
rect 295760 41420 295766 41432
rect 296530 41420 296536 41432
rect 296588 41420 296594 41472
rect 298646 41420 298652 41472
rect 298704 41460 298710 41472
rect 299382 41460 299388 41472
rect 298704 41432 299388 41460
rect 298704 41420 298710 41432
rect 299382 41420 299388 41432
rect 299440 41420 299446 41472
rect 299566 41420 299572 41472
rect 299624 41460 299630 41472
rect 300762 41460 300768 41472
rect 299624 41432 300768 41460
rect 299624 41420 299630 41432
rect 300762 41420 300768 41432
rect 300820 41420 300826 41472
rect 302510 41420 302516 41472
rect 302568 41460 302574 41472
rect 303522 41460 303528 41472
rect 302568 41432 303528 41460
rect 302568 41420 302574 41432
rect 303522 41420 303528 41432
rect 303580 41420 303586 41472
rect 305454 41420 305460 41472
rect 305512 41460 305518 41472
rect 306282 41460 306288 41472
rect 305512 41432 306288 41460
rect 305512 41420 305518 41432
rect 306282 41420 306288 41432
rect 306340 41420 306346 41472
rect 306466 41420 306472 41472
rect 306524 41460 306530 41472
rect 307570 41460 307576 41472
rect 306524 41432 307576 41460
rect 306524 41420 306530 41432
rect 307570 41420 307576 41432
rect 307628 41420 307634 41472
rect 309410 41420 309416 41472
rect 309468 41460 309474 41472
rect 310330 41460 310336 41472
rect 309468 41432 310336 41460
rect 309468 41420 309474 41432
rect 310330 41420 310336 41432
rect 310388 41420 310394 41472
rect 312354 41420 312360 41472
rect 312412 41460 312418 41472
rect 313182 41460 313188 41472
rect 312412 41432 313188 41460
rect 312412 41420 312418 41432
rect 313182 41420 313188 41432
rect 313240 41420 313246 41472
rect 313274 41420 313280 41472
rect 313332 41460 313338 41472
rect 314562 41460 314568 41472
rect 313332 41432 314568 41460
rect 313332 41420 313338 41432
rect 314562 41420 314568 41432
rect 314620 41420 314626 41472
rect 316218 41420 316224 41472
rect 316276 41460 316282 41472
rect 317230 41460 317236 41472
rect 316276 41432 317236 41460
rect 316276 41420 316282 41432
rect 317230 41420 317236 41432
rect 317288 41420 317294 41472
rect 319162 41420 319168 41472
rect 319220 41460 319226 41472
rect 320082 41460 320088 41472
rect 319220 41432 320088 41460
rect 319220 41420 319226 41432
rect 320082 41420 320088 41432
rect 320140 41420 320146 41472
rect 320174 41420 320180 41472
rect 320232 41460 320238 41472
rect 321462 41460 321468 41472
rect 320232 41432 321468 41460
rect 320232 41420 320238 41432
rect 321462 41420 321468 41432
rect 321520 41420 321526 41472
rect 323118 41420 323124 41472
rect 323176 41460 323182 41472
rect 324222 41460 324228 41472
rect 323176 41432 324228 41460
rect 323176 41420 323182 41432
rect 324222 41420 324228 41432
rect 324280 41420 324286 41472
rect 326062 41420 326068 41472
rect 326120 41460 326126 41472
rect 326890 41460 326896 41472
rect 326120 41432 326896 41460
rect 326120 41420 326126 41432
rect 326890 41420 326896 41432
rect 326948 41420 326954 41472
rect 329006 41420 329012 41472
rect 329064 41460 329070 41472
rect 329742 41460 329748 41472
rect 329064 41432 329748 41460
rect 329064 41420 329070 41432
rect 329742 41420 329748 41432
rect 329800 41420 329806 41472
rect 329926 41420 329932 41472
rect 329984 41460 329990 41472
rect 331030 41460 331036 41472
rect 329984 41432 331036 41460
rect 329984 41420 329990 41432
rect 331030 41420 331036 41432
rect 331088 41420 331094 41472
rect 332870 41420 332876 41472
rect 332928 41460 332934 41472
rect 333790 41460 333796 41472
rect 332928 41432 333796 41460
rect 332928 41420 332934 41432
rect 333790 41420 333796 41432
rect 333848 41420 333854 41472
rect 335814 41420 335820 41472
rect 335872 41460 335878 41472
rect 336642 41460 336648 41472
rect 335872 41432 336648 41460
rect 335872 41420 335878 41432
rect 336642 41420 336648 41432
rect 336700 41420 336706 41472
rect 336826 41420 336832 41472
rect 336884 41460 336890 41472
rect 338022 41460 338028 41472
rect 336884 41432 338028 41460
rect 336884 41420 336890 41432
rect 338022 41420 338028 41432
rect 338080 41420 338086 41472
rect 339770 41420 339776 41472
rect 339828 41460 339834 41472
rect 340782 41460 340788 41472
rect 339828 41432 340788 41460
rect 339828 41420 339834 41432
rect 340782 41420 340788 41432
rect 340840 41420 340846 41472
rect 342714 41420 342720 41472
rect 342772 41460 342778 41472
rect 343542 41460 343548 41472
rect 342772 41432 343548 41460
rect 342772 41420 342778 41432
rect 343542 41420 343548 41432
rect 343600 41420 343606 41472
rect 343634 41420 343640 41472
rect 343692 41460 343698 41472
rect 344922 41460 344928 41472
rect 343692 41432 344928 41460
rect 343692 41420 343698 41432
rect 344922 41420 344928 41432
rect 344980 41420 344986 41472
rect 346578 41420 346584 41472
rect 346636 41460 346642 41472
rect 347682 41460 347688 41472
rect 346636 41432 347688 41460
rect 346636 41420 346642 41432
rect 347682 41420 347688 41432
rect 347740 41420 347746 41472
rect 349522 41420 349528 41472
rect 349580 41460 349586 41472
rect 350442 41460 350448 41472
rect 349580 41432 350448 41460
rect 349580 41420 349586 41432
rect 350442 41420 350448 41432
rect 350500 41420 350506 41472
rect 357434 41420 357440 41472
rect 357492 41460 357498 41472
rect 358722 41460 358728 41472
rect 357492 41432 358728 41460
rect 357492 41420 357498 41432
rect 358722 41420 358728 41432
rect 358780 41420 358786 41472
rect 360286 41420 360292 41472
rect 360344 41460 360350 41472
rect 361482 41460 361488 41472
rect 360344 41432 361488 41460
rect 360344 41420 360350 41432
rect 361482 41420 361488 41432
rect 361540 41420 361546 41472
rect 363230 41420 363236 41472
rect 363288 41460 363294 41472
rect 364242 41460 364248 41472
rect 363288 41432 364248 41460
rect 363288 41420 363294 41432
rect 364242 41420 364248 41432
rect 364300 41420 364306 41472
rect 366174 41420 366180 41472
rect 366232 41460 366238 41472
rect 367002 41460 367008 41472
rect 366232 41432 367008 41460
rect 366232 41420 366238 41432
rect 367002 41420 367008 41432
rect 367060 41420 367066 41472
rect 367186 41420 367192 41472
rect 367244 41460 367250 41472
rect 368382 41460 368388 41472
rect 367244 41432 368388 41460
rect 367244 41420 367250 41432
rect 368382 41420 368388 41432
rect 368440 41420 368446 41472
rect 370130 41420 370136 41472
rect 370188 41460 370194 41472
rect 371142 41460 371148 41472
rect 370188 41432 371148 41460
rect 370188 41420 370194 41432
rect 371142 41420 371148 41432
rect 371200 41420 371206 41472
rect 373074 41420 373080 41472
rect 373132 41460 373138 41472
rect 373902 41460 373908 41472
rect 373132 41432 373908 41460
rect 373132 41420 373138 41432
rect 373902 41420 373908 41432
rect 373960 41420 373966 41472
rect 380894 41420 380900 41472
rect 380952 41460 380958 41472
rect 382182 41460 382188 41472
rect 380952 41432 382188 41460
rect 380952 41420 380958 41432
rect 382182 41420 382188 41432
rect 382240 41420 382246 41472
rect 383838 41420 383844 41472
rect 383896 41460 383902 41472
rect 384942 41460 384948 41472
rect 383896 41432 384948 41460
rect 383896 41420 383902 41432
rect 384942 41420 384948 41432
rect 385000 41420 385006 41472
rect 386782 41420 386788 41472
rect 386840 41460 386846 41472
rect 387702 41460 387708 41472
rect 386840 41432 387708 41460
rect 386840 41420 386846 41432
rect 387702 41420 387708 41432
rect 387760 41420 387766 41472
rect 387794 41420 387800 41472
rect 387852 41460 387858 41472
rect 389082 41460 389088 41472
rect 387852 41432 389088 41460
rect 387852 41420 387858 41432
rect 389082 41420 389088 41432
rect 389140 41420 389146 41472
rect 389726 41420 389732 41472
rect 389784 41460 389790 41472
rect 390462 41460 390468 41472
rect 389784 41432 390468 41460
rect 389784 41420 389790 41432
rect 390462 41420 390468 41432
rect 390520 41420 390526 41472
rect 390738 41420 390744 41472
rect 390796 41460 390802 41472
rect 391842 41460 391848 41472
rect 390796 41432 391848 41460
rect 390796 41420 390802 41432
rect 391842 41420 391848 41432
rect 391900 41420 391906 41472
rect 393590 41420 393596 41472
rect 393648 41460 393654 41472
rect 394602 41460 394608 41472
rect 393648 41432 394608 41460
rect 393648 41420 393654 41432
rect 394602 41420 394608 41432
rect 394660 41420 394666 41472
rect 397546 41420 397552 41472
rect 397604 41460 397610 41472
rect 398650 41460 398656 41472
rect 397604 41432 398656 41460
rect 397604 41420 397610 41432
rect 398650 41420 398656 41432
rect 398708 41420 398714 41472
rect 399404 41324 399432 41500
rect 436738 41488 436744 41540
rect 436796 41528 436802 41540
rect 443638 41528 443644 41540
rect 436796 41500 443644 41528
rect 436796 41488 436802 41500
rect 443638 41488 443644 41500
rect 443696 41488 443702 41540
rect 410242 41420 410248 41472
rect 410300 41460 410306 41472
rect 411162 41460 411168 41472
rect 410300 41432 411168 41460
rect 410300 41420 410306 41432
rect 411162 41420 411168 41432
rect 411220 41420 411226 41472
rect 420086 41420 420092 41472
rect 420144 41460 420150 41472
rect 420822 41460 420828 41472
rect 420144 41432 420828 41460
rect 420144 41420 420150 41432
rect 420822 41420 420828 41432
rect 420880 41420 420886 41472
rect 421098 41420 421104 41472
rect 421156 41460 421162 41472
rect 422110 41460 422116 41472
rect 421156 41432 422116 41460
rect 421156 41420 421162 41432
rect 422110 41420 422116 41432
rect 422168 41420 422174 41472
rect 424042 41420 424048 41472
rect 424100 41460 424106 41472
rect 424870 41460 424876 41472
rect 424100 41432 424876 41460
rect 424100 41420 424106 41432
rect 424870 41420 424876 41432
rect 424928 41420 424934 41472
rect 426894 41420 426900 41472
rect 426952 41460 426958 41472
rect 427722 41460 427728 41472
rect 426952 41432 427728 41460
rect 426952 41420 426958 41432
rect 427722 41420 427728 41432
rect 427780 41420 427786 41472
rect 427906 41420 427912 41472
rect 427964 41460 427970 41472
rect 429102 41460 429108 41472
rect 427964 41432 429108 41460
rect 427964 41420 427970 41432
rect 429102 41420 429108 41432
rect 429160 41420 429166 41472
rect 430850 41420 430856 41472
rect 430908 41460 430914 41472
rect 431862 41460 431868 41472
rect 430908 41432 431868 41460
rect 430908 41420 430914 41432
rect 431862 41420 431868 41432
rect 431920 41420 431926 41472
rect 433794 41420 433800 41472
rect 433852 41460 433858 41472
rect 434622 41460 434628 41472
rect 433852 41432 434628 41460
rect 433852 41420 433858 41432
rect 434622 41420 434628 41432
rect 434680 41420 434686 41472
rect 437750 41420 437756 41472
rect 437808 41460 437814 41472
rect 438762 41460 438768 41472
rect 437808 41432 438768 41460
rect 437808 41420 437814 41432
rect 438762 41420 438768 41432
rect 438820 41420 438826 41472
rect 441614 41420 441620 41472
rect 441672 41460 441678 41472
rect 442810 41460 442816 41472
rect 441672 41432 442816 41460
rect 441672 41420 441678 41432
rect 442810 41420 442816 41432
rect 442868 41420 442874 41472
rect 444558 41420 444564 41472
rect 444616 41460 444622 41472
rect 445662 41460 445668 41472
rect 444616 41432 445668 41460
rect 444616 41420 444622 41432
rect 445662 41420 445668 41432
rect 445720 41420 445726 41472
rect 447502 41420 447508 41472
rect 447560 41460 447566 41472
rect 448422 41460 448428 41472
rect 447560 41432 448428 41460
rect 447560 41420 447566 41432
rect 448422 41420 448428 41432
rect 448480 41420 448486 41472
rect 448514 41420 448520 41472
rect 448572 41460 448578 41472
rect 449710 41460 449716 41472
rect 448572 41432 449716 41460
rect 448572 41420 448578 41432
rect 449710 41420 449716 41432
rect 449768 41420 449774 41472
rect 450446 41420 450452 41472
rect 450504 41460 450510 41472
rect 451182 41460 451188 41472
rect 450504 41432 451188 41460
rect 450504 41420 450510 41432
rect 451182 41420 451188 41432
rect 451240 41420 451246 41472
rect 451458 41420 451464 41472
rect 451516 41460 451522 41472
rect 452562 41460 452568 41472
rect 451516 41432 452568 41460
rect 451516 41420 451522 41432
rect 452562 41420 452568 41432
rect 452620 41420 452626 41472
rect 454402 41420 454408 41472
rect 454460 41460 454466 41472
rect 455322 41460 455328 41472
rect 454460 41432 455328 41460
rect 454460 41420 454466 41432
rect 455322 41420 455328 41432
rect 455380 41420 455386 41472
rect 465166 41420 465172 41472
rect 465224 41460 465230 41472
rect 466270 41460 466276 41472
rect 465224 41432 466276 41460
rect 465224 41420 465230 41432
rect 466270 41420 466276 41432
rect 466328 41420 466334 41472
rect 468110 41420 468116 41472
rect 468168 41460 468174 41472
rect 469122 41460 469128 41472
rect 468168 41432 469128 41460
rect 468168 41420 468174 41432
rect 469122 41420 469128 41432
rect 469180 41420 469186 41472
rect 471054 41420 471060 41472
rect 471112 41460 471118 41472
rect 471882 41460 471888 41472
rect 471112 41432 471888 41460
rect 471112 41420 471118 41432
rect 471882 41420 471888 41432
rect 471940 41420 471946 41472
rect 474918 41420 474924 41472
rect 474976 41460 474982 41472
rect 476022 41460 476028 41472
rect 474976 41432 476028 41460
rect 474976 41420 474982 41432
rect 476022 41420 476028 41432
rect 476080 41420 476086 41472
rect 480806 41420 480812 41472
rect 480864 41460 480870 41472
rect 481542 41460 481548 41472
rect 480864 41432 481548 41460
rect 480864 41420 480870 41432
rect 481542 41420 481548 41432
rect 481600 41420 481606 41472
rect 481818 41420 481824 41472
rect 481876 41460 481882 41472
rect 482922 41460 482928 41472
rect 481876 41432 482928 41460
rect 481876 41420 481882 41432
rect 482922 41420 482928 41432
rect 482980 41420 482986 41472
rect 488626 41420 488632 41472
rect 488684 41460 488690 41472
rect 489730 41460 489736 41472
rect 488684 41432 489736 41460
rect 488684 41420 488690 41432
rect 489730 41420 489736 41432
rect 489788 41420 489794 41472
rect 491570 41420 491576 41472
rect 491628 41460 491634 41472
rect 492490 41460 492496 41472
rect 491628 41432 492496 41460
rect 491628 41420 491634 41432
rect 492490 41420 492496 41432
rect 492548 41420 492554 41472
rect 494514 41420 494520 41472
rect 494572 41460 494578 41472
rect 495342 41460 495348 41472
rect 494572 41432 495348 41460
rect 494572 41420 494578 41432
rect 495342 41420 495348 41432
rect 495400 41420 495406 41472
rect 498470 41420 498476 41472
rect 498528 41460 498534 41472
rect 499482 41460 499488 41472
rect 498528 41432 499488 41460
rect 498528 41420 498534 41432
rect 499482 41420 499488 41432
rect 499540 41420 499546 41472
rect 505278 41420 505284 41472
rect 505336 41460 505342 41472
rect 506382 41460 506388 41472
rect 505336 41432 506388 41460
rect 505336 41420 505342 41432
rect 506382 41420 506388 41432
rect 506440 41420 506446 41472
rect 509234 41420 509240 41472
rect 509292 41460 509298 41472
rect 510430 41460 510436 41472
rect 509292 41432 510436 41460
rect 509292 41420 509298 41432
rect 510430 41420 510436 41432
rect 510488 41420 510494 41472
rect 511166 41420 511172 41472
rect 511224 41460 511230 41472
rect 511902 41460 511908 41472
rect 511224 41432 511908 41460
rect 511224 41420 511230 41432
rect 511902 41420 511908 41432
rect 511960 41420 511966 41472
rect 512178 41420 512184 41472
rect 512236 41460 512242 41472
rect 513282 41460 513288 41472
rect 512236 41432 513288 41460
rect 512236 41420 512242 41432
rect 513282 41420 513288 41432
rect 513340 41420 513346 41472
rect 515122 41420 515128 41472
rect 515180 41460 515186 41472
rect 515950 41460 515956 41472
rect 515180 41432 515956 41460
rect 515180 41420 515186 41432
rect 515950 41420 515956 41432
rect 516008 41420 516014 41472
rect 521930 41420 521936 41472
rect 521988 41460 521994 41472
rect 522942 41460 522948 41472
rect 521988 41432 522948 41460
rect 521988 41420 521994 41432
rect 522942 41420 522948 41432
rect 523000 41420 523006 41472
rect 399478 41324 399484 41336
rect 399404 41296 399484 41324
rect 399478 41284 399484 41296
rect 399536 41284 399542 41336
rect 238846 39992 238852 40044
rect 238904 40032 238910 40044
rect 239582 40032 239588 40044
rect 238904 40004 239588 40032
rect 238904 39992 238910 40004
rect 239582 39992 239588 40004
rect 239640 39992 239646 40044
rect 108942 38672 108948 38684
rect 108903 38644 108948 38672
rect 108942 38632 108948 38644
rect 109000 38632 109006 38684
rect 31662 38604 31668 38616
rect 31623 38576 31668 38604
rect 31662 38564 31668 38576
rect 31720 38564 31726 38616
rect 53285 38607 53343 38613
rect 53285 38573 53297 38607
rect 53331 38604 53343 38607
rect 53374 38604 53380 38616
rect 53331 38576 53380 38604
rect 53331 38573 53343 38576
rect 53285 38567 53343 38573
rect 53374 38564 53380 38576
rect 53432 38564 53438 38616
rect 73522 38604 73528 38616
rect 73483 38576 73528 38604
rect 73522 38564 73528 38576
rect 73580 38564 73586 38616
rect 75730 38564 75736 38616
rect 75788 38604 75794 38616
rect 75822 38604 75828 38616
rect 75788 38576 75828 38604
rect 75788 38564 75794 38576
rect 75822 38564 75828 38576
rect 75880 38564 75886 38616
rect 244274 38564 244280 38616
rect 244332 38604 244338 38616
rect 244366 38604 244372 38616
rect 244332 38576 244372 38604
rect 244332 38564 244338 38576
rect 244366 38564 244372 38576
rect 244424 38564 244430 38616
rect 245933 38607 245991 38613
rect 245933 38573 245945 38607
rect 245979 38604 245991 38607
rect 246022 38604 246028 38616
rect 245979 38576 246028 38604
rect 245979 38573 245991 38576
rect 245933 38567 245991 38573
rect 246022 38564 246028 38576
rect 246080 38564 246086 38616
rect 108942 38536 108948 38548
rect 108903 38508 108948 38536
rect 108942 38496 108948 38508
rect 109000 38496 109006 38548
rect 75730 37204 75736 37256
rect 75788 37244 75794 37256
rect 244366 37244 244372 37256
rect 75788 37216 75833 37244
rect 244327 37216 244372 37244
rect 75788 37204 75794 37216
rect 244366 37204 244372 37216
rect 244424 37204 244430 37256
rect 433426 37244 433432 37256
rect 433387 37216 433432 37244
rect 433426 37204 433432 37216
rect 433484 37204 433490 37256
rect 241606 35912 241612 35964
rect 241664 35952 241670 35964
rect 242526 35952 242532 35964
rect 241664 35924 242532 35952
rect 241664 35912 241670 35924
rect 242526 35912 242532 35924
rect 242584 35912 242590 35964
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 25498 35884 25504 35896
rect 3476 35856 25504 35884
rect 3476 35844 3482 35856
rect 25498 35844 25504 35856
rect 25556 35844 25562 35896
rect 175001 35887 175059 35893
rect 175001 35853 175013 35887
rect 175047 35884 175059 35887
rect 175182 35884 175188 35896
rect 175047 35856 175188 35884
rect 175047 35853 175059 35856
rect 175001 35847 175059 35853
rect 175182 35844 175188 35856
rect 175240 35844 175246 35896
rect 56870 31764 56876 31816
rect 56928 31804 56934 31816
rect 57422 31804 57428 31816
rect 56928 31776 57428 31804
rect 56928 31764 56934 31776
rect 57422 31764 57428 31776
rect 57480 31764 57486 31816
rect 31662 29016 31668 29028
rect 31623 28988 31668 29016
rect 31662 28976 31668 28988
rect 31720 28976 31726 29028
rect 53282 29016 53288 29028
rect 53243 28988 53288 29016
rect 53282 28976 53288 28988
rect 53340 28976 53346 29028
rect 73525 29019 73583 29025
rect 73525 28985 73537 29019
rect 73571 29016 73583 29019
rect 73614 29016 73620 29028
rect 73571 28988 73620 29016
rect 73571 28985 73583 28988
rect 73525 28979 73583 28985
rect 73614 28976 73620 28988
rect 73672 28976 73678 29028
rect 96614 28976 96620 29028
rect 96672 29016 96678 29028
rect 97534 29016 97540 29028
rect 96672 28988 97540 29016
rect 96672 28976 96678 28988
rect 97534 28976 97540 28988
rect 97592 28976 97598 29028
rect 108942 29016 108948 29028
rect 108903 28988 108948 29016
rect 108942 28976 108948 28988
rect 109000 28976 109006 29028
rect 174998 29016 175004 29028
rect 174959 28988 175004 29016
rect 174998 28976 175004 28988
rect 175056 28976 175062 29028
rect 245930 29016 245936 29028
rect 245891 28988 245936 29016
rect 245930 28976 245936 28988
rect 245988 28976 245994 29028
rect 75733 27659 75791 27665
rect 75733 27625 75745 27659
rect 75779 27656 75791 27659
rect 75822 27656 75828 27668
rect 75779 27628 75828 27656
rect 75779 27625 75791 27628
rect 75733 27619 75791 27625
rect 75822 27616 75828 27628
rect 75880 27616 75886 27668
rect 244274 27616 244280 27668
rect 244332 27656 244338 27668
rect 244369 27659 244427 27665
rect 244369 27656 244381 27659
rect 244332 27628 244381 27656
rect 244332 27616 244338 27628
rect 244369 27625 244381 27628
rect 244415 27625 244427 27659
rect 433426 27656 433432 27668
rect 433387 27628 433432 27656
rect 244369 27619 244427 27625
rect 433426 27616 433432 27628
rect 433484 27616 433490 27668
rect 117406 27548 117412 27600
rect 117464 27588 117470 27600
rect 117685 27591 117743 27597
rect 117685 27588 117697 27591
rect 117464 27560 117697 27588
rect 117464 27548 117470 27560
rect 117685 27557 117697 27560
rect 117731 27557 117743 27591
rect 117685 27551 117743 27557
rect 120166 27548 120172 27600
rect 120224 27588 120230 27600
rect 120445 27591 120503 27597
rect 120445 27588 120457 27591
rect 120224 27560 120457 27588
rect 120224 27548 120230 27560
rect 120445 27557 120457 27560
rect 120491 27557 120503 27591
rect 120445 27551 120503 27557
rect 244274 22760 244280 22772
rect 244235 22732 244280 22760
rect 244274 22720 244280 22732
rect 244332 22720 244338 22772
rect 52546 22108 52552 22160
rect 52604 22148 52610 22160
rect 53282 22148 53288 22160
rect 52604 22120 53288 22148
rect 52604 22108 52610 22120
rect 53282 22108 53288 22120
rect 53340 22108 53346 22160
rect 174998 22148 175004 22160
rect 174832 22120 175004 22148
rect 174832 22092 174860 22120
rect 174998 22108 175004 22120
rect 175056 22108 175062 22160
rect 174814 22040 174820 22092
rect 174872 22040 174878 22092
rect 245838 22040 245844 22092
rect 245896 22080 245902 22092
rect 246022 22080 246028 22092
rect 245896 22052 246028 22080
rect 245896 22040 245902 22052
rect 246022 22040 246028 22052
rect 246080 22040 246086 22092
rect 75457 20995 75515 21001
rect 75457 20961 75469 20995
rect 75503 20992 75515 20995
rect 75822 20992 75828 21004
rect 75503 20964 75828 20992
rect 75503 20961 75515 20964
rect 75457 20955 75515 20961
rect 75822 20952 75828 20964
rect 75880 20952 75886 21004
rect 100662 19524 100668 19576
rect 100720 19524 100726 19576
rect 100680 19440 100708 19524
rect 100662 19388 100668 19440
rect 100720 19388 100726 19440
rect 96614 19320 96620 19372
rect 96672 19360 96678 19372
rect 96706 19360 96712 19372
rect 96672 19332 96712 19360
rect 96672 19320 96678 19332
rect 96706 19320 96712 19332
rect 96764 19320 96770 19372
rect 31478 19252 31484 19304
rect 31536 19292 31542 19304
rect 31662 19292 31668 19304
rect 31536 19264 31668 19292
rect 31536 19252 31542 19264
rect 31662 19252 31668 19264
rect 31720 19252 31726 19304
rect 108758 19252 108764 19304
rect 108816 19292 108822 19304
rect 108942 19292 108948 19304
rect 108816 19264 108948 19292
rect 108816 19252 108822 19264
rect 108942 19252 108948 19264
rect 109000 19252 109006 19304
rect 246022 19292 246028 19304
rect 245983 19264 246028 19292
rect 246022 19252 246028 19264
rect 246080 19252 246086 19304
rect 404449 19295 404507 19301
rect 404449 19261 404461 19295
rect 404495 19292 404507 19295
rect 404722 19292 404728 19304
rect 404495 19264 404728 19292
rect 404495 19261 404507 19264
rect 404449 19255 404507 19261
rect 404722 19252 404728 19264
rect 404780 19252 404786 19304
rect 433426 17932 433432 17944
rect 433387 17904 433432 17932
rect 433426 17892 433432 17904
rect 433484 17892 433490 17944
rect 522298 17892 522304 17944
rect 522356 17932 522362 17944
rect 579798 17932 579804 17944
rect 522356 17904 579804 17932
rect 522356 17892 522362 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 120442 12424 120448 12436
rect 120403 12396 120448 12424
rect 120442 12384 120448 12396
rect 120500 12384 120506 12436
rect 125318 12384 125324 12436
rect 125376 12424 125382 12436
rect 125502 12424 125508 12436
rect 125376 12396 125508 12424
rect 125376 12384 125382 12396
rect 125502 12384 125508 12396
rect 125560 12384 125566 12436
rect 252278 12384 252284 12436
rect 252336 12424 252342 12436
rect 252462 12424 252468 12436
rect 252336 12396 252468 12424
rect 252336 12384 252342 12396
rect 252462 12384 252468 12396
rect 252520 12384 252526 12436
rect 75454 9704 75460 9716
rect 75415 9676 75460 9704
rect 75454 9664 75460 9676
rect 75512 9664 75518 9716
rect 117682 9704 117688 9716
rect 117643 9676 117688 9704
rect 117682 9664 117688 9676
rect 117740 9664 117746 9716
rect 244277 9707 244335 9713
rect 244277 9673 244289 9707
rect 244323 9704 244335 9707
rect 244366 9704 244372 9716
rect 244323 9676 244372 9704
rect 244323 9673 244335 9676
rect 244277 9667 244335 9673
rect 244366 9664 244372 9676
rect 244424 9664 244430 9716
rect 246022 9704 246028 9716
rect 245983 9676 246028 9704
rect 246022 9664 246028 9676
rect 246080 9664 246086 9716
rect 404446 9704 404452 9716
rect 404407 9676 404452 9704
rect 404446 9664 404452 9676
rect 404504 9664 404510 9716
rect 31481 9639 31539 9645
rect 31481 9605 31493 9639
rect 31527 9636 31539 9639
rect 31662 9636 31668 9648
rect 31527 9608 31668 9636
rect 31527 9605 31539 9608
rect 31481 9599 31539 9605
rect 31662 9596 31668 9608
rect 31720 9596 31726 9648
rect 100481 9639 100539 9645
rect 100481 9605 100493 9639
rect 100527 9636 100539 9639
rect 100662 9636 100668 9648
rect 100527 9608 100668 9636
rect 100527 9605 100539 9608
rect 100481 9599 100539 9605
rect 100662 9596 100668 9608
rect 100720 9596 100726 9648
rect 108761 9639 108819 9645
rect 108761 9605 108773 9639
rect 108807 9636 108819 9639
rect 108942 9636 108948 9648
rect 108807 9608 108948 9636
rect 108807 9605 108819 9608
rect 108761 9599 108819 9605
rect 108942 9596 108948 9608
rect 109000 9596 109006 9648
rect 433426 8412 433432 8424
rect 433387 8384 433432 8412
rect 433426 8372 433432 8384
rect 433484 8372 433490 8424
rect 433426 8236 433432 8288
rect 433484 8276 433490 8288
rect 433521 8279 433579 8285
rect 433521 8276 433533 8279
rect 433484 8248 433533 8276
rect 433484 8236 433490 8248
rect 433521 8245 433533 8248
rect 433567 8245 433579 8279
rect 433521 8239 433579 8245
rect 471882 6536 471888 6588
rect 471940 6576 471946 6588
rect 519078 6576 519084 6588
rect 471940 6548 519084 6576
rect 471940 6536 471946 6548
rect 519078 6536 519084 6548
rect 519136 6536 519142 6588
rect 474642 6468 474648 6520
rect 474700 6508 474706 6520
rect 522666 6508 522672 6520
rect 474700 6480 522672 6508
rect 474700 6468 474706 6480
rect 522666 6468 522672 6480
rect 522724 6468 522730 6520
rect 477402 6400 477408 6452
rect 477460 6440 477466 6452
rect 526254 6440 526260 6452
rect 477460 6412 526260 6440
rect 477460 6400 477466 6412
rect 526254 6400 526260 6412
rect 526312 6400 526318 6452
rect 513282 6332 513288 6384
rect 513340 6372 513346 6384
rect 569034 6372 569040 6384
rect 513340 6344 569040 6372
rect 513340 6332 513346 6344
rect 569034 6332 569040 6344
rect 569092 6332 569098 6384
rect 515950 6264 515956 6316
rect 516008 6304 516014 6316
rect 572622 6304 572628 6316
rect 516008 6276 572628 6304
rect 516008 6264 516014 6276
rect 572622 6264 572628 6276
rect 572680 6264 572686 6316
rect 506290 6196 506296 6248
rect 506348 6236 506354 6248
rect 561950 6236 561956 6248
rect 506348 6208 561956 6236
rect 506348 6196 506354 6208
rect 561950 6196 561956 6208
rect 562008 6196 562014 6248
rect 469122 6128 469128 6180
rect 469180 6168 469186 6180
rect 515582 6168 515588 6180
rect 469180 6140 515588 6168
rect 469180 6128 469186 6140
rect 515582 6128 515588 6140
rect 515640 6128 515646 6180
rect 518802 6128 518808 6180
rect 518860 6168 518866 6180
rect 576210 6168 576216 6180
rect 518860 6140 576216 6168
rect 518860 6128 518866 6140
rect 576210 6128 576216 6140
rect 576268 6128 576274 6180
rect 466270 5448 466276 5500
rect 466328 5488 466334 5500
rect 511994 5488 512000 5500
rect 466328 5460 512000 5488
rect 466328 5448 466334 5460
rect 511994 5448 512000 5460
rect 512052 5448 512058 5500
rect 452580 5392 454080 5420
rect 340506 5312 340512 5364
rect 340564 5352 340570 5364
rect 340782 5352 340788 5364
rect 340564 5324 340788 5352
rect 340564 5312 340570 5324
rect 340782 5312 340788 5324
rect 340840 5312 340846 5364
rect 422110 5312 422116 5364
rect 422168 5352 422174 5364
rect 437385 5355 437443 5361
rect 437385 5352 437397 5355
rect 422168 5324 437397 5352
rect 422168 5312 422174 5324
rect 437385 5321 437397 5324
rect 437431 5321 437443 5355
rect 437385 5315 437443 5321
rect 437477 5355 437535 5361
rect 437477 5321 437489 5355
rect 437523 5352 437535 5355
rect 442997 5355 443055 5361
rect 442997 5352 443009 5355
rect 437523 5324 443009 5352
rect 437523 5321 437535 5324
rect 437477 5315 437535 5321
rect 442997 5321 443009 5324
rect 443043 5321 443055 5355
rect 442997 5315 443055 5321
rect 445573 5355 445631 5361
rect 445573 5321 445585 5355
rect 445619 5352 445631 5355
rect 452580 5352 452608 5392
rect 454052 5361 454080 5392
rect 480162 5380 480168 5432
rect 480220 5420 480226 5432
rect 529842 5420 529848 5432
rect 480220 5392 529848 5420
rect 480220 5380 480226 5392
rect 529842 5380 529848 5392
rect 529900 5380 529906 5432
rect 445619 5324 452608 5352
rect 454037 5355 454095 5361
rect 445619 5321 445631 5324
rect 445573 5315 445631 5321
rect 454037 5321 454049 5355
rect 454083 5321 454095 5355
rect 454037 5315 454095 5321
rect 489730 5312 489736 5364
rect 489788 5352 489794 5364
rect 540514 5352 540520 5364
rect 489788 5324 540520 5352
rect 489788 5312 489794 5324
rect 540514 5312 540520 5324
rect 540572 5312 540578 5364
rect 37366 5244 37372 5296
rect 37424 5284 37430 5296
rect 73246 5284 73252 5296
rect 37424 5256 73252 5284
rect 37424 5244 37430 5256
rect 73246 5244 73252 5256
rect 73304 5244 73310 5296
rect 456702 5244 456708 5296
rect 456760 5284 456766 5296
rect 462317 5287 462375 5293
rect 462317 5284 462329 5287
rect 456760 5256 462329 5284
rect 456760 5244 456766 5256
rect 462317 5253 462329 5256
rect 462363 5253 462375 5287
rect 462317 5247 462375 5253
rect 482830 5244 482836 5296
rect 482888 5284 482894 5296
rect 533430 5284 533436 5296
rect 482888 5256 533436 5284
rect 482888 5244 482894 5256
rect 533430 5244 533436 5256
rect 533488 5244 533494 5296
rect 33870 5176 33876 5228
rect 33928 5216 33934 5228
rect 70486 5216 70492 5228
rect 33928 5188 70492 5216
rect 33928 5176 33934 5188
rect 70486 5176 70492 5188
rect 70544 5176 70550 5228
rect 398650 5176 398656 5228
rect 398708 5216 398714 5228
rect 429930 5216 429936 5228
rect 398708 5188 429936 5216
rect 398708 5176 398714 5188
rect 429930 5176 429936 5188
rect 429988 5176 429994 5228
rect 442997 5219 443055 5225
rect 442997 5185 443009 5219
rect 443043 5216 443055 5219
rect 445573 5219 445631 5225
rect 445573 5216 445585 5219
rect 443043 5188 445585 5216
rect 443043 5185 443055 5188
rect 442997 5179 443055 5185
rect 445573 5185 445585 5188
rect 445619 5185 445631 5219
rect 445573 5179 445631 5185
rect 445662 5176 445668 5228
rect 445720 5216 445726 5228
rect 486970 5216 486976 5228
rect 445720 5188 486976 5216
rect 445720 5176 445726 5188
rect 486970 5176 486976 5188
rect 487028 5176 487034 5228
rect 495342 5176 495348 5228
rect 495400 5216 495406 5228
rect 547690 5216 547696 5228
rect 495400 5188 547696 5216
rect 495400 5176 495406 5188
rect 547690 5176 547696 5188
rect 547748 5176 547754 5228
rect 30282 5108 30288 5160
rect 30340 5148 30346 5160
rect 67634 5148 67640 5160
rect 30340 5120 67640 5148
rect 30340 5108 30346 5120
rect 67634 5108 67640 5120
rect 67692 5108 67698 5160
rect 404262 5108 404268 5160
rect 404320 5148 404326 5160
rect 437014 5148 437020 5160
rect 404320 5120 437020 5148
rect 404320 5108 404326 5120
rect 437014 5108 437020 5120
rect 437072 5108 437078 5160
rect 442810 5108 442816 5160
rect 442868 5148 442874 5160
rect 483474 5148 483480 5160
rect 442868 5120 483480 5148
rect 442868 5108 442874 5120
rect 483474 5108 483480 5120
rect 483532 5108 483538 5160
rect 485682 5108 485688 5160
rect 485740 5148 485746 5160
rect 536926 5148 536932 5160
rect 485740 5120 536932 5148
rect 485740 5108 485746 5120
rect 536926 5108 536932 5120
rect 536984 5108 536990 5160
rect 26694 5040 26700 5092
rect 26752 5080 26758 5092
rect 64874 5080 64880 5092
rect 26752 5052 64880 5080
rect 26752 5040 26758 5052
rect 64874 5040 64880 5052
rect 64932 5040 64938 5092
rect 407022 5040 407028 5092
rect 407080 5080 407086 5092
rect 440602 5080 440608 5092
rect 407080 5052 440608 5080
rect 407080 5040 407086 5052
rect 440602 5040 440608 5052
rect 440660 5040 440666 5092
rect 448422 5040 448428 5092
rect 448480 5080 448486 5092
rect 490558 5080 490564 5092
rect 448480 5052 490564 5080
rect 448480 5040 448486 5052
rect 490558 5040 490564 5052
rect 490616 5040 490622 5092
rect 492490 5040 492496 5092
rect 492548 5080 492554 5092
rect 544102 5080 544108 5092
rect 492548 5052 544108 5080
rect 492548 5040 492554 5052
rect 544102 5040 544108 5052
rect 544160 5040 544166 5092
rect 22002 4972 22008 5024
rect 22060 5012 22066 5024
rect 60734 5012 60740 5024
rect 22060 4984 60740 5012
rect 22060 4972 22066 4984
rect 60734 4972 60740 4984
rect 60792 4972 60798 5024
rect 409782 4972 409788 5024
rect 409840 5012 409846 5024
rect 444190 5012 444196 5024
rect 409840 4984 444196 5012
rect 409840 4972 409846 4984
rect 444190 4972 444196 4984
rect 444248 4972 444254 5024
rect 453942 4972 453948 5024
rect 454000 5012 454006 5024
rect 497734 5012 497740 5024
rect 454000 4984 497740 5012
rect 454000 4972 454006 4984
rect 497734 4972 497740 4984
rect 497792 4972 497798 5024
rect 498102 4972 498108 5024
rect 498160 5012 498166 5024
rect 551186 5012 551192 5024
rect 498160 4984 551192 5012
rect 498160 4972 498166 4984
rect 551186 4972 551192 4984
rect 551244 4972 551250 5024
rect 17218 4904 17224 4956
rect 17276 4944 17282 4956
rect 56686 4944 56692 4956
rect 17276 4916 56692 4944
rect 17276 4904 17282 4916
rect 56686 4904 56692 4916
rect 56744 4904 56750 4956
rect 415302 4904 415308 4956
rect 415360 4944 415366 4956
rect 451274 4944 451280 4956
rect 415360 4916 451280 4944
rect 415360 4904 415366 4916
rect 451274 4904 451280 4916
rect 451332 4904 451338 4956
rect 454037 4947 454095 4953
rect 454037 4913 454049 4947
rect 454083 4944 454095 4947
rect 458450 4944 458456 4956
rect 454083 4916 458456 4944
rect 454083 4913 454095 4916
rect 454037 4907 454095 4913
rect 458450 4904 458456 4916
rect 458508 4904 458514 4956
rect 462317 4947 462375 4953
rect 462317 4913 462329 4947
rect 462363 4944 462375 4947
rect 501230 4944 501236 4956
rect 462363 4916 501236 4944
rect 462363 4913 462375 4916
rect 462317 4907 462375 4913
rect 501230 4904 501236 4916
rect 501288 4904 501294 4956
rect 503622 4904 503628 4956
rect 503680 4944 503686 4956
rect 558362 4944 558368 4956
rect 503680 4916 558368 4944
rect 503680 4904 503686 4916
rect 558362 4904 558368 4916
rect 558420 4904 558426 4956
rect 12434 4836 12440 4888
rect 12492 4876 12498 4888
rect 52638 4876 52644 4888
rect 12492 4848 52644 4876
rect 12492 4836 12498 4848
rect 52638 4836 52644 4848
rect 52696 4836 52702 4888
rect 412542 4836 412548 4888
rect 412600 4876 412606 4888
rect 447778 4876 447784 4888
rect 412600 4848 447784 4876
rect 412600 4836 412606 4848
rect 447778 4836 447784 4848
rect 447836 4836 447842 4888
rect 451182 4836 451188 4888
rect 451240 4876 451246 4888
rect 494146 4876 494152 4888
rect 451240 4848 494152 4876
rect 451240 4836 451246 4848
rect 494146 4836 494152 4848
rect 494204 4836 494210 4888
rect 500862 4836 500868 4888
rect 500920 4876 500926 4888
rect 554774 4876 554780 4888
rect 500920 4848 554780 4876
rect 500920 4836 500926 4848
rect 554774 4836 554780 4848
rect 554832 4836 554838 4888
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 49786 4808 49792 4820
rect 7708 4780 49792 4808
rect 7708 4768 7714 4780
rect 49786 4768 49792 4780
rect 49844 4768 49850 4820
rect 73062 4768 73068 4820
rect 73120 4808 73126 4820
rect 103606 4808 103612 4820
rect 73120 4780 103612 4808
rect 73120 4768 73126 4780
rect 103606 4768 103612 4780
rect 103664 4768 103670 4820
rect 391750 4768 391756 4820
rect 391808 4808 391814 4820
rect 422754 4808 422760 4820
rect 391808 4780 422760 4808
rect 391808 4768 391814 4780
rect 422754 4768 422760 4780
rect 422812 4768 422818 4820
rect 424870 4768 424876 4820
rect 424928 4808 424934 4820
rect 462038 4808 462044 4820
rect 424928 4780 462044 4808
rect 424928 4768 424934 4780
rect 462038 4768 462044 4780
rect 462096 4768 462102 4820
rect 462222 4768 462228 4820
rect 462280 4808 462286 4820
rect 508406 4808 508412 4820
rect 462280 4780 508412 4808
rect 462280 4768 462286 4780
rect 508406 4768 508412 4780
rect 508464 4768 508470 4820
rect 510430 4768 510436 4820
rect 510488 4808 510494 4820
rect 565538 4808 565544 4820
rect 510488 4780 565544 4808
rect 510488 4768 510494 4780
rect 565538 4768 565544 4780
rect 565596 4768 565602 4820
rect 459462 4700 459468 4752
rect 459520 4740 459526 4752
rect 504818 4740 504824 4752
rect 459520 4712 504824 4740
rect 459520 4700 459526 4712
rect 504818 4700 504824 4712
rect 504876 4700 504882 4752
rect 115937 4403 115995 4409
rect 115937 4369 115949 4403
rect 115983 4400 115995 4403
rect 120442 4400 120448 4412
rect 115983 4372 120448 4400
rect 115983 4369 115995 4372
rect 115937 4363 115995 4369
rect 120442 4360 120448 4372
rect 120500 4360 120506 4412
rect 437477 4199 437535 4205
rect 437477 4165 437489 4199
rect 437523 4196 437535 4199
rect 445481 4199 445539 4205
rect 445481 4196 445493 4199
rect 437523 4168 445493 4196
rect 437523 4165 437535 4168
rect 437477 4159 437535 4165
rect 445481 4165 445493 4168
rect 445527 4165 445539 4199
rect 445481 4159 445539 4165
rect 16022 4088 16028 4140
rect 16080 4128 16086 4140
rect 16482 4128 16488 4140
rect 16080 4100 16488 4128
rect 16080 4088 16086 4100
rect 16482 4088 16488 4100
rect 16540 4088 16546 4140
rect 18322 4088 18328 4140
rect 18380 4128 18386 4140
rect 19242 4128 19248 4140
rect 18380 4100 19248 4128
rect 18380 4088 18386 4100
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 19518 4088 19524 4140
rect 19576 4128 19582 4140
rect 20622 4128 20628 4140
rect 19576 4100 20628 4128
rect 19576 4088 19582 4100
rect 20622 4088 20628 4100
rect 20680 4088 20686 4140
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 21910 4128 21916 4140
rect 20772 4100 21916 4128
rect 20772 4088 20778 4100
rect 21910 4088 21916 4100
rect 21968 4088 21974 4140
rect 36170 4088 36176 4140
rect 36228 4128 36234 4140
rect 36228 4100 39436 4128
rect 36228 4088 36234 4100
rect 29086 4020 29092 4072
rect 29144 4060 29150 4072
rect 39298 4060 39304 4072
rect 29144 4032 39304 4060
rect 29144 4020 29150 4032
rect 39298 4020 39304 4032
rect 39356 4020 39362 4072
rect 39408 4060 39436 4100
rect 54018 4088 54024 4140
rect 54076 4128 54082 4140
rect 55122 4128 55128 4140
rect 54076 4100 55128 4128
rect 54076 4088 54082 4100
rect 55122 4088 55128 4100
rect 55180 4088 55186 4140
rect 59998 4088 60004 4140
rect 60056 4128 60062 4140
rect 60642 4128 60648 4140
rect 60056 4100 60648 4128
rect 60056 4088 60062 4100
rect 60642 4088 60648 4100
rect 60700 4088 60706 4140
rect 71866 4088 71872 4140
rect 71924 4128 71930 4140
rect 73798 4128 73804 4140
rect 71924 4100 73804 4128
rect 71924 4088 71930 4100
rect 73798 4088 73804 4100
rect 73856 4088 73862 4140
rect 75181 4131 75239 4137
rect 75181 4097 75193 4131
rect 75227 4128 75239 4131
rect 80698 4128 80704 4140
rect 75227 4100 80704 4128
rect 75227 4097 75239 4100
rect 75181 4091 75239 4097
rect 80698 4088 80704 4100
rect 80756 4088 80762 4140
rect 84930 4088 84936 4140
rect 84988 4128 84994 4140
rect 85482 4128 85488 4140
rect 84988 4100 85488 4128
rect 84988 4088 84994 4100
rect 85482 4088 85488 4100
rect 85540 4088 85546 4140
rect 86126 4088 86132 4140
rect 86184 4128 86190 4140
rect 86862 4128 86868 4140
rect 86184 4100 86868 4128
rect 86184 4088 86190 4100
rect 86862 4088 86868 4100
rect 86920 4088 86926 4140
rect 93302 4088 93308 4140
rect 93360 4128 93366 4140
rect 93762 4128 93768 4140
rect 93360 4100 93768 4128
rect 93360 4088 93366 4100
rect 93762 4088 93768 4100
rect 93820 4088 93826 4140
rect 96890 4088 96896 4140
rect 96948 4128 96954 4140
rect 97902 4128 97908 4140
rect 96948 4100 97908 4128
rect 96948 4088 96954 4100
rect 97902 4088 97908 4100
rect 97960 4088 97966 4140
rect 102778 4088 102784 4140
rect 102836 4128 102842 4140
rect 103422 4128 103428 4140
rect 102836 4100 103428 4128
rect 102836 4088 102842 4100
rect 103422 4088 103428 4100
rect 103480 4088 103486 4140
rect 106366 4088 106372 4140
rect 106424 4128 106430 4140
rect 107470 4128 107476 4140
rect 106424 4100 107476 4128
rect 106424 4088 106430 4100
rect 107470 4088 107476 4100
rect 107528 4088 107534 4140
rect 111150 4088 111156 4140
rect 111208 4128 111214 4140
rect 111702 4128 111708 4140
rect 111208 4100 111708 4128
rect 111208 4088 111214 4100
rect 111702 4088 111708 4100
rect 111760 4088 111766 4140
rect 112346 4088 112352 4140
rect 112404 4128 112410 4140
rect 113082 4128 113088 4140
rect 112404 4100 113088 4128
rect 112404 4088 112410 4100
rect 113082 4088 113088 4100
rect 113140 4088 113146 4140
rect 113542 4088 113548 4140
rect 113600 4128 113606 4140
rect 114462 4128 114468 4140
rect 113600 4100 114468 4128
rect 113600 4088 113606 4100
rect 114462 4088 114468 4100
rect 114520 4088 114526 4140
rect 115934 4088 115940 4140
rect 115992 4128 115998 4140
rect 117222 4128 117228 4140
rect 115992 4100 117228 4128
rect 115992 4088 115998 4100
rect 117222 4088 117228 4100
rect 117280 4088 117286 4140
rect 119430 4088 119436 4140
rect 119488 4128 119494 4140
rect 119982 4128 119988 4140
rect 119488 4100 119988 4128
rect 119488 4088 119494 4100
rect 119982 4088 119988 4100
rect 120040 4088 120046 4140
rect 127802 4088 127808 4140
rect 127860 4128 127866 4140
rect 128262 4128 128268 4140
rect 127860 4100 128268 4128
rect 127860 4088 127866 4100
rect 128262 4088 128268 4100
rect 128320 4088 128326 4140
rect 170582 4088 170588 4140
rect 170640 4128 170646 4140
rect 171042 4128 171048 4140
rect 170640 4100 171048 4128
rect 170640 4088 170646 4100
rect 171042 4088 171048 4100
rect 171100 4088 171106 4140
rect 171778 4088 171784 4140
rect 171836 4128 171842 4140
rect 172422 4128 172428 4140
rect 171836 4100 172428 4128
rect 171836 4088 171842 4100
rect 172422 4088 172428 4100
rect 172480 4088 172486 4140
rect 238386 4088 238392 4140
rect 238444 4128 238450 4140
rect 238846 4128 238852 4140
rect 238444 4100 238852 4128
rect 238444 4088 238450 4100
rect 238846 4088 238852 4100
rect 238904 4088 238910 4140
rect 240778 4088 240784 4140
rect 240836 4128 240842 4140
rect 241422 4128 241428 4140
rect 240836 4100 241428 4128
rect 240836 4088 240842 4100
rect 241422 4088 241428 4100
rect 241480 4088 241486 4140
rect 246022 4088 246028 4140
rect 246080 4128 246086 4140
rect 246758 4128 246764 4140
rect 246080 4100 246764 4128
rect 246080 4088 246086 4100
rect 246758 4088 246764 4100
rect 246816 4088 246822 4140
rect 247034 4088 247040 4140
rect 247092 4128 247098 4140
rect 247954 4128 247960 4140
rect 247092 4100 247960 4128
rect 247092 4088 247098 4100
rect 247954 4088 247960 4100
rect 248012 4088 248018 4140
rect 248506 4088 248512 4140
rect 248564 4128 248570 4140
rect 249150 4128 249156 4140
rect 248564 4100 249156 4128
rect 248564 4088 248570 4100
rect 249150 4088 249156 4100
rect 249208 4088 249214 4140
rect 249702 4088 249708 4140
rect 249760 4128 249766 4140
rect 250346 4128 250352 4140
rect 249760 4100 250352 4128
rect 249760 4088 249766 4100
rect 250346 4088 250352 4100
rect 250404 4088 250410 4140
rect 252554 4088 252560 4140
rect 252612 4128 252618 4140
rect 253842 4128 253848 4140
rect 252612 4100 253848 4128
rect 252612 4088 252618 4100
rect 253842 4088 253848 4100
rect 253900 4088 253906 4140
rect 266998 4088 267004 4140
rect 267056 4128 267062 4140
rect 268102 4128 268108 4140
rect 267056 4100 268108 4128
rect 267056 4088 267062 4100
rect 268102 4088 268108 4100
rect 268160 4088 268166 4140
rect 303522 4088 303528 4140
rect 303580 4128 303586 4140
rect 314378 4128 314384 4140
rect 303580 4100 314384 4128
rect 303580 4088 303586 4100
rect 314378 4088 314384 4100
rect 314436 4088 314442 4140
rect 314562 4088 314568 4140
rect 314620 4128 314626 4140
rect 327626 4128 327632 4140
rect 314620 4100 327632 4128
rect 314620 4088 314626 4100
rect 327626 4088 327632 4100
rect 327684 4088 327690 4140
rect 328362 4088 328368 4140
rect 328420 4128 328426 4140
rect 345474 4128 345480 4140
rect 328420 4100 345480 4128
rect 328420 4088 328426 4100
rect 345474 4088 345480 4100
rect 345532 4088 345538 4140
rect 346302 4088 346308 4140
rect 346360 4128 346366 4140
rect 366910 4128 366916 4140
rect 346360 4100 366916 4128
rect 346360 4088 346366 4100
rect 366910 4088 366916 4100
rect 366968 4088 366974 4140
rect 368382 4088 368388 4140
rect 368440 4128 368446 4140
rect 393038 4128 393044 4140
rect 368440 4100 393044 4128
rect 368440 4088 368446 4100
rect 393038 4088 393044 4100
rect 393096 4088 393102 4140
rect 394602 4088 394608 4140
rect 394660 4128 394666 4140
rect 425146 4128 425152 4140
rect 394660 4100 425152 4128
rect 394660 4088 394666 4100
rect 425146 4088 425152 4100
rect 425204 4088 425210 4140
rect 427722 4088 427728 4140
rect 427780 4128 427786 4140
rect 427780 4100 432644 4128
rect 427780 4088 427786 4100
rect 68278 4060 68284 4072
rect 39408 4032 68284 4060
rect 68278 4020 68284 4032
rect 68336 4020 68342 4072
rect 69474 4020 69480 4072
rect 69532 4060 69538 4072
rect 100846 4060 100852 4072
rect 69532 4032 100852 4060
rect 69532 4020 69538 4032
rect 100846 4020 100852 4032
rect 100904 4020 100910 4072
rect 252278 4020 252284 4072
rect 252336 4060 252342 4072
rect 252646 4060 252652 4072
rect 252336 4032 252652 4060
rect 252336 4020 252342 4032
rect 252646 4020 252652 4032
rect 252704 4020 252710 4072
rect 289722 4020 289728 4072
rect 289780 4060 289786 4072
rect 297910 4060 297916 4072
rect 289780 4032 297916 4060
rect 289780 4020 289786 4032
rect 297910 4020 297916 4032
rect 297968 4020 297974 4072
rect 310330 4020 310336 4072
rect 310388 4060 310394 4072
rect 322750 4060 322756 4072
rect 310388 4032 322756 4060
rect 310388 4020 310394 4032
rect 322750 4020 322756 4032
rect 322808 4020 322814 4072
rect 325602 4020 325608 4072
rect 325660 4060 325666 4072
rect 341886 4060 341892 4072
rect 325660 4032 341892 4060
rect 325660 4020 325666 4032
rect 341886 4020 341892 4032
rect 341944 4020 341950 4072
rect 344922 4020 344928 4072
rect 344980 4060 344986 4072
rect 364518 4060 364524 4072
rect 344980 4032 364524 4060
rect 344980 4020 344986 4032
rect 364518 4020 364524 4032
rect 364576 4020 364582 4072
rect 371142 4020 371148 4072
rect 371200 4060 371206 4072
rect 396626 4060 396632 4072
rect 371200 4032 396632 4060
rect 371200 4020 371206 4032
rect 396626 4020 396632 4032
rect 396684 4020 396690 4072
rect 398742 4020 398748 4072
rect 398800 4060 398806 4072
rect 431126 4060 431132 4072
rect 398800 4032 431132 4060
rect 398800 4020 398806 4032
rect 431126 4020 431132 4032
rect 431184 4020 431190 4072
rect 432616 4060 432644 4100
rect 433978 4088 433984 4140
rect 434036 4128 434042 4140
rect 435818 4128 435824 4140
rect 434036 4100 435824 4128
rect 434036 4088 434042 4100
rect 435818 4088 435824 4100
rect 435876 4088 435882 4140
rect 436002 4088 436008 4140
rect 436060 4128 436066 4140
rect 476298 4128 476304 4140
rect 436060 4100 476304 4128
rect 436060 4088 436066 4100
rect 476298 4088 476304 4100
rect 476356 4088 476362 4140
rect 499482 4088 499488 4140
rect 499540 4128 499546 4140
rect 552382 4128 552388 4140
rect 499540 4100 552388 4128
rect 499540 4088 499546 4100
rect 552382 4088 552388 4100
rect 552440 4088 552446 4140
rect 440053 4063 440111 4069
rect 440053 4060 440065 4063
rect 432616 4032 440065 4060
rect 440053 4029 440065 4032
rect 440099 4029 440111 4063
rect 440053 4023 440111 4029
rect 440142 4020 440148 4072
rect 440200 4060 440206 4072
rect 481082 4060 481088 4072
rect 440200 4032 481088 4060
rect 440200 4020 440206 4032
rect 481082 4020 481088 4032
rect 481140 4020 481146 4072
rect 492582 4020 492588 4072
rect 492640 4060 492646 4072
rect 545298 4060 545304 4072
rect 492640 4032 545304 4060
rect 492640 4020 492646 4032
rect 545298 4020 545304 4032
rect 545356 4020 545362 4072
rect 545758 4020 545764 4072
rect 545816 4060 545822 4072
rect 571426 4060 571432 4072
rect 545816 4032 571432 4060
rect 545816 4020 545822 4032
rect 571426 4020 571432 4032
rect 571484 4020 571490 4072
rect 25498 3952 25504 4004
rect 25556 3992 25562 4004
rect 57238 3992 57244 4004
rect 25556 3964 57244 3992
rect 25556 3952 25562 3964
rect 57238 3952 57244 3964
rect 57296 3952 57302 4004
rect 65978 3952 65984 4004
rect 66036 3992 66042 4004
rect 96798 3992 96804 4004
rect 66036 3964 96804 3992
rect 66036 3952 66042 3964
rect 96798 3952 96804 3964
rect 96856 3952 96862 4004
rect 295242 3952 295248 4004
rect 295300 3992 295306 4004
rect 304994 3992 305000 4004
rect 295300 3964 305000 3992
rect 295300 3952 295306 3964
rect 304994 3952 305000 3964
rect 305052 3952 305058 4004
rect 307570 3952 307576 4004
rect 307628 3992 307634 4004
rect 319254 3992 319260 4004
rect 307628 3964 319260 3992
rect 307628 3952 307634 3964
rect 319254 3952 319260 3964
rect 319312 3952 319318 4004
rect 326982 3952 326988 4004
rect 327040 3992 327046 4004
rect 344278 3992 344284 4004
rect 327040 3964 344284 3992
rect 327040 3952 327046 3964
rect 344278 3952 344284 3964
rect 344336 3952 344342 4004
rect 350442 3952 350448 4004
rect 350500 3992 350506 4004
rect 371602 3992 371608 4004
rect 350500 3964 371608 3992
rect 350500 3952 350506 3964
rect 371602 3952 371608 3964
rect 371660 3952 371666 4004
rect 373902 3952 373908 4004
rect 373960 3992 373966 4004
rect 395893 3995 395951 4001
rect 395893 3992 395905 3995
rect 373960 3964 395905 3992
rect 373960 3952 373966 3964
rect 395893 3961 395905 3964
rect 395939 3961 395951 3995
rect 395893 3955 395951 3961
rect 395982 3952 395988 4004
rect 396040 3992 396046 4004
rect 401413 3995 401471 4001
rect 401413 3992 401425 3995
rect 396040 3964 401425 3992
rect 396040 3952 396046 3964
rect 401413 3961 401425 3964
rect 401459 3961 401471 3995
rect 401413 3955 401471 3961
rect 401502 3952 401508 4004
rect 401560 3992 401566 4004
rect 423033 3995 423091 4001
rect 423033 3992 423045 3995
rect 401560 3964 423045 3992
rect 401560 3952 401566 3964
rect 423033 3961 423045 3964
rect 423079 3961 423091 3995
rect 423033 3955 423091 3961
rect 429102 3952 429108 4004
rect 429160 3992 429166 4004
rect 432417 3995 432475 4001
rect 432417 3992 432429 3995
rect 429160 3964 432429 3992
rect 429160 3952 429166 3964
rect 432417 3961 432429 3964
rect 432463 3961 432475 3995
rect 432417 3955 432475 3961
rect 433242 3952 433248 4004
rect 433300 3992 433306 4004
rect 438581 3995 438639 4001
rect 438581 3992 438593 3995
rect 433300 3964 438593 3992
rect 433300 3952 433306 3964
rect 438581 3961 438593 3964
rect 438627 3961 438639 3995
rect 438581 3955 438639 3961
rect 438670 3952 438676 4004
rect 438728 3992 438734 4004
rect 479886 3992 479892 4004
rect 438728 3964 479892 3992
rect 438728 3952 438734 3964
rect 479886 3952 479892 3964
rect 479944 3952 479950 4004
rect 493962 3952 493968 4004
rect 494020 3992 494026 4004
rect 546494 3992 546500 4004
rect 494020 3964 546500 3992
rect 494020 3952 494026 3964
rect 546494 3952 546500 3964
rect 546552 3952 546558 4004
rect 547138 3952 547144 4004
rect 547196 3992 547202 4004
rect 578602 3992 578608 4004
rect 547196 3964 578608 3992
rect 547196 3952 547202 3964
rect 578602 3952 578608 3964
rect 578660 3952 578666 4004
rect 24302 3884 24308 3936
rect 24360 3924 24366 3936
rect 59906 3924 59912 3936
rect 24360 3896 59912 3924
rect 24360 3884 24366 3896
rect 59906 3884 59912 3896
rect 59964 3884 59970 3936
rect 62390 3884 62396 3936
rect 62448 3924 62454 3936
rect 93946 3924 93952 3936
rect 62448 3896 93952 3924
rect 62448 3884 62454 3896
rect 93946 3884 93952 3896
rect 94004 3884 94010 3936
rect 98086 3884 98092 3936
rect 98144 3924 98150 3936
rect 124306 3924 124312 3936
rect 98144 3896 124312 3924
rect 98144 3884 98150 3896
rect 124306 3884 124312 3896
rect 124364 3884 124370 3936
rect 293862 3884 293868 3936
rect 293920 3924 293926 3936
rect 303798 3924 303804 3936
rect 293920 3896 303804 3924
rect 293920 3884 293926 3896
rect 303798 3884 303804 3896
rect 303856 3884 303862 3936
rect 313182 3884 313188 3936
rect 313240 3924 313246 3936
rect 326430 3924 326436 3936
rect 313240 3896 326436 3924
rect 313240 3884 313246 3896
rect 326430 3884 326436 3896
rect 326488 3884 326494 3936
rect 331030 3884 331036 3936
rect 331088 3924 331094 3936
rect 347866 3924 347872 3936
rect 331088 3896 347872 3924
rect 331088 3884 331094 3896
rect 347866 3884 347872 3896
rect 347924 3884 347930 3936
rect 349062 3884 349068 3936
rect 349120 3924 349126 3936
rect 370406 3924 370412 3936
rect 349120 3896 370412 3924
rect 349120 3884 349126 3896
rect 370406 3884 370412 3896
rect 370464 3884 370470 3936
rect 372522 3884 372528 3936
rect 372580 3924 372586 3936
rect 399018 3924 399024 3936
rect 372580 3896 399024 3924
rect 372580 3884 372586 3896
rect 399018 3884 399024 3896
rect 399076 3884 399082 3936
rect 402238 3884 402244 3936
rect 402296 3924 402302 3936
rect 402790 3924 402796 3936
rect 402296 3896 402796 3924
rect 402296 3884 402302 3896
rect 402790 3884 402796 3896
rect 402848 3884 402854 3936
rect 422849 3927 422907 3933
rect 422849 3924 422861 3927
rect 411088 3896 422861 3924
rect 14826 3816 14832 3868
rect 14884 3856 14890 3868
rect 50338 3856 50344 3868
rect 14884 3828 50344 3856
rect 14884 3816 14890 3828
rect 50338 3816 50344 3828
rect 50396 3816 50402 3868
rect 55214 3816 55220 3868
rect 55272 3856 55278 3868
rect 82541 3859 82599 3865
rect 82541 3856 82553 3859
rect 55272 3828 82553 3856
rect 55272 3816 55278 3828
rect 82541 3825 82553 3828
rect 82587 3825 82599 3859
rect 82541 3819 82599 3825
rect 82630 3816 82636 3868
rect 82688 3856 82694 3868
rect 83458 3856 83464 3868
rect 82688 3828 83464 3856
rect 82688 3816 82694 3828
rect 83458 3816 83464 3828
rect 83516 3816 83522 3868
rect 101582 3816 101588 3868
rect 101640 3856 101646 3868
rect 127066 3856 127072 3868
rect 101640 3828 127072 3856
rect 101640 3816 101646 3828
rect 127066 3816 127072 3828
rect 127124 3816 127130 3868
rect 273162 3816 273168 3868
rect 273220 3856 273226 3868
rect 278866 3856 278872 3868
rect 273220 3828 278872 3856
rect 273220 3816 273226 3828
rect 278866 3816 278872 3828
rect 278924 3816 278930 3868
rect 285582 3816 285588 3868
rect 285640 3856 285646 3868
rect 293126 3856 293132 3868
rect 285640 3828 293132 3856
rect 285640 3816 285646 3828
rect 293126 3816 293132 3828
rect 293184 3816 293190 3868
rect 293770 3816 293776 3868
rect 293828 3856 293834 3868
rect 302602 3856 302608 3868
rect 293828 3828 302608 3856
rect 293828 3816 293834 3828
rect 302602 3816 302608 3828
rect 302660 3816 302666 3868
rect 303430 3816 303436 3868
rect 303488 3856 303494 3868
rect 315758 3856 315764 3868
rect 303488 3828 315764 3856
rect 303488 3816 303494 3828
rect 315758 3816 315764 3828
rect 315816 3816 315822 3868
rect 315942 3816 315948 3868
rect 316000 3856 316006 3868
rect 330018 3856 330024 3868
rect 316000 3828 330024 3856
rect 316000 3816 316006 3828
rect 330018 3816 330024 3828
rect 330076 3816 330082 3868
rect 336642 3816 336648 3868
rect 336700 3856 336706 3868
rect 354950 3856 354956 3868
rect 336700 3828 354956 3856
rect 336700 3816 336706 3828
rect 354950 3816 354956 3828
rect 355008 3816 355014 3868
rect 355962 3816 355968 3868
rect 356020 3856 356026 3868
rect 378778 3856 378784 3868
rect 356020 3828 378784 3856
rect 356020 3816 356026 3828
rect 378778 3816 378784 3828
rect 378836 3816 378842 3868
rect 379422 3816 379428 3868
rect 379480 3856 379486 3868
rect 407298 3856 407304 3868
rect 379480 3828 407304 3856
rect 379480 3816 379486 3828
rect 407298 3816 407304 3828
rect 407356 3816 407362 3868
rect 16500 3760 27016 3788
rect 6454 3612 6460 3664
rect 6512 3652 6518 3664
rect 16500 3652 16528 3760
rect 6512 3624 16528 3652
rect 22020 3692 26924 3720
rect 6512 3612 6518 3624
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 22020 3584 22048 3692
rect 2924 3556 22048 3584
rect 26896 3584 26924 3692
rect 26988 3652 27016 3760
rect 39758 3748 39764 3800
rect 39816 3788 39822 3800
rect 76098 3788 76104 3800
rect 39816 3760 76104 3788
rect 39816 3748 39822 3760
rect 76098 3748 76104 3760
rect 76156 3748 76162 3800
rect 79042 3748 79048 3800
rect 79100 3788 79106 3800
rect 79962 3788 79968 3800
rect 79100 3760 79968 3788
rect 79100 3748 79106 3760
rect 79962 3748 79968 3760
rect 80020 3748 80026 3800
rect 80238 3748 80244 3800
rect 80296 3788 80302 3800
rect 109034 3788 109040 3800
rect 80296 3760 109040 3788
rect 80296 3748 80302 3760
rect 109034 3748 109040 3760
rect 109092 3748 109098 3800
rect 277302 3748 277308 3800
rect 277360 3788 277366 3800
rect 282454 3788 282460 3800
rect 277360 3760 282460 3788
rect 277360 3748 277366 3760
rect 282454 3748 282460 3760
rect 282512 3748 282518 3800
rect 284202 3748 284208 3800
rect 284260 3788 284266 3800
rect 291930 3788 291936 3800
rect 284260 3760 291936 3788
rect 284260 3748 284266 3760
rect 291930 3748 291936 3760
rect 291988 3748 291994 3800
rect 292482 3748 292488 3800
rect 292540 3788 292546 3800
rect 301406 3788 301412 3800
rect 292540 3760 301412 3788
rect 292540 3748 292546 3760
rect 301406 3748 301412 3760
rect 301464 3748 301470 3800
rect 302142 3748 302148 3800
rect 302200 3788 302206 3800
rect 313366 3788 313372 3800
rect 302200 3760 313372 3788
rect 302200 3748 302206 3760
rect 313366 3748 313372 3760
rect 313424 3748 313430 3800
rect 314470 3748 314476 3800
rect 314528 3788 314534 3800
rect 328822 3788 328828 3800
rect 314528 3760 328828 3788
rect 314528 3748 314534 3760
rect 328822 3748 328828 3760
rect 328880 3748 328886 3800
rect 335262 3748 335268 3800
rect 335320 3788 335326 3800
rect 353754 3788 353760 3800
rect 335320 3760 353760 3788
rect 335320 3748 335326 3760
rect 353754 3748 353760 3760
rect 353812 3748 353818 3800
rect 354582 3748 354588 3800
rect 354640 3788 354646 3800
rect 377582 3788 377588 3800
rect 354640 3760 377588 3788
rect 354640 3748 354646 3760
rect 377582 3748 377588 3760
rect 377640 3748 377646 3800
rect 378042 3748 378048 3800
rect 378100 3788 378106 3800
rect 406102 3788 406108 3800
rect 378100 3760 406108 3788
rect 378100 3748 378106 3760
rect 406102 3748 406108 3760
rect 406160 3748 406166 3800
rect 408402 3748 408408 3800
rect 408460 3788 408466 3800
rect 411088 3788 411116 3896
rect 422849 3893 422861 3896
rect 422895 3893 422907 3927
rect 422849 3887 422907 3893
rect 422941 3927 422999 3933
rect 422941 3893 422953 3927
rect 422987 3924 422999 3927
rect 431681 3927 431739 3933
rect 431681 3924 431693 3927
rect 422987 3896 431693 3924
rect 422987 3893 422999 3896
rect 422941 3887 422999 3893
rect 431681 3893 431693 3896
rect 431727 3893 431739 3927
rect 431681 3887 431739 3893
rect 432601 3927 432659 3933
rect 432601 3893 432613 3927
rect 432647 3924 432659 3927
rect 441798 3924 441804 3936
rect 432647 3896 441804 3924
rect 432647 3893 432659 3896
rect 432601 3887 432659 3893
rect 441798 3884 441804 3896
rect 441856 3884 441862 3936
rect 443638 3884 443644 3936
rect 443696 3924 443702 3936
rect 449621 3927 449679 3933
rect 449621 3924 449633 3927
rect 443696 3896 449633 3924
rect 443696 3884 443702 3896
rect 449621 3893 449633 3896
rect 449667 3893 449679 3927
rect 449621 3887 449679 3893
rect 449802 3884 449808 3936
rect 449860 3924 449866 3936
rect 451829 3927 451887 3933
rect 451829 3924 451841 3927
rect 449860 3896 451841 3924
rect 449860 3884 449866 3896
rect 451829 3893 451841 3896
rect 451875 3893 451887 3927
rect 451829 3887 451887 3893
rect 451918 3884 451924 3936
rect 451976 3924 451982 3936
rect 453666 3924 453672 3936
rect 451976 3896 453672 3924
rect 451976 3884 451982 3896
rect 453666 3884 453672 3896
rect 453724 3884 453730 3936
rect 453761 3927 453819 3933
rect 453761 3893 453773 3927
rect 453807 3924 453819 3927
rect 457254 3924 457260 3936
rect 453807 3896 457260 3924
rect 453807 3893 453819 3896
rect 453761 3887 453819 3893
rect 457254 3884 457260 3896
rect 457312 3884 457318 3936
rect 457349 3927 457407 3933
rect 457349 3893 457361 3927
rect 457395 3924 457407 3927
rect 495342 3924 495348 3936
rect 457395 3896 495348 3924
rect 457395 3893 457407 3896
rect 457349 3887 457407 3893
rect 495342 3884 495348 3896
rect 495400 3884 495406 3936
rect 508498 3884 508504 3936
rect 508556 3924 508562 3936
rect 510798 3924 510804 3936
rect 508556 3896 510804 3924
rect 508556 3884 508562 3896
rect 510798 3884 510804 3896
rect 510856 3884 510862 3936
rect 514021 3927 514079 3933
rect 514021 3893 514033 3927
rect 514067 3924 514079 3927
rect 559558 3924 559564 3936
rect 514067 3896 559564 3924
rect 514067 3893 514079 3896
rect 514021 3887 514079 3893
rect 559558 3884 559564 3896
rect 559616 3884 559622 3936
rect 411162 3816 411168 3868
rect 411220 3856 411226 3868
rect 445386 3856 445392 3868
rect 411220 3828 445392 3856
rect 411220 3816 411226 3828
rect 445386 3816 445392 3828
rect 445444 3816 445450 3868
rect 445481 3859 445539 3865
rect 445481 3825 445493 3859
rect 445527 3856 445539 3859
rect 452470 3856 452476 3868
rect 445527 3828 452476 3856
rect 445527 3825 445539 3828
rect 445481 3819 445539 3825
rect 452470 3816 452476 3828
rect 452528 3816 452534 3868
rect 491754 3856 491760 3868
rect 452580 3828 491760 3856
rect 408460 3760 411116 3788
rect 408460 3748 408466 3760
rect 416682 3748 416688 3800
rect 416740 3788 416746 3800
rect 422941 3791 422999 3797
rect 422941 3788 422953 3791
rect 416740 3760 422953 3788
rect 416740 3748 416746 3760
rect 422941 3757 422953 3760
rect 422987 3757 422999 3791
rect 422941 3751 422999 3757
rect 423033 3791 423091 3797
rect 423033 3757 423045 3791
rect 423079 3788 423091 3791
rect 431221 3791 431279 3797
rect 431221 3788 431233 3791
rect 423079 3760 431233 3788
rect 423079 3757 423091 3760
rect 423033 3751 423091 3757
rect 431221 3757 431233 3760
rect 431267 3757 431279 3791
rect 431221 3751 431279 3757
rect 431681 3791 431739 3797
rect 431681 3757 431693 3791
rect 431727 3788 431739 3791
rect 437477 3791 437535 3797
rect 437477 3788 437489 3791
rect 431727 3760 437489 3788
rect 431727 3757 431739 3760
rect 431681 3751 431739 3757
rect 437477 3757 437489 3760
rect 437523 3757 437535 3791
rect 437477 3751 437535 3757
rect 449710 3748 449716 3800
rect 449768 3788 449774 3800
rect 452580 3788 452608 3828
rect 491754 3816 491760 3828
rect 491812 3816 491818 3868
rect 501598 3816 501604 3868
rect 501656 3856 501662 3868
rect 501656 3828 506244 3856
rect 501656 3816 501662 3828
rect 449768 3760 452608 3788
rect 452657 3791 452715 3797
rect 449768 3748 449774 3760
rect 452657 3757 452669 3791
rect 452703 3788 452715 3791
rect 452703 3760 453988 3788
rect 452703 3757 452715 3760
rect 452657 3751 452715 3757
rect 27890 3680 27896 3732
rect 27948 3720 27954 3732
rect 28902 3720 28908 3732
rect 27948 3692 28908 3720
rect 27948 3680 27954 3692
rect 28902 3680 28908 3692
rect 28960 3680 28966 3732
rect 32674 3680 32680 3732
rect 32732 3720 32738 3732
rect 70394 3720 70400 3732
rect 32732 3692 70400 3720
rect 32732 3680 32738 3692
rect 70394 3680 70400 3692
rect 70452 3680 70458 3732
rect 76650 3680 76656 3732
rect 76708 3720 76714 3732
rect 106274 3720 106280 3732
rect 76708 3692 106280 3720
rect 76708 3680 76714 3692
rect 106274 3680 106280 3692
rect 106332 3680 106338 3732
rect 115937 3723 115995 3729
rect 115937 3720 115949 3723
rect 106384 3692 115949 3720
rect 40589 3655 40647 3661
rect 40589 3652 40601 3655
rect 26988 3624 40601 3652
rect 40589 3621 40601 3624
rect 40635 3621 40647 3655
rect 45646 3652 45652 3664
rect 40589 3615 40647 3621
rect 40696 3624 45652 3652
rect 40696 3584 40724 3624
rect 45646 3612 45652 3624
rect 45704 3612 45710 3664
rect 56413 3655 56471 3661
rect 56413 3621 56425 3655
rect 56459 3652 56471 3655
rect 56502 3652 56508 3664
rect 56459 3624 56508 3652
rect 56459 3621 56471 3624
rect 56413 3615 56471 3621
rect 56502 3612 56508 3624
rect 56560 3612 56566 3664
rect 58802 3612 58808 3664
rect 58860 3652 58866 3664
rect 91094 3652 91100 3664
rect 58860 3624 91100 3652
rect 58860 3612 58866 3624
rect 91094 3612 91100 3624
rect 91152 3612 91158 3664
rect 94498 3612 94504 3664
rect 94556 3652 94562 3664
rect 106384 3652 106412 3692
rect 115937 3689 115949 3692
rect 115983 3689 115995 3723
rect 115937 3683 115995 3689
rect 121822 3680 121828 3732
rect 121880 3720 121886 3732
rect 122742 3720 122748 3732
rect 121880 3692 122748 3720
rect 121880 3680 121886 3692
rect 122742 3680 122748 3692
rect 122800 3680 122806 3732
rect 227714 3680 227720 3732
rect 227772 3720 227778 3732
rect 230566 3720 230572 3732
rect 227772 3692 230572 3720
rect 227772 3680 227778 3692
rect 230566 3680 230572 3692
rect 230624 3680 230630 3732
rect 267642 3680 267648 3732
rect 267700 3720 267706 3732
rect 271690 3720 271696 3732
rect 267700 3692 271696 3720
rect 267700 3680 267706 3692
rect 271690 3680 271696 3692
rect 271748 3680 271754 3732
rect 300670 3680 300676 3732
rect 300728 3720 300734 3732
rect 312170 3720 312176 3732
rect 300728 3692 312176 3720
rect 300728 3680 300734 3692
rect 312170 3680 312176 3692
rect 312228 3680 312234 3732
rect 317230 3680 317236 3732
rect 317288 3720 317294 3732
rect 331214 3720 331220 3732
rect 317288 3692 331220 3720
rect 317288 3680 317294 3692
rect 331214 3680 331220 3692
rect 331272 3680 331278 3732
rect 333882 3680 333888 3732
rect 333940 3720 333946 3732
rect 352558 3720 352564 3732
rect 333940 3692 352564 3720
rect 333940 3680 333946 3692
rect 352558 3680 352564 3692
rect 352616 3680 352622 3732
rect 358722 3680 358728 3732
rect 358780 3720 358786 3732
rect 381170 3720 381176 3732
rect 358780 3692 381176 3720
rect 358780 3680 358786 3692
rect 381170 3680 381176 3692
rect 381228 3680 381234 3732
rect 382090 3680 382096 3732
rect 382148 3720 382154 3732
rect 410886 3720 410892 3732
rect 382148 3692 410892 3720
rect 382148 3680 382154 3692
rect 410886 3680 410892 3692
rect 410944 3680 410950 3732
rect 413922 3680 413928 3732
rect 413980 3720 413986 3732
rect 448974 3720 448980 3732
rect 413980 3692 448980 3720
rect 413980 3680 413986 3692
rect 448974 3680 448980 3692
rect 449032 3680 449038 3732
rect 449621 3723 449679 3729
rect 449621 3689 449633 3723
rect 449667 3720 449679 3723
rect 451737 3723 451795 3729
rect 451737 3720 451749 3723
rect 449667 3692 451749 3720
rect 449667 3689 449679 3692
rect 449621 3683 449679 3689
rect 451737 3689 451749 3692
rect 451783 3689 451795 3723
rect 453761 3723 453819 3729
rect 453761 3720 453773 3723
rect 451737 3683 451795 3689
rect 451844 3692 453773 3720
rect 94556 3624 106412 3652
rect 94556 3612 94562 3624
rect 123018 3612 123024 3664
rect 123076 3652 123082 3664
rect 124122 3652 124128 3664
rect 123076 3624 124128 3652
rect 123076 3612 123082 3624
rect 124122 3612 124128 3624
rect 124180 3612 124186 3664
rect 275922 3612 275928 3664
rect 275980 3652 275986 3664
rect 281258 3652 281264 3664
rect 275980 3624 281264 3652
rect 275980 3612 275986 3624
rect 281258 3612 281264 3624
rect 281316 3612 281322 3664
rect 284110 3612 284116 3664
rect 284168 3652 284174 3664
rect 290734 3652 290740 3664
rect 284168 3624 290740 3652
rect 284168 3612 284174 3624
rect 290734 3612 290740 3624
rect 290792 3612 290798 3664
rect 291010 3612 291016 3664
rect 291068 3652 291074 3664
rect 300302 3652 300308 3664
rect 291068 3624 300308 3652
rect 291068 3612 291074 3624
rect 300302 3612 300308 3624
rect 300360 3612 300366 3664
rect 300762 3612 300768 3664
rect 300820 3652 300826 3664
rect 310974 3652 310980 3664
rect 300820 3624 310980 3652
rect 300820 3612 300826 3624
rect 310974 3612 310980 3624
rect 311032 3612 311038 3664
rect 311802 3612 311808 3664
rect 311860 3652 311866 3664
rect 325234 3652 325240 3664
rect 311860 3624 325240 3652
rect 311860 3612 311866 3624
rect 325234 3612 325240 3624
rect 325292 3612 325298 3664
rect 326890 3612 326896 3664
rect 326948 3652 326954 3664
rect 343082 3652 343088 3664
rect 326948 3624 343088 3652
rect 326948 3612 326954 3624
rect 343082 3612 343088 3624
rect 343140 3612 343146 3664
rect 343542 3612 343548 3664
rect 343600 3652 343606 3664
rect 363322 3652 363328 3664
rect 343600 3624 363328 3652
rect 343600 3612 343606 3624
rect 363322 3612 363328 3624
rect 363380 3612 363386 3664
rect 364242 3612 364248 3664
rect 364300 3652 364306 3664
rect 388254 3652 388260 3664
rect 364300 3624 388260 3652
rect 364300 3612 364306 3624
rect 388254 3612 388260 3624
rect 388312 3612 388318 3664
rect 390462 3612 390468 3664
rect 390520 3652 390526 3664
rect 420362 3652 420368 3664
rect 390520 3624 420368 3652
rect 390520 3612 390526 3624
rect 420362 3612 420368 3624
rect 420420 3612 420426 3664
rect 420822 3612 420828 3664
rect 420880 3652 420886 3664
rect 451844 3652 451872 3692
rect 453761 3689 453773 3692
rect 453807 3689 453819 3723
rect 453960 3720 453988 3760
rect 455322 3748 455328 3800
rect 455380 3788 455386 3800
rect 498930 3788 498936 3800
rect 455380 3760 498936 3788
rect 455380 3748 455386 3760
rect 498930 3748 498936 3760
rect 498988 3748 498994 3800
rect 499390 3748 499396 3800
rect 499448 3788 499454 3800
rect 506109 3791 506167 3797
rect 506109 3788 506121 3791
rect 499448 3760 506121 3788
rect 499448 3748 499454 3760
rect 506109 3757 506121 3760
rect 506155 3757 506167 3791
rect 506109 3751 506167 3757
rect 492950 3720 492956 3732
rect 453960 3692 492956 3720
rect 453761 3683 453819 3689
rect 492950 3680 492956 3692
rect 493008 3680 493014 3732
rect 494698 3680 494704 3732
rect 494756 3720 494762 3732
rect 496538 3720 496544 3732
rect 494756 3692 496544 3720
rect 494756 3680 494762 3692
rect 496538 3680 496544 3692
rect 496596 3680 496602 3732
rect 502426 3680 502432 3732
rect 502484 3720 502490 3732
rect 503622 3720 503628 3732
rect 502484 3692 503628 3720
rect 502484 3680 502490 3692
rect 503622 3680 503628 3692
rect 503680 3680 503686 3732
rect 505002 3680 505008 3732
rect 505060 3720 505066 3732
rect 506216 3720 506244 3828
rect 506382 3816 506388 3868
rect 506440 3856 506446 3868
rect 560754 3856 560760 3868
rect 506440 3828 560760 3856
rect 506440 3816 506446 3828
rect 560754 3816 560760 3828
rect 560812 3816 560818 3868
rect 506293 3791 506351 3797
rect 506293 3757 506305 3791
rect 506339 3788 506351 3791
rect 553578 3788 553584 3800
rect 506339 3760 553584 3788
rect 506339 3757 506351 3760
rect 506293 3751 506351 3757
rect 553578 3748 553584 3760
rect 553636 3748 553642 3800
rect 509602 3720 509608 3732
rect 505060 3692 506152 3720
rect 506216 3692 509608 3720
rect 505060 3680 505066 3692
rect 420880 3624 451872 3652
rect 451921 3655 451979 3661
rect 420880 3612 420886 3624
rect 451921 3621 451933 3655
rect 451967 3652 451979 3655
rect 459554 3652 459560 3664
rect 451967 3624 459560 3652
rect 451967 3621 451979 3624
rect 451921 3615 451979 3621
rect 459554 3612 459560 3624
rect 459612 3612 459618 3664
rect 502334 3652 502340 3664
rect 459664 3624 502340 3652
rect 46198 3584 46204 3596
rect 26896 3556 40724 3584
rect 40788 3556 46204 3584
rect 2924 3544 2930 3556
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 40589 3519 40647 3525
rect 624 3488 39436 3516
rect 624 3476 630 3488
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 39408 3448 39436 3488
rect 40589 3485 40601 3519
rect 40635 3516 40647 3519
rect 40788 3516 40816 3556
rect 46198 3544 46204 3556
rect 46256 3544 46262 3596
rect 46934 3544 46940 3596
rect 46992 3584 46998 3596
rect 75181 3587 75239 3593
rect 75181 3584 75193 3587
rect 46992 3556 75193 3584
rect 46992 3544 46998 3556
rect 75181 3553 75193 3556
rect 75227 3553 75239 3587
rect 82449 3587 82507 3593
rect 82449 3584 82461 3587
rect 75181 3547 75239 3553
rect 75288 3556 82461 3584
rect 40635 3488 40816 3516
rect 40635 3485 40647 3488
rect 40589 3479 40647 3485
rect 43346 3476 43352 3528
rect 43404 3516 43410 3528
rect 44082 3516 44088 3528
rect 43404 3488 44088 3516
rect 43404 3476 43410 3488
rect 44082 3476 44088 3488
rect 44140 3476 44146 3528
rect 44542 3476 44548 3528
rect 44600 3516 44606 3528
rect 45462 3516 45468 3528
rect 44600 3488 45468 3516
rect 44600 3476 44606 3488
rect 45462 3476 45468 3488
rect 45520 3476 45526 3528
rect 45738 3476 45744 3528
rect 45796 3516 45802 3528
rect 46842 3516 46848 3528
rect 45796 3488 46848 3516
rect 45796 3476 45802 3488
rect 46842 3476 46848 3488
rect 46900 3476 46906 3528
rect 50522 3476 50528 3528
rect 50580 3516 50586 3528
rect 50982 3516 50988 3528
rect 50580 3488 50988 3516
rect 50580 3476 50586 3488
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 51626 3476 51632 3528
rect 51684 3516 51690 3528
rect 75288 3516 75316 3556
rect 82449 3553 82461 3556
rect 82495 3553 82507 3587
rect 82449 3547 82507 3553
rect 82541 3587 82599 3593
rect 82541 3553 82553 3587
rect 82587 3584 82599 3587
rect 88334 3584 88340 3596
rect 82587 3556 88340 3584
rect 82587 3553 82599 3556
rect 82541 3547 82599 3553
rect 88334 3544 88340 3556
rect 88392 3544 88398 3596
rect 89714 3544 89720 3596
rect 89772 3584 89778 3596
rect 91002 3584 91008 3596
rect 89772 3556 91008 3584
rect 89772 3544 89778 3556
rect 91002 3544 91008 3556
rect 91060 3544 91066 3596
rect 117682 3584 117688 3596
rect 91112 3556 117688 3584
rect 51684 3488 75316 3516
rect 51684 3476 51690 3488
rect 90910 3476 90916 3528
rect 90968 3516 90974 3528
rect 91112 3516 91140 3556
rect 117682 3544 117688 3556
rect 117740 3544 117746 3596
rect 150434 3544 150440 3596
rect 150492 3584 150498 3596
rect 151630 3584 151636 3596
rect 150492 3556 151636 3584
rect 150492 3544 150498 3556
rect 151630 3544 151636 3556
rect 151688 3544 151694 3596
rect 158714 3544 158720 3596
rect 158772 3584 158778 3596
rect 159910 3584 159916 3596
rect 158772 3556 159916 3584
rect 158772 3544 158778 3556
rect 159910 3544 159916 3556
rect 159968 3544 159974 3596
rect 183738 3544 183744 3596
rect 183796 3584 183802 3596
rect 184842 3584 184848 3596
rect 183796 3556 184848 3584
rect 183796 3544 183802 3556
rect 184842 3544 184848 3556
rect 184900 3544 184906 3596
rect 201494 3544 201500 3596
rect 201552 3584 201558 3596
rect 202690 3584 202696 3596
rect 201552 3556 202696 3584
rect 201552 3544 201558 3556
rect 202690 3544 202696 3556
rect 202748 3544 202754 3596
rect 235994 3544 236000 3596
rect 236052 3584 236058 3596
rect 237374 3584 237380 3596
rect 236052 3556 237380 3584
rect 236052 3544 236058 3556
rect 237374 3544 237380 3556
rect 237432 3544 237438 3596
rect 263502 3544 263508 3596
rect 263560 3584 263566 3596
rect 266998 3584 267004 3596
rect 263560 3556 267004 3584
rect 263560 3544 263566 3556
rect 266998 3544 267004 3556
rect 267056 3544 267062 3596
rect 270402 3544 270408 3596
rect 270460 3584 270466 3596
rect 274082 3584 274088 3596
rect 270460 3556 274088 3584
rect 270460 3544 270466 3556
rect 274082 3544 274088 3556
rect 274140 3544 274146 3596
rect 279970 3544 279976 3596
rect 280028 3584 280034 3596
rect 280028 3556 286088 3584
rect 280028 3544 280034 3556
rect 114646 3516 114652 3528
rect 90968 3488 91140 3516
rect 91204 3488 114652 3516
rect 90968 3476 90974 3488
rect 42886 3448 42892 3460
rect 1728 3420 35940 3448
rect 39408 3420 42892 3448
rect 1728 3408 1734 3420
rect 8846 3340 8852 3392
rect 8904 3380 8910 3392
rect 9582 3380 9588 3392
rect 8904 3352 9588 3380
rect 8904 3340 8910 3352
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 10042 3340 10048 3392
rect 10100 3380 10106 3392
rect 10962 3380 10968 3392
rect 10100 3352 10968 3380
rect 10100 3340 10106 3352
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11238 3340 11244 3392
rect 11296 3380 11302 3392
rect 12342 3380 12348 3392
rect 11296 3352 12348 3380
rect 11296 3340 11302 3352
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 34974 3340 34980 3392
rect 35032 3380 35038 3392
rect 35802 3380 35808 3392
rect 35032 3352 35808 3380
rect 35032 3340 35038 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 35912 3244 35940 3420
rect 42886 3408 42892 3420
rect 42944 3408 42950 3460
rect 52822 3408 52828 3460
rect 52880 3448 52886 3460
rect 53742 3448 53748 3460
rect 52880 3420 53748 3448
rect 52880 3408 52886 3420
rect 53742 3408 53748 3420
rect 53800 3408 53806 3460
rect 61194 3408 61200 3460
rect 61252 3448 61258 3460
rect 62022 3448 62028 3460
rect 61252 3420 62028 3448
rect 61252 3408 61258 3420
rect 62022 3408 62028 3420
rect 62080 3408 62086 3460
rect 63586 3408 63592 3460
rect 63644 3448 63650 3460
rect 64782 3448 64788 3460
rect 63644 3420 64788 3448
rect 63644 3408 63650 3420
rect 64782 3408 64788 3420
rect 64840 3408 64846 3460
rect 68278 3408 68284 3460
rect 68336 3448 68342 3460
rect 68922 3448 68928 3460
rect 68336 3420 68928 3448
rect 68336 3408 68342 3420
rect 68922 3408 68928 3420
rect 68980 3408 68986 3460
rect 81434 3408 81440 3460
rect 81492 3448 81498 3460
rect 82722 3448 82728 3460
rect 81492 3420 82728 3448
rect 81492 3408 81498 3420
rect 82722 3408 82728 3420
rect 82780 3408 82786 3460
rect 91204 3448 91232 3488
rect 114646 3476 114652 3488
rect 114704 3476 114710 3528
rect 114738 3476 114744 3528
rect 114796 3516 114802 3528
rect 115842 3516 115848 3528
rect 114796 3488 115848 3516
rect 114796 3476 114802 3488
rect 115842 3476 115848 3488
rect 115900 3476 115906 3528
rect 130194 3476 130200 3528
rect 130252 3516 130258 3528
rect 131022 3516 131028 3528
rect 130252 3488 131028 3516
rect 130252 3476 130258 3488
rect 131022 3476 131028 3488
rect 131080 3476 131086 3528
rect 131390 3476 131396 3528
rect 131448 3516 131454 3528
rect 132402 3516 132408 3528
rect 131448 3488 132408 3516
rect 131448 3476 131454 3488
rect 132402 3476 132408 3488
rect 132460 3476 132466 3528
rect 132586 3476 132592 3528
rect 132644 3516 132650 3528
rect 133690 3516 133696 3528
rect 132644 3488 133696 3516
rect 132644 3476 132650 3488
rect 133690 3476 133696 3488
rect 133748 3476 133754 3528
rect 137278 3476 137284 3528
rect 137336 3516 137342 3528
rect 137922 3516 137928 3528
rect 137336 3488 137928 3516
rect 137336 3476 137342 3488
rect 137922 3476 137928 3488
rect 137980 3476 137986 3528
rect 138474 3476 138480 3528
rect 138532 3516 138538 3528
rect 139302 3516 139308 3528
rect 138532 3488 139308 3516
rect 138532 3476 138538 3488
rect 139302 3476 139308 3488
rect 139360 3476 139366 3528
rect 139670 3476 139676 3528
rect 139728 3516 139734 3528
rect 140682 3516 140688 3528
rect 139728 3488 140688 3516
rect 139728 3476 139734 3488
rect 140682 3476 140688 3488
rect 140740 3476 140746 3528
rect 140866 3476 140872 3528
rect 140924 3516 140930 3528
rect 141970 3516 141976 3528
rect 140924 3488 141976 3516
rect 140924 3476 140930 3488
rect 141970 3476 141976 3488
rect 142028 3476 142034 3528
rect 145650 3476 145656 3528
rect 145708 3516 145714 3528
rect 146202 3516 146208 3528
rect 145708 3488 146208 3516
rect 145708 3476 145714 3488
rect 146202 3476 146208 3488
rect 146260 3476 146266 3528
rect 146846 3476 146852 3528
rect 146904 3516 146910 3528
rect 147582 3516 147588 3528
rect 146904 3488 147588 3516
rect 146904 3476 146910 3488
rect 147582 3476 147588 3488
rect 147640 3476 147646 3528
rect 148042 3476 148048 3528
rect 148100 3516 148106 3528
rect 148962 3516 148968 3528
rect 148100 3488 148968 3516
rect 148100 3476 148106 3488
rect 148962 3476 148968 3488
rect 149020 3476 149026 3528
rect 149238 3476 149244 3528
rect 149296 3516 149302 3528
rect 150342 3516 150348 3528
rect 149296 3488 150348 3516
rect 149296 3476 149302 3488
rect 150342 3476 150348 3488
rect 150400 3476 150406 3528
rect 153930 3476 153936 3528
rect 153988 3516 153994 3528
rect 154482 3516 154488 3528
rect 153988 3488 154488 3516
rect 153988 3476 153994 3488
rect 154482 3476 154488 3488
rect 154540 3476 154546 3528
rect 155126 3476 155132 3528
rect 155184 3516 155190 3528
rect 155862 3516 155868 3528
rect 155184 3488 155868 3516
rect 155184 3476 155190 3488
rect 155862 3476 155868 3488
rect 155920 3476 155926 3528
rect 156322 3476 156328 3528
rect 156380 3516 156386 3528
rect 157242 3516 157248 3528
rect 156380 3488 157248 3516
rect 156380 3476 156386 3488
rect 157242 3476 157248 3488
rect 157300 3476 157306 3528
rect 162302 3476 162308 3528
rect 162360 3516 162366 3528
rect 162762 3516 162768 3528
rect 162360 3488 162768 3516
rect 162360 3476 162366 3488
rect 162762 3476 162768 3488
rect 162820 3476 162826 3528
rect 163498 3476 163504 3528
rect 163556 3516 163562 3528
rect 164142 3516 164148 3528
rect 163556 3488 164148 3516
rect 163556 3476 163562 3488
rect 164142 3476 164148 3488
rect 164200 3476 164206 3528
rect 165890 3476 165896 3528
rect 165948 3516 165954 3528
rect 166902 3516 166908 3528
rect 165948 3488 166908 3516
rect 165948 3476 165954 3488
rect 166902 3476 166908 3488
rect 166960 3476 166966 3528
rect 172974 3476 172980 3528
rect 173032 3516 173038 3528
rect 173802 3516 173808 3528
rect 173032 3488 173808 3516
rect 173032 3476 173038 3488
rect 173802 3476 173808 3488
rect 173860 3476 173866 3528
rect 180150 3476 180156 3528
rect 180208 3516 180214 3528
rect 180702 3516 180708 3528
rect 180208 3488 180708 3516
rect 180208 3476 180214 3488
rect 180702 3476 180708 3488
rect 180760 3476 180766 3528
rect 182542 3476 182548 3528
rect 182600 3516 182606 3528
rect 183462 3516 183468 3528
rect 182600 3488 183468 3516
rect 182600 3476 182606 3488
rect 183462 3476 183468 3488
rect 183520 3476 183526 3528
rect 188430 3476 188436 3528
rect 188488 3516 188494 3528
rect 188982 3516 188988 3528
rect 188488 3488 188988 3516
rect 188488 3476 188494 3488
rect 188982 3476 188988 3488
rect 189040 3476 189046 3528
rect 189626 3476 189632 3528
rect 189684 3516 189690 3528
rect 190362 3516 190368 3528
rect 189684 3488 190368 3516
rect 189684 3476 189690 3488
rect 190362 3476 190368 3488
rect 190420 3476 190426 3528
rect 192018 3476 192024 3528
rect 192076 3516 192082 3528
rect 193122 3516 193128 3528
rect 192076 3488 193128 3516
rect 192076 3476 192082 3488
rect 193122 3476 193128 3488
rect 193180 3476 193186 3528
rect 193214 3476 193220 3528
rect 193272 3516 193278 3528
rect 194502 3516 194508 3528
rect 193272 3488 194508 3516
rect 193272 3476 193278 3488
rect 194502 3476 194508 3488
rect 194560 3476 194566 3528
rect 196802 3476 196808 3528
rect 196860 3516 196866 3528
rect 197262 3516 197268 3528
rect 196860 3488 197268 3516
rect 196860 3476 196866 3488
rect 197262 3476 197268 3488
rect 197320 3476 197326 3528
rect 197998 3476 198004 3528
rect 198056 3516 198062 3528
rect 198642 3516 198648 3528
rect 198056 3488 198648 3516
rect 198056 3476 198062 3488
rect 198642 3476 198648 3488
rect 198700 3476 198706 3528
rect 199194 3476 199200 3528
rect 199252 3516 199258 3528
rect 200022 3516 200028 3528
rect 199252 3488 200028 3516
rect 199252 3476 199258 3488
rect 200022 3476 200028 3488
rect 200080 3476 200086 3528
rect 200390 3476 200396 3528
rect 200448 3516 200454 3528
rect 201402 3516 201408 3528
rect 200448 3488 201408 3516
rect 200448 3476 200454 3488
rect 201402 3476 201408 3488
rect 201460 3476 201466 3528
rect 205082 3476 205088 3528
rect 205140 3516 205146 3528
rect 205542 3516 205548 3528
rect 205140 3488 205548 3516
rect 205140 3476 205146 3488
rect 205542 3476 205548 3488
rect 205600 3476 205606 3528
rect 207474 3476 207480 3528
rect 207532 3516 207538 3528
rect 208302 3516 208308 3528
rect 207532 3488 208308 3516
rect 207532 3476 207538 3488
rect 208302 3476 208308 3488
rect 208360 3476 208366 3528
rect 208670 3476 208676 3528
rect 208728 3516 208734 3528
rect 209682 3516 209688 3528
rect 208728 3488 209688 3516
rect 208728 3476 208734 3488
rect 209682 3476 209688 3488
rect 209740 3476 209746 3528
rect 209866 3476 209872 3528
rect 209924 3516 209930 3528
rect 210970 3516 210976 3528
rect 209924 3488 210976 3516
rect 209924 3476 209930 3488
rect 210970 3476 210976 3488
rect 211028 3476 211034 3528
rect 214650 3476 214656 3528
rect 214708 3516 214714 3528
rect 215202 3516 215208 3528
rect 214708 3488 215208 3516
rect 214708 3476 214714 3488
rect 215202 3476 215208 3488
rect 215260 3476 215266 3528
rect 215846 3476 215852 3528
rect 215904 3516 215910 3528
rect 216582 3516 216588 3528
rect 215904 3488 216588 3516
rect 215904 3476 215910 3488
rect 216582 3476 216588 3488
rect 216640 3476 216646 3528
rect 217042 3476 217048 3528
rect 217100 3516 217106 3528
rect 217962 3516 217968 3528
rect 217100 3488 217968 3516
rect 217100 3476 217106 3488
rect 217962 3476 217968 3488
rect 218020 3476 218026 3528
rect 222930 3476 222936 3528
rect 222988 3516 222994 3528
rect 223482 3516 223488 3528
rect 222988 3488 223488 3516
rect 222988 3476 222994 3488
rect 223482 3476 223488 3488
rect 223540 3476 223546 3528
rect 224126 3476 224132 3528
rect 224184 3516 224190 3528
rect 224862 3516 224868 3528
rect 224184 3488 224868 3516
rect 224184 3476 224190 3488
rect 224862 3476 224868 3488
rect 224920 3476 224926 3528
rect 225322 3476 225328 3528
rect 225380 3516 225386 3528
rect 226242 3516 226248 3528
rect 225380 3488 226248 3516
rect 225380 3476 225386 3488
rect 226242 3476 226248 3488
rect 226300 3476 226306 3528
rect 231302 3476 231308 3528
rect 231360 3516 231366 3528
rect 231762 3516 231768 3528
rect 231360 3488 231768 3516
rect 231360 3476 231366 3488
rect 231762 3476 231768 3488
rect 231820 3476 231826 3528
rect 232498 3476 232504 3528
rect 232556 3516 232562 3528
rect 233142 3516 233148 3528
rect 232556 3488 233148 3516
rect 232556 3476 232562 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 233694 3476 233700 3528
rect 233752 3516 233758 3528
rect 234522 3516 234528 3528
rect 233752 3488 234528 3516
rect 233752 3476 233758 3488
rect 234522 3476 234528 3488
rect 234580 3476 234586 3528
rect 234798 3476 234804 3528
rect 234856 3516 234862 3528
rect 236178 3516 236184 3528
rect 234856 3488 236184 3516
rect 234856 3476 234862 3488
rect 236178 3476 236184 3488
rect 236236 3476 236242 3528
rect 239582 3476 239588 3528
rect 239640 3516 239646 3528
rect 240042 3516 240048 3528
rect 239640 3488 240048 3516
rect 239640 3476 239646 3488
rect 240042 3476 240048 3488
rect 240100 3476 240106 3528
rect 255222 3476 255228 3528
rect 255280 3516 255286 3528
rect 256234 3516 256240 3528
rect 255280 3488 256240 3516
rect 255280 3476 255286 3488
rect 256234 3476 256240 3488
rect 256292 3476 256298 3528
rect 258718 3476 258724 3528
rect 258776 3516 258782 3528
rect 259822 3516 259828 3528
rect 258776 3488 259828 3516
rect 258776 3476 258782 3488
rect 259822 3476 259828 3488
rect 259880 3476 259886 3528
rect 261478 3476 261484 3528
rect 261536 3516 261542 3528
rect 262214 3516 262220 3528
rect 261536 3488 262220 3516
rect 261536 3476 261542 3488
rect 262214 3476 262220 3488
rect 262272 3476 262278 3528
rect 263410 3476 263416 3528
rect 263468 3516 263474 3528
rect 265802 3516 265808 3528
rect 263468 3488 265808 3516
rect 263468 3476 263474 3488
rect 265802 3476 265808 3488
rect 265860 3476 265866 3528
rect 266262 3476 266268 3528
rect 266320 3516 266326 3528
rect 270494 3516 270500 3528
rect 266320 3488 270500 3516
rect 266320 3476 266326 3488
rect 270494 3476 270500 3488
rect 270552 3476 270558 3528
rect 280062 3476 280068 3528
rect 280120 3516 280126 3528
rect 285950 3516 285956 3528
rect 280120 3488 285956 3516
rect 280120 3476 280126 3488
rect 285950 3476 285956 3488
rect 286008 3476 286014 3528
rect 286060 3516 286088 3556
rect 286870 3544 286876 3596
rect 286928 3584 286934 3596
rect 294322 3584 294328 3596
rect 286928 3556 294328 3584
rect 286928 3544 286934 3556
rect 294322 3544 294328 3556
rect 294380 3544 294386 3596
rect 298002 3544 298008 3596
rect 298060 3584 298066 3596
rect 308582 3584 308588 3596
rect 298060 3556 308588 3584
rect 298060 3544 298066 3556
rect 308582 3544 308588 3556
rect 308640 3544 308646 3596
rect 309042 3544 309048 3596
rect 309100 3584 309106 3596
rect 321646 3584 321652 3596
rect 309100 3556 321652 3584
rect 309100 3544 309106 3556
rect 321646 3544 321652 3556
rect 321704 3544 321710 3596
rect 322842 3544 322848 3596
rect 322900 3584 322906 3596
rect 338298 3584 338304 3596
rect 322900 3556 338304 3584
rect 322900 3544 322906 3556
rect 338298 3544 338304 3556
rect 338356 3544 338362 3596
rect 339402 3544 339408 3596
rect 339460 3584 339466 3596
rect 358538 3584 358544 3596
rect 339460 3556 358544 3584
rect 339460 3544 339466 3556
rect 358538 3544 358544 3556
rect 358596 3544 358602 3596
rect 361390 3544 361396 3596
rect 361448 3584 361454 3596
rect 385862 3584 385868 3596
rect 361448 3556 385868 3584
rect 361448 3544 361454 3556
rect 385862 3544 385868 3556
rect 385920 3544 385926 3596
rect 387702 3544 387708 3596
rect 387760 3584 387766 3596
rect 416866 3584 416872 3596
rect 387760 3556 416872 3584
rect 387760 3544 387766 3556
rect 416866 3544 416872 3556
rect 416924 3544 416930 3596
rect 419442 3544 419448 3596
rect 419500 3584 419506 3596
rect 456058 3584 456064 3596
rect 419500 3556 456064 3584
rect 419500 3544 419506 3556
rect 456058 3544 456064 3556
rect 456116 3544 456122 3596
rect 458082 3544 458088 3596
rect 458140 3584 458146 3596
rect 459664 3584 459692 3624
rect 502334 3612 502340 3624
rect 502392 3612 502398 3664
rect 506014 3652 506020 3664
rect 502444 3624 506020 3652
rect 458140 3556 459692 3584
rect 458140 3544 458146 3556
rect 460842 3544 460848 3596
rect 460900 3584 460906 3596
rect 502444 3584 502472 3624
rect 506014 3612 506020 3624
rect 506072 3612 506078 3664
rect 506124 3652 506152 3692
rect 509602 3680 509608 3692
rect 509660 3680 509666 3732
rect 511902 3680 511908 3732
rect 511960 3720 511966 3732
rect 518161 3723 518219 3729
rect 511960 3692 518112 3720
rect 511960 3680 511966 3692
rect 514021 3655 514079 3661
rect 514021 3652 514033 3655
rect 506124 3624 514033 3652
rect 514021 3621 514033 3624
rect 514067 3621 514079 3655
rect 514021 3615 514079 3621
rect 516042 3612 516048 3664
rect 516100 3652 516106 3664
rect 518084 3652 518112 3692
rect 518161 3689 518173 3723
rect 518207 3720 518219 3723
rect 566734 3720 566740 3732
rect 518207 3692 566740 3720
rect 518207 3689 518219 3692
rect 518161 3683 518219 3689
rect 566734 3680 566740 3692
rect 566792 3680 566798 3732
rect 567838 3652 567844 3664
rect 516100 3624 518020 3652
rect 518084 3624 567844 3652
rect 516100 3612 516106 3624
rect 460900 3556 502472 3584
rect 511077 3587 511135 3593
rect 460900 3544 460906 3556
rect 511077 3553 511089 3587
rect 511123 3584 511135 3587
rect 517882 3584 517888 3596
rect 511123 3556 517888 3584
rect 511123 3553 511135 3556
rect 511077 3547 511135 3553
rect 517882 3544 517888 3556
rect 517940 3544 517946 3596
rect 517992 3584 518020 3624
rect 567838 3612 567844 3624
rect 567896 3612 567902 3664
rect 573818 3584 573824 3596
rect 517992 3556 573824 3584
rect 573818 3544 573824 3556
rect 573876 3544 573882 3596
rect 287146 3516 287152 3528
rect 286060 3488 287152 3516
rect 287146 3476 287152 3488
rect 287204 3476 287210 3528
rect 288342 3476 288348 3528
rect 288400 3516 288406 3528
rect 296714 3516 296720 3528
rect 288400 3488 296720 3516
rect 288400 3476 288406 3488
rect 296714 3476 296720 3488
rect 296772 3476 296778 3528
rect 299382 3476 299388 3528
rect 299440 3516 299446 3528
rect 309778 3516 309784 3528
rect 299440 3488 309784 3516
rect 299440 3476 299446 3488
rect 309778 3476 309784 3488
rect 309836 3476 309842 3528
rect 310422 3476 310428 3528
rect 310480 3516 310486 3528
rect 324038 3516 324044 3528
rect 310480 3488 324044 3516
rect 310480 3476 310486 3488
rect 324038 3476 324044 3488
rect 324096 3476 324102 3528
rect 324130 3476 324136 3528
rect 324188 3516 324194 3528
rect 340690 3516 340696 3528
rect 324188 3488 340696 3516
rect 324188 3476 324194 3488
rect 340690 3476 340696 3488
rect 340748 3476 340754 3528
rect 340782 3476 340788 3528
rect 340840 3516 340846 3528
rect 360930 3516 360936 3528
rect 340840 3488 360936 3516
rect 340840 3476 340846 3488
rect 360930 3476 360936 3488
rect 360988 3476 360994 3528
rect 364150 3476 364156 3528
rect 364208 3516 364214 3528
rect 389450 3516 389456 3528
rect 364208 3488 389456 3516
rect 364208 3476 364214 3488
rect 389450 3476 389456 3488
rect 389508 3476 389514 3528
rect 393222 3476 393228 3528
rect 393280 3516 393286 3528
rect 423950 3516 423956 3528
rect 393280 3488 423956 3516
rect 393280 3476 393286 3488
rect 423950 3476 423956 3488
rect 424008 3476 424014 3528
rect 424962 3476 424968 3528
rect 425020 3516 425026 3528
rect 425020 3488 461900 3516
rect 425020 3476 425026 3488
rect 89824 3420 91232 3448
rect 94332 3420 104204 3448
rect 48130 3340 48136 3392
rect 48188 3380 48194 3392
rect 82998 3380 83004 3392
rect 48188 3352 83004 3380
rect 48188 3340 48194 3352
rect 82998 3340 83004 3352
rect 83056 3340 83062 3392
rect 85666 3380 85672 3392
rect 83108 3352 85672 3380
rect 42150 3272 42156 3324
rect 42208 3312 42214 3324
rect 42702 3312 42708 3324
rect 42208 3284 42708 3312
rect 42208 3272 42214 3284
rect 42702 3272 42708 3284
rect 42760 3272 42766 3324
rect 82449 3315 82507 3321
rect 82449 3281 82461 3315
rect 82495 3312 82507 3315
rect 83108 3312 83136 3352
rect 85666 3340 85672 3352
rect 85724 3340 85730 3392
rect 87322 3340 87328 3392
rect 87380 3380 87386 3392
rect 89824 3380 89852 3420
rect 87380 3352 89852 3380
rect 87380 3340 87386 3352
rect 82495 3284 83136 3312
rect 82495 3281 82507 3284
rect 82449 3275 82507 3281
rect 83826 3272 83832 3324
rect 83884 3312 83890 3324
rect 94332 3312 94360 3420
rect 104176 3380 104204 3420
rect 105170 3408 105176 3460
rect 105228 3448 105234 3460
rect 106182 3448 106188 3460
rect 105228 3420 106188 3448
rect 105228 3408 105234 3420
rect 106182 3408 106188 3420
rect 106240 3408 106246 3460
rect 126606 3408 126612 3460
rect 126664 3448 126670 3460
rect 147766 3448 147772 3460
rect 126664 3420 147772 3448
rect 126664 3408 126670 3420
rect 147766 3408 147772 3420
rect 147824 3408 147830 3460
rect 164694 3408 164700 3460
rect 164752 3448 164758 3460
rect 165522 3448 165528 3460
rect 164752 3420 165528 3448
rect 164752 3408 164758 3420
rect 165522 3408 165528 3420
rect 165580 3408 165586 3460
rect 259362 3408 259368 3460
rect 259420 3448 259426 3460
rect 261018 3448 261024 3460
rect 259420 3420 261024 3448
rect 259420 3408 259426 3420
rect 261018 3408 261024 3420
rect 261076 3408 261082 3460
rect 266170 3408 266176 3460
rect 266228 3448 266234 3460
rect 269298 3448 269304 3460
rect 266228 3420 269304 3448
rect 266228 3408 266234 3420
rect 269298 3408 269304 3420
rect 269356 3408 269362 3460
rect 270310 3408 270316 3460
rect 270368 3448 270374 3460
rect 275278 3448 275284 3460
rect 270368 3420 275284 3448
rect 270368 3408 270374 3420
rect 275278 3408 275284 3420
rect 275336 3408 275342 3460
rect 277210 3408 277216 3460
rect 277268 3448 277274 3460
rect 283650 3448 283656 3460
rect 277268 3420 283656 3448
rect 277268 3408 277274 3420
rect 283650 3408 283656 3420
rect 283708 3408 283714 3460
rect 286962 3408 286968 3460
rect 287020 3448 287026 3460
rect 295518 3448 295524 3460
rect 287020 3420 295524 3448
rect 287020 3408 287026 3420
rect 295518 3408 295524 3420
rect 295576 3408 295582 3460
rect 296622 3408 296628 3460
rect 296680 3448 296686 3460
rect 307386 3448 307392 3460
rect 296680 3420 307392 3448
rect 296680 3408 296686 3420
rect 307386 3408 307392 3420
rect 307444 3408 307450 3460
rect 307662 3408 307668 3460
rect 307720 3448 307726 3460
rect 320450 3448 320456 3460
rect 307720 3420 320456 3448
rect 307720 3408 307726 3420
rect 320450 3408 320456 3420
rect 320508 3408 320514 3460
rect 321370 3408 321376 3460
rect 321428 3448 321434 3460
rect 337102 3448 337108 3460
rect 321428 3420 337108 3448
rect 321428 3408 321434 3420
rect 337102 3408 337108 3420
rect 337160 3408 337166 3460
rect 337930 3408 337936 3460
rect 337988 3448 337994 3460
rect 357342 3448 357348 3460
rect 337988 3420 357348 3448
rect 337988 3408 337994 3420
rect 357342 3408 357348 3420
rect 357400 3408 357406 3460
rect 358630 3408 358636 3460
rect 358688 3448 358694 3460
rect 382366 3448 382372 3460
rect 358688 3420 382372 3448
rect 358688 3408 358694 3420
rect 382366 3408 382372 3420
rect 382424 3408 382430 3460
rect 384850 3408 384856 3460
rect 384908 3448 384914 3460
rect 414474 3448 414480 3460
rect 384908 3420 414480 3448
rect 384908 3408 384914 3420
rect 414474 3408 414480 3420
rect 414532 3408 414538 3460
rect 422202 3408 422208 3460
rect 422260 3448 422266 3460
rect 451921 3451 451979 3457
rect 451921 3448 451933 3451
rect 422260 3420 451933 3448
rect 422260 3408 422266 3420
rect 451921 3417 451933 3420
rect 451967 3417 451979 3451
rect 451921 3411 451979 3417
rect 452562 3408 452568 3460
rect 452620 3448 452626 3460
rect 457349 3451 457407 3457
rect 457349 3448 457361 3451
rect 452620 3420 457361 3448
rect 452620 3408 452626 3420
rect 457349 3417 457361 3420
rect 457395 3417 457407 3451
rect 457349 3411 457407 3417
rect 459646 3408 459652 3460
rect 459704 3448 459710 3460
rect 460842 3448 460848 3460
rect 459704 3420 460848 3448
rect 459704 3408 459710 3420
rect 460842 3408 460848 3420
rect 460900 3408 460906 3460
rect 461872 3448 461900 3488
rect 462958 3476 462964 3528
rect 463016 3516 463022 3528
rect 464430 3516 464436 3528
rect 463016 3488 464436 3516
rect 463016 3476 463022 3488
rect 464430 3476 464436 3488
rect 464488 3476 464494 3528
rect 466362 3476 466368 3528
rect 466420 3516 466426 3528
rect 466420 3488 511212 3516
rect 466420 3476 466426 3488
rect 463234 3448 463240 3460
rect 461872 3420 463240 3448
rect 463234 3408 463240 3420
rect 463292 3408 463298 3460
rect 464338 3408 464344 3460
rect 464396 3448 464402 3460
rect 467926 3448 467932 3460
rect 464396 3420 467932 3448
rect 464396 3408 464402 3420
rect 467926 3408 467932 3420
rect 467984 3408 467990 3460
rect 468478 3408 468484 3460
rect 468536 3448 468542 3460
rect 469217 3451 469275 3457
rect 469217 3448 469229 3451
rect 468536 3420 469229 3448
rect 468536 3408 468542 3420
rect 469217 3417 469229 3420
rect 469263 3417 469275 3451
rect 469217 3411 469275 3417
rect 470502 3408 470508 3460
rect 470560 3448 470566 3460
rect 511077 3451 511135 3457
rect 511077 3448 511089 3451
rect 470560 3420 511089 3448
rect 470560 3408 470566 3420
rect 511077 3417 511089 3420
rect 511123 3417 511135 3451
rect 511184 3448 511212 3488
rect 512638 3476 512644 3528
rect 512696 3516 512702 3528
rect 514386 3516 514392 3528
rect 512696 3488 514392 3516
rect 512696 3476 512702 3488
rect 514386 3476 514392 3488
rect 514444 3476 514450 3528
rect 517422 3476 517428 3528
rect 517480 3516 517486 3528
rect 575014 3516 575020 3528
rect 517480 3488 575020 3516
rect 517480 3476 517486 3488
rect 575014 3476 575020 3488
rect 575072 3476 575078 3528
rect 513190 3448 513196 3460
rect 511184 3420 513196 3448
rect 511077 3411 511135 3417
rect 513190 3408 513196 3420
rect 513248 3408 513254 3460
rect 522942 3408 522948 3460
rect 523000 3448 523006 3460
rect 580994 3448 581000 3460
rect 523000 3420 581000 3448
rect 523000 3408 523006 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 111886 3380 111892 3392
rect 104176 3352 111892 3380
rect 111886 3340 111892 3352
rect 111944 3340 111950 3392
rect 120626 3340 120632 3392
rect 120684 3380 120690 3392
rect 121362 3380 121368 3392
rect 120684 3352 121368 3380
rect 120684 3340 120690 3352
rect 121362 3340 121368 3352
rect 121420 3340 121426 3392
rect 260742 3340 260748 3392
rect 260800 3380 260806 3392
rect 263410 3380 263416 3392
rect 260800 3352 263416 3380
rect 260800 3340 260806 3352
rect 263410 3340 263416 3352
rect 263468 3340 263474 3392
rect 281442 3340 281448 3392
rect 281500 3380 281506 3392
rect 288342 3380 288348 3392
rect 281500 3352 288348 3380
rect 281500 3340 281506 3352
rect 288342 3340 288348 3352
rect 288400 3340 288406 3392
rect 296530 3340 296536 3392
rect 296588 3380 296594 3392
rect 306190 3380 306196 3392
rect 296588 3352 306196 3380
rect 296588 3340 296594 3352
rect 306190 3340 306196 3352
rect 306248 3340 306254 3392
rect 306282 3340 306288 3392
rect 306340 3380 306346 3392
rect 318058 3380 318064 3392
rect 306340 3352 318064 3380
rect 306340 3340 306346 3352
rect 318058 3340 318064 3352
rect 318116 3340 318122 3392
rect 329742 3340 329748 3392
rect 329800 3380 329806 3392
rect 346670 3380 346676 3392
rect 329800 3352 346676 3380
rect 329800 3340 329806 3352
rect 346670 3340 346676 3352
rect 346728 3340 346734 3392
rect 347682 3340 347688 3392
rect 347740 3380 347746 3392
rect 368014 3380 368020 3392
rect 347740 3352 368020 3380
rect 347740 3340 347746 3352
rect 368014 3340 368020 3352
rect 368072 3340 368078 3392
rect 369762 3340 369768 3392
rect 369820 3380 369826 3392
rect 395430 3380 395436 3392
rect 369820 3352 395436 3380
rect 369820 3340 369826 3352
rect 395430 3340 395436 3352
rect 395488 3340 395494 3392
rect 395893 3383 395951 3389
rect 395893 3349 395905 3383
rect 395939 3380 395951 3383
rect 400214 3380 400220 3392
rect 395939 3352 400220 3380
rect 395939 3349 395951 3352
rect 395893 3343 395951 3349
rect 400214 3340 400220 3352
rect 400272 3340 400278 3392
rect 401413 3383 401471 3389
rect 401413 3349 401425 3383
rect 401459 3380 401471 3383
rect 427538 3380 427544 3392
rect 401459 3352 427544 3380
rect 401459 3349 401471 3352
rect 401413 3343 401471 3349
rect 427538 3340 427544 3352
rect 427596 3340 427602 3392
rect 431221 3383 431279 3389
rect 431221 3349 431233 3383
rect 431267 3380 431279 3383
rect 434622 3380 434628 3392
rect 431267 3352 434628 3380
rect 431267 3349 431279 3352
rect 431221 3343 431279 3349
rect 434622 3340 434628 3352
rect 434680 3340 434686 3392
rect 434717 3383 434775 3389
rect 434717 3349 434729 3383
rect 434763 3380 434775 3383
rect 471514 3380 471520 3392
rect 434763 3352 471520 3380
rect 434763 3349 434775 3352
rect 434717 3343 434775 3349
rect 471514 3340 471520 3352
rect 471572 3340 471578 3392
rect 486418 3340 486424 3392
rect 486476 3380 486482 3392
rect 489362 3380 489368 3392
rect 486476 3352 489368 3380
rect 486476 3340 486482 3352
rect 489362 3340 489368 3352
rect 489420 3340 489426 3392
rect 489822 3340 489828 3392
rect 489880 3380 489886 3392
rect 539505 3383 539563 3389
rect 539505 3380 539517 3383
rect 489880 3352 539517 3380
rect 489880 3340 489886 3352
rect 539505 3349 539517 3352
rect 539551 3349 539563 3383
rect 539505 3343 539563 3349
rect 540238 3340 540244 3392
rect 540296 3380 540302 3392
rect 542906 3380 542912 3392
rect 540296 3352 542912 3380
rect 540296 3340 540302 3352
rect 542906 3340 542912 3352
rect 542964 3340 542970 3392
rect 544378 3340 544384 3392
rect 544436 3380 544442 3392
rect 564342 3380 564348 3392
rect 544436 3352 564348 3380
rect 544436 3340 544442 3352
rect 564342 3340 564348 3352
rect 564400 3340 564406 3392
rect 83884 3284 94360 3312
rect 83884 3272 83890 3284
rect 157518 3272 157524 3324
rect 157576 3312 157582 3324
rect 158622 3312 158628 3324
rect 157576 3284 158628 3312
rect 157576 3272 157582 3284
rect 158622 3272 158628 3284
rect 158680 3272 158686 3324
rect 175366 3272 175372 3324
rect 175424 3312 175430 3324
rect 176470 3312 176476 3324
rect 175424 3284 176476 3312
rect 175424 3272 175430 3284
rect 176470 3272 176476 3284
rect 176528 3272 176534 3324
rect 226518 3272 226524 3324
rect 226576 3312 226582 3324
rect 227622 3312 227628 3324
rect 226576 3284 227628 3312
rect 226576 3272 226582 3284
rect 227622 3272 227628 3284
rect 227680 3272 227686 3324
rect 256602 3272 256608 3324
rect 256660 3312 256666 3324
rect 258626 3312 258632 3324
rect 256660 3284 258632 3312
rect 256660 3272 256666 3284
rect 258626 3272 258632 3284
rect 258684 3272 258690 3324
rect 272518 3272 272524 3324
rect 272576 3312 272582 3324
rect 276474 3312 276480 3324
rect 272576 3284 276480 3312
rect 272576 3272 272582 3284
rect 276474 3272 276480 3284
rect 276532 3272 276538 3324
rect 278682 3272 278688 3324
rect 278740 3312 278746 3324
rect 284754 3312 284760 3324
rect 278740 3284 284760 3312
rect 278740 3272 278746 3284
rect 284754 3272 284760 3284
rect 284812 3272 284818 3324
rect 304902 3272 304908 3324
rect 304960 3312 304966 3324
rect 316954 3312 316960 3324
rect 304960 3284 316960 3312
rect 304960 3272 304966 3284
rect 316954 3272 316960 3284
rect 317012 3272 317018 3324
rect 317322 3272 317328 3324
rect 317380 3312 317386 3324
rect 332410 3312 332416 3324
rect 317380 3284 332416 3312
rect 317380 3272 317386 3284
rect 332410 3272 332416 3284
rect 332468 3272 332474 3324
rect 333790 3272 333796 3324
rect 333848 3312 333854 3324
rect 351362 3312 351368 3324
rect 333848 3284 351368 3312
rect 333848 3272 333854 3284
rect 351362 3272 351368 3284
rect 351420 3272 351426 3324
rect 351822 3272 351828 3324
rect 351880 3312 351886 3324
rect 373994 3312 374000 3324
rect 351880 3284 374000 3312
rect 351880 3272 351886 3284
rect 373994 3272 374000 3284
rect 374052 3272 374058 3324
rect 375282 3272 375288 3324
rect 375340 3312 375346 3324
rect 402514 3312 402520 3324
rect 375340 3284 402520 3312
rect 375340 3272 375346 3284
rect 402514 3272 402520 3284
rect 402572 3272 402578 3324
rect 402790 3272 402796 3324
rect 402848 3312 402854 3324
rect 432322 3312 432328 3324
rect 402848 3284 432328 3312
rect 402848 3272 402854 3284
rect 432322 3272 432328 3284
rect 432380 3272 432386 3324
rect 432417 3315 432475 3321
rect 432417 3281 432429 3315
rect 432463 3312 432475 3315
rect 434809 3315 434867 3321
rect 434809 3312 434821 3315
rect 432463 3284 434821 3312
rect 432463 3281 432475 3284
rect 432417 3275 432475 3281
rect 434809 3281 434821 3284
rect 434855 3281 434867 3315
rect 434809 3275 434867 3281
rect 438762 3272 438768 3324
rect 438820 3312 438826 3324
rect 442169 3315 442227 3321
rect 442169 3312 442181 3315
rect 438820 3284 442181 3312
rect 438820 3272 438826 3284
rect 442169 3281 442181 3284
rect 442215 3281 442227 3315
rect 442169 3275 442227 3281
rect 442258 3272 442264 3324
rect 442316 3312 442322 3324
rect 473906 3312 473912 3324
rect 442316 3284 473912 3312
rect 442316 3272 442322 3284
rect 473906 3272 473912 3284
rect 473964 3272 473970 3324
rect 476022 3272 476028 3324
rect 476080 3312 476086 3324
rect 523862 3312 523868 3324
rect 476080 3284 523868 3312
rect 476080 3272 476086 3284
rect 523862 3272 523868 3284
rect 523920 3272 523926 3324
rect 530578 3272 530584 3324
rect 530636 3312 530642 3324
rect 534534 3312 534540 3324
rect 530636 3284 534540 3312
rect 530636 3272 530642 3284
rect 534534 3272 534540 3284
rect 534592 3272 534598 3324
rect 534629 3315 534687 3321
rect 534629 3281 534641 3315
rect 534675 3312 534687 3315
rect 579798 3312 579804 3324
rect 534675 3284 579804 3312
rect 534675 3281 534687 3284
rect 534629 3275 534687 3281
rect 579798 3272 579804 3284
rect 579856 3272 579862 3324
rect 44266 3244 44272 3256
rect 35912 3216 44272 3244
rect 44266 3204 44272 3216
rect 44324 3204 44330 3256
rect 70670 3204 70676 3256
rect 70728 3244 70734 3256
rect 71682 3244 71688 3256
rect 70728 3216 71688 3244
rect 70728 3204 70734 3216
rect 71682 3204 71688 3216
rect 71740 3204 71746 3256
rect 95694 3204 95700 3256
rect 95752 3244 95758 3256
rect 96522 3244 96528 3256
rect 95752 3216 96528 3244
rect 95752 3204 95758 3216
rect 96522 3204 96528 3216
rect 96580 3204 96586 3256
rect 324222 3204 324228 3256
rect 324280 3244 324286 3256
rect 339494 3244 339500 3256
rect 324280 3216 339500 3244
rect 324280 3204 324286 3216
rect 339494 3204 339500 3216
rect 339552 3204 339558 3256
rect 342162 3204 342168 3256
rect 342220 3244 342226 3256
rect 362126 3244 362132 3256
rect 342220 3216 362132 3244
rect 342220 3204 342226 3216
rect 362126 3204 362132 3216
rect 362184 3204 362190 3256
rect 376662 3204 376668 3256
rect 376720 3244 376726 3256
rect 403710 3244 403716 3256
rect 376720 3216 403716 3244
rect 376720 3204 376726 3216
rect 403710 3204 403716 3216
rect 403768 3204 403774 3256
rect 405642 3204 405648 3256
rect 405700 3244 405706 3256
rect 438210 3244 438216 3256
rect 405700 3216 438216 3244
rect 405700 3204 405706 3216
rect 438210 3204 438216 3216
rect 438268 3204 438274 3256
rect 438581 3247 438639 3253
rect 438581 3213 438593 3247
rect 438627 3244 438639 3247
rect 442445 3247 442503 3253
rect 438627 3216 442396 3244
rect 438627 3213 438639 3216
rect 438581 3207 438639 3213
rect 77846 3136 77852 3188
rect 77904 3176 77910 3188
rect 78582 3176 78588 3188
rect 77904 3148 78588 3176
rect 77904 3136 77910 3148
rect 78582 3136 78588 3148
rect 78640 3136 78646 3188
rect 88518 3136 88524 3188
rect 88576 3176 88582 3188
rect 89622 3176 89628 3188
rect 88576 3148 89628 3176
rect 88576 3136 88582 3148
rect 89622 3136 89628 3148
rect 89680 3136 89686 3188
rect 103974 3136 103980 3188
rect 104032 3176 104038 3188
rect 104802 3176 104808 3188
rect 104032 3148 104808 3176
rect 104032 3136 104038 3148
rect 104802 3136 104808 3148
rect 104860 3136 104866 3188
rect 124214 3136 124220 3188
rect 124272 3176 124278 3188
rect 125410 3176 125416 3188
rect 124272 3148 125416 3176
rect 124272 3136 124278 3148
rect 125410 3136 125416 3148
rect 125468 3136 125474 3188
rect 269022 3136 269028 3188
rect 269080 3176 269086 3188
rect 272886 3176 272892 3188
rect 269080 3148 272892 3176
rect 269080 3136 269086 3148
rect 272886 3136 272892 3148
rect 272944 3136 272950 3188
rect 318702 3136 318708 3188
rect 318760 3176 318766 3188
rect 333606 3176 333612 3188
rect 318760 3148 333612 3176
rect 318760 3136 318766 3148
rect 333606 3136 333612 3148
rect 333664 3136 333670 3188
rect 338022 3136 338028 3188
rect 338080 3176 338086 3188
rect 356146 3176 356152 3188
rect 338080 3148 356152 3176
rect 338080 3136 338086 3148
rect 356146 3136 356152 3148
rect 356204 3136 356210 3188
rect 367002 3136 367008 3188
rect 367060 3176 367066 3188
rect 391842 3176 391848 3188
rect 367060 3148 391848 3176
rect 367060 3136 367066 3148
rect 391842 3136 391848 3148
rect 391900 3136 391906 3188
rect 421558 3176 421564 3188
rect 391952 3148 421564 3176
rect 64782 3068 64788 3120
rect 64840 3108 64846 3120
rect 66898 3108 66904 3120
rect 64840 3080 66904 3108
rect 64840 3068 64846 3080
rect 66898 3068 66904 3080
rect 66956 3068 66962 3120
rect 167086 3068 167092 3120
rect 167144 3108 167150 3120
rect 168282 3108 168288 3120
rect 167144 3080 168288 3108
rect 167144 3068 167150 3080
rect 168282 3068 168288 3080
rect 168340 3068 168346 3120
rect 181346 3068 181352 3120
rect 181404 3108 181410 3120
rect 182082 3108 182088 3120
rect 181404 3080 182088 3108
rect 181404 3068 181410 3080
rect 182082 3068 182088 3080
rect 182140 3068 182146 3120
rect 262122 3068 262128 3120
rect 262180 3108 262186 3120
rect 264606 3108 264612 3120
rect 262180 3080 264612 3108
rect 262180 3068 262186 3080
rect 264606 3068 264612 3080
rect 264664 3068 264670 3120
rect 273070 3068 273076 3120
rect 273128 3108 273134 3120
rect 277670 3108 277676 3120
rect 273128 3080 277676 3108
rect 273128 3068 273134 3080
rect 277670 3068 277676 3080
rect 277728 3068 277734 3120
rect 320082 3068 320088 3120
rect 320140 3108 320146 3120
rect 334710 3108 334716 3120
rect 320140 3080 334716 3108
rect 320140 3068 320146 3080
rect 334710 3068 334716 3080
rect 334768 3068 334774 3120
rect 340506 3068 340512 3120
rect 340564 3108 340570 3120
rect 359734 3108 359740 3120
rect 340564 3080 359740 3108
rect 340564 3068 340570 3080
rect 359734 3068 359740 3080
rect 359792 3068 359798 3120
rect 361482 3068 361488 3120
rect 361540 3108 361546 3120
rect 384666 3108 384672 3120
rect 361540 3080 384672 3108
rect 361540 3068 361546 3080
rect 384666 3068 384672 3080
rect 384724 3068 384730 3120
rect 391750 3068 391756 3120
rect 391808 3108 391814 3120
rect 391952 3108 391980 3148
rect 421558 3136 421564 3148
rect 421616 3136 421622 3188
rect 422849 3179 422907 3185
rect 422849 3145 422861 3179
rect 422895 3176 422907 3179
rect 432601 3179 432659 3185
rect 432601 3176 432613 3179
rect 422895 3148 432613 3176
rect 422895 3145 422907 3148
rect 422849 3139 422907 3145
rect 432601 3145 432613 3148
rect 432647 3145 432659 3179
rect 432601 3139 432659 3145
rect 432693 3179 432751 3185
rect 432693 3145 432705 3179
rect 432739 3176 432751 3179
rect 434441 3179 434499 3185
rect 434441 3176 434453 3179
rect 432739 3148 434453 3176
rect 432739 3145 432751 3148
rect 432693 3139 432751 3145
rect 434441 3145 434453 3148
rect 434487 3145 434499 3179
rect 434441 3139 434499 3145
rect 434530 3136 434536 3188
rect 434588 3176 434594 3188
rect 442258 3176 442264 3188
rect 434588 3148 442264 3176
rect 434588 3136 434594 3148
rect 442258 3136 442264 3148
rect 442316 3136 442322 3188
rect 442368 3176 442396 3216
rect 442445 3213 442457 3247
rect 442491 3244 442503 3247
rect 478690 3244 478696 3256
rect 442491 3216 478696 3244
rect 442491 3213 442503 3216
rect 442445 3207 442503 3213
rect 478690 3204 478696 3216
rect 478748 3204 478754 3256
rect 483750 3204 483756 3256
rect 483808 3244 483814 3256
rect 488166 3244 488172 3256
rect 483808 3216 488172 3244
rect 483808 3204 483814 3216
rect 488166 3204 488172 3216
rect 488224 3204 488230 3256
rect 488442 3204 488448 3256
rect 488500 3244 488506 3256
rect 539318 3244 539324 3256
rect 488500 3216 539324 3244
rect 488500 3204 488506 3216
rect 539318 3204 539324 3216
rect 539376 3204 539382 3256
rect 539505 3247 539563 3253
rect 539505 3213 539517 3247
rect 539551 3244 539563 3247
rect 541710 3244 541716 3256
rect 539551 3216 541716 3244
rect 539551 3213 539563 3216
rect 539505 3207 539563 3213
rect 541710 3204 541716 3216
rect 541768 3204 541774 3256
rect 577406 3244 577412 3256
rect 541820 3216 577412 3244
rect 472710 3176 472716 3188
rect 442368 3148 472716 3176
rect 472710 3136 472716 3148
rect 472768 3136 472774 3188
rect 482922 3136 482928 3188
rect 482980 3176 482986 3188
rect 532234 3176 532240 3188
rect 482980 3148 532240 3176
rect 482980 3136 482986 3148
rect 532234 3136 532240 3148
rect 532292 3136 532298 3188
rect 391808 3080 391980 3108
rect 391808 3068 391814 3080
rect 399570 3068 399576 3120
rect 399628 3108 399634 3120
rect 428734 3108 428740 3120
rect 399628 3080 428740 3108
rect 399628 3068 399634 3080
rect 428734 3068 428740 3080
rect 428792 3068 428798 3120
rect 431770 3068 431776 3120
rect 431828 3108 431834 3120
rect 434717 3111 434775 3117
rect 434717 3108 434729 3111
rect 431828 3080 434729 3108
rect 431828 3068 431834 3080
rect 434717 3077 434729 3080
rect 434763 3077 434775 3111
rect 434717 3071 434775 3077
rect 434809 3111 434867 3117
rect 434809 3077 434821 3111
rect 434855 3108 434867 3111
rect 466822 3108 466828 3120
rect 434855 3080 466828 3108
rect 434855 3077 434867 3080
rect 434809 3071 434867 3077
rect 466822 3068 466828 3080
rect 466880 3068 466886 3120
rect 467098 3068 467104 3120
rect 467156 3108 467162 3120
rect 475102 3108 475108 3120
rect 467156 3080 475108 3108
rect 467156 3068 467162 3080
rect 475102 3068 475108 3080
rect 475160 3068 475166 3120
rect 481542 3068 481548 3120
rect 481600 3108 481606 3120
rect 531038 3108 531044 3120
rect 481600 3080 531044 3108
rect 481600 3068 481606 3080
rect 531038 3068 531044 3080
rect 531096 3068 531102 3120
rect 537570 3068 537576 3120
rect 537628 3108 537634 3120
rect 538769 3111 538827 3117
rect 538769 3108 538781 3111
rect 537628 3080 538781 3108
rect 537628 3068 537634 3080
rect 538769 3077 538781 3080
rect 538815 3077 538827 3111
rect 538769 3071 538827 3077
rect 538858 3068 538864 3120
rect 538916 3108 538922 3120
rect 541820 3108 541848 3216
rect 577406 3204 577412 3216
rect 577464 3204 577470 3256
rect 541897 3179 541955 3185
rect 541897 3145 541909 3179
rect 541943 3176 541955 3179
rect 570230 3176 570236 3188
rect 541943 3148 570236 3176
rect 541943 3145 541955 3148
rect 541897 3139 541955 3145
rect 570230 3136 570236 3148
rect 570288 3136 570294 3188
rect 563146 3108 563152 3120
rect 538916 3080 541848 3108
rect 543016 3080 563152 3108
rect 538916 3068 538922 3080
rect 128998 3000 129004 3052
rect 129056 3040 129062 3052
rect 129642 3040 129648 3052
rect 129056 3012 129648 3040
rect 129056 3000 129062 3012
rect 129642 3000 129648 3012
rect 129700 3000 129706 3052
rect 174170 3000 174176 3052
rect 174228 3040 174234 3052
rect 174814 3040 174820 3052
rect 174228 3012 174820 3040
rect 174228 3000 174234 3012
rect 174814 3000 174820 3012
rect 174872 3000 174878 3052
rect 190822 3000 190828 3052
rect 190880 3040 190886 3052
rect 191742 3040 191748 3052
rect 190880 3012 191748 3040
rect 190880 3000 190886 3012
rect 191742 3000 191748 3012
rect 191800 3000 191806 3052
rect 206278 3000 206284 3052
rect 206336 3040 206342 3052
rect 206922 3040 206928 3052
rect 206336 3012 206928 3040
rect 206336 3000 206342 3012
rect 206922 3000 206928 3012
rect 206980 3000 206986 3052
rect 218146 3000 218152 3052
rect 218204 3040 218210 3052
rect 219342 3040 219348 3052
rect 218204 3012 219348 3040
rect 218204 3000 218210 3012
rect 219342 3000 219348 3012
rect 219400 3000 219406 3052
rect 282822 3000 282828 3052
rect 282880 3040 282886 3052
rect 289538 3040 289544 3052
rect 282880 3012 289544 3040
rect 282880 3000 282886 3012
rect 289538 3000 289544 3012
rect 289596 3000 289602 3052
rect 332502 3000 332508 3052
rect 332560 3040 332566 3052
rect 350258 3040 350264 3052
rect 332560 3012 350264 3040
rect 332560 3000 332566 3012
rect 350258 3000 350264 3012
rect 350316 3000 350322 3052
rect 353202 3000 353208 3052
rect 353260 3040 353266 3052
rect 375190 3040 375196 3052
rect 353260 3012 375196 3040
rect 353260 3000 353266 3012
rect 375190 3000 375196 3012
rect 375248 3000 375254 3052
rect 389082 3000 389088 3052
rect 389140 3040 389146 3052
rect 417970 3040 417976 3052
rect 389140 3012 417976 3040
rect 389140 3000 389146 3012
rect 417970 3000 417976 3012
rect 418028 3000 418034 3052
rect 430482 3000 430488 3052
rect 430540 3040 430546 3052
rect 441430 3040 441436 3052
rect 430540 3012 441436 3040
rect 430540 3000 430546 3012
rect 441430 3000 441436 3012
rect 441488 3000 441494 3052
rect 441525 3043 441583 3049
rect 441525 3009 441537 3043
rect 441571 3040 441583 3043
rect 470318 3040 470324 3052
rect 441571 3012 470324 3040
rect 441571 3009 441583 3012
rect 441525 3003 441583 3009
rect 470318 3000 470324 3012
rect 470376 3000 470382 3052
rect 478138 3000 478144 3052
rect 478196 3040 478202 3052
rect 516778 3040 516784 3052
rect 478196 3012 516784 3040
rect 478196 3000 478202 3012
rect 516778 3000 516784 3012
rect 516836 3000 516842 3052
rect 529198 3000 529204 3052
rect 529256 3040 529262 3052
rect 534629 3043 534687 3049
rect 534629 3040 534641 3043
rect 529256 3012 534641 3040
rect 529256 3000 529262 3012
rect 534629 3009 534641 3012
rect 534675 3009 534687 3043
rect 534629 3003 534687 3009
rect 537478 3000 537484 3052
rect 537536 3040 537542 3052
rect 543016 3040 543044 3080
rect 563146 3068 563152 3080
rect 563204 3068 563210 3120
rect 537536 3012 543044 3040
rect 543093 3043 543151 3049
rect 537536 3000 537542 3012
rect 543093 3009 543105 3043
rect 543139 3040 543151 3043
rect 555970 3040 555976 3052
rect 543139 3012 555976 3040
rect 543139 3009 543151 3012
rect 543093 3003 543151 3009
rect 555970 3000 555976 3012
rect 556028 3000 556034 3052
rect 274542 2932 274548 2984
rect 274600 2972 274606 2984
rect 280062 2972 280068 2984
rect 274600 2944 280068 2972
rect 274600 2932 274606 2944
rect 280062 2932 280068 2944
rect 280120 2932 280126 2984
rect 291102 2932 291108 2984
rect 291160 2972 291166 2984
rect 299106 2972 299112 2984
rect 291160 2944 299112 2972
rect 291160 2932 291166 2944
rect 299106 2932 299112 2944
rect 299164 2932 299170 2984
rect 331122 2932 331128 2984
rect 331180 2972 331186 2984
rect 349062 2972 349068 2984
rect 331180 2944 349068 2972
rect 331180 2932 331186 2944
rect 349062 2932 349068 2944
rect 349120 2932 349126 2984
rect 384942 2932 384948 2984
rect 385000 2972 385006 2984
rect 413278 2972 413284 2984
rect 385000 2944 413284 2972
rect 385000 2932 385006 2944
rect 413278 2932 413284 2944
rect 413336 2932 413342 2984
rect 422938 2932 422944 2984
rect 422996 2972 423002 2984
rect 431773 2975 431831 2981
rect 431773 2972 431785 2975
rect 422996 2944 431785 2972
rect 422996 2932 423002 2944
rect 431773 2941 431785 2944
rect 431819 2941 431831 2975
rect 431773 2935 431831 2941
rect 431862 2932 431868 2984
rect 431920 2972 431926 2984
rect 434441 2975 434499 2981
rect 434441 2972 434453 2975
rect 431920 2944 434453 2972
rect 431920 2932 431926 2944
rect 434441 2941 434453 2944
rect 434487 2941 434499 2975
rect 434441 2935 434499 2941
rect 434533 2975 434591 2981
rect 434533 2941 434545 2975
rect 434579 2972 434591 2975
rect 434717 2975 434775 2981
rect 434717 2972 434729 2975
rect 434579 2944 434729 2972
rect 434579 2941 434591 2944
rect 434533 2935 434591 2941
rect 434717 2941 434729 2944
rect 434763 2941 434775 2975
rect 434717 2935 434775 2941
rect 447042 2932 447048 2984
rect 447100 2972 447106 2984
rect 469122 2972 469128 2984
rect 447100 2944 469128 2972
rect 447100 2932 447106 2944
rect 469122 2932 469128 2944
rect 469180 2932 469186 2984
rect 469217 2975 469275 2981
rect 469217 2941 469229 2975
rect 469263 2972 469275 2975
rect 482278 2972 482284 2984
rect 469263 2944 482284 2972
rect 469263 2941 469275 2944
rect 469217 2935 469275 2941
rect 482278 2932 482284 2944
rect 482336 2932 482342 2984
rect 483658 2932 483664 2984
rect 483716 2972 483722 2984
rect 520274 2972 520280 2984
rect 483716 2944 520280 2972
rect 483716 2932 483722 2944
rect 520274 2932 520280 2944
rect 520332 2932 520338 2984
rect 531958 2932 531964 2984
rect 532016 2972 532022 2984
rect 538122 2972 538128 2984
rect 532016 2944 538128 2972
rect 532016 2932 532022 2944
rect 538122 2932 538128 2944
rect 538180 2932 538186 2984
rect 538769 2975 538827 2981
rect 538769 2941 538781 2975
rect 538815 2972 538827 2975
rect 541529 2975 541587 2981
rect 541529 2972 541541 2975
rect 538815 2944 541541 2972
rect 538815 2941 538827 2944
rect 538769 2935 538827 2941
rect 541529 2941 541541 2944
rect 541575 2941 541587 2975
rect 541529 2935 541587 2941
rect 541618 2932 541624 2984
rect 541676 2972 541682 2984
rect 542817 2975 542875 2981
rect 542817 2972 542829 2975
rect 541676 2944 542829 2972
rect 541676 2932 541682 2944
rect 542817 2941 542829 2944
rect 542863 2941 542875 2975
rect 548886 2972 548892 2984
rect 542817 2935 542875 2941
rect 543016 2944 548892 2972
rect 136082 2864 136088 2916
rect 136140 2904 136146 2916
rect 136542 2904 136548 2916
rect 136140 2876 136548 2904
rect 136140 2864 136146 2876
rect 136542 2864 136548 2876
rect 136600 2864 136606 2916
rect 321462 2864 321468 2916
rect 321520 2904 321526 2916
rect 335906 2904 335912 2916
rect 321520 2876 335912 2904
rect 321520 2864 321526 2876
rect 335906 2864 335912 2876
rect 335964 2864 335970 2916
rect 382182 2864 382188 2916
rect 382240 2904 382246 2916
rect 409690 2904 409696 2916
rect 382240 2876 409696 2904
rect 382240 2864 382246 2876
rect 409690 2864 409696 2876
rect 409748 2864 409754 2916
rect 440053 2907 440111 2913
rect 440053 2873 440065 2907
rect 440099 2904 440111 2907
rect 465626 2904 465632 2916
rect 440099 2876 465632 2904
rect 440099 2873 440111 2876
rect 440053 2867 440111 2873
rect 465626 2864 465632 2876
rect 465684 2864 465690 2916
rect 496078 2864 496084 2916
rect 496136 2904 496142 2916
rect 525058 2904 525064 2916
rect 496136 2876 525064 2904
rect 496136 2864 496142 2876
rect 525058 2864 525064 2876
rect 525116 2864 525122 2916
rect 534718 2864 534724 2916
rect 534776 2904 534782 2916
rect 542909 2907 542967 2913
rect 542909 2904 542921 2907
rect 534776 2876 542921 2904
rect 534776 2864 534782 2876
rect 542909 2873 542921 2876
rect 542955 2873 542967 2907
rect 542909 2867 542967 2873
rect 23106 2796 23112 2848
rect 23164 2836 23170 2848
rect 23382 2836 23388 2848
rect 23164 2808 23388 2836
rect 23164 2796 23170 2808
rect 23382 2796 23388 2808
rect 23440 2796 23446 2848
rect 57609 2839 57667 2845
rect 57609 2805 57621 2839
rect 57655 2836 57667 2839
rect 57882 2836 57888 2848
rect 57655 2808 57888 2836
rect 57655 2805 57667 2808
rect 57609 2799 57667 2805
rect 57882 2796 57888 2808
rect 57940 2796 57946 2848
rect 92106 2796 92112 2848
rect 92164 2836 92170 2848
rect 92382 2836 92388 2848
rect 92164 2808 92388 2836
rect 92164 2796 92170 2808
rect 92382 2796 92388 2808
rect 92440 2796 92446 2848
rect 109954 2796 109960 2848
rect 110012 2836 110018 2848
rect 110322 2836 110328 2848
rect 110012 2808 110328 2836
rect 110012 2796 110018 2808
rect 110322 2796 110328 2808
rect 110380 2796 110386 2848
rect 118234 2796 118240 2848
rect 118292 2836 118298 2848
rect 118602 2836 118608 2848
rect 118292 2808 118608 2836
rect 118292 2796 118298 2808
rect 118602 2796 118608 2808
rect 118660 2796 118666 2848
rect 169386 2796 169392 2848
rect 169444 2836 169450 2848
rect 169662 2836 169668 2848
rect 169444 2808 169668 2836
rect 169444 2796 169450 2808
rect 169662 2796 169668 2808
rect 169720 2796 169726 2848
rect 417418 2796 417424 2848
rect 417476 2836 417482 2848
rect 431865 2839 431923 2845
rect 431865 2836 431877 2839
rect 417476 2808 431877 2836
rect 417476 2796 417482 2808
rect 431865 2805 431877 2808
rect 431911 2805 431923 2839
rect 450170 2836 450176 2848
rect 431865 2799 431923 2805
rect 431972 2808 450176 2836
rect 431773 2703 431831 2709
rect 431773 2669 431785 2703
rect 431819 2700 431831 2703
rect 431972 2700 432000 2808
rect 450170 2796 450176 2808
rect 450228 2796 450234 2848
rect 451737 2839 451795 2845
rect 451737 2805 451749 2839
rect 451783 2836 451795 2839
rect 477494 2836 477500 2848
rect 451783 2808 477500 2836
rect 451783 2805 451795 2808
rect 451737 2799 451795 2805
rect 477494 2796 477500 2808
rect 477552 2796 477558 2848
rect 510522 2796 510528 2848
rect 510580 2836 510586 2848
rect 518161 2839 518219 2845
rect 518161 2836 518173 2839
rect 510580 2808 518173 2836
rect 510580 2796 510586 2808
rect 518161 2805 518173 2808
rect 518207 2805 518219 2839
rect 518161 2799 518219 2805
rect 533338 2796 533344 2848
rect 533396 2836 533402 2848
rect 543016 2836 543044 2944
rect 548886 2932 548892 2944
rect 548944 2932 548950 2984
rect 543182 2864 543188 2916
rect 543240 2904 543246 2916
rect 557166 2904 557172 2916
rect 543240 2876 557172 2904
rect 543240 2864 543246 2876
rect 557166 2864 557172 2876
rect 557224 2864 557230 2916
rect 550082 2836 550088 2848
rect 533396 2808 543044 2836
rect 543108 2808 550088 2836
rect 533396 2796 533402 2808
rect 434441 2771 434499 2777
rect 434441 2737 434453 2771
rect 434487 2768 434499 2771
rect 441525 2771 441583 2777
rect 441525 2768 441537 2771
rect 434487 2740 441537 2768
rect 434487 2737 434499 2740
rect 434441 2731 434499 2737
rect 441525 2737 441537 2740
rect 441571 2737 441583 2771
rect 441525 2731 441583 2737
rect 542817 2771 542875 2777
rect 542817 2737 542829 2771
rect 542863 2768 542875 2771
rect 543108 2768 543136 2808
rect 550082 2796 550088 2808
rect 550140 2796 550146 2848
rect 542863 2740 543136 2768
rect 542863 2737 542875 2740
rect 542817 2731 542875 2737
rect 431819 2672 432000 2700
rect 431819 2669 431831 2672
rect 431773 2663 431831 2669
rect 434717 2295 434775 2301
rect 434717 2261 434729 2295
rect 434763 2292 434775 2295
rect 439406 2292 439412 2304
rect 434763 2264 439412 2292
rect 434763 2261 434775 2264
rect 434717 2255 434775 2261
rect 439406 2252 439412 2264
rect 439464 2252 439470 2304
rect 404446 620 404452 672
rect 404504 660 404510 672
rect 404504 632 404952 660
rect 404504 620 404510 632
rect 404924 604 404952 632
rect 31478 592 31484 604
rect 31439 564 31484 592
rect 31478 552 31484 564
rect 31536 552 31542 604
rect 40954 552 40960 604
rect 41012 592 41018 604
rect 41322 592 41328 604
rect 41012 564 41328 592
rect 41012 552 41018 564
rect 41322 552 41328 564
rect 41380 552 41386 604
rect 56410 592 56416 604
rect 56371 564 56416 592
rect 56410 552 56416 564
rect 56468 552 56474 604
rect 57606 592 57612 604
rect 57567 564 57612 592
rect 57606 552 57612 564
rect 57664 552 57670 604
rect 74258 552 74264 604
rect 74316 592 74322 604
rect 74442 592 74448 604
rect 74316 564 74448 592
rect 74316 552 74322 564
rect 74442 552 74448 564
rect 74500 552 74506 604
rect 100478 592 100484 604
rect 100439 564 100484 592
rect 100478 552 100484 564
rect 100536 552 100542 604
rect 108758 592 108764 604
rect 108719 564 108764 592
rect 108758 552 108764 564
rect 108816 552 108822 604
rect 254026 552 254032 604
rect 254084 592 254090 604
rect 255038 592 255044 604
rect 254084 564 255044 592
rect 254084 552 254090 564
rect 255038 552 255044 564
rect 255096 552 255102 604
rect 256694 552 256700 604
rect 256752 592 256758 604
rect 257430 592 257436 604
rect 256752 564 257436 592
rect 256752 552 256758 564
rect 257430 552 257436 564
rect 257488 552 257494 604
rect 368566 552 368572 604
rect 368624 592 368630 604
rect 369210 592 369216 604
rect 368624 564 369216 592
rect 368624 552 368630 564
rect 369210 552 369216 564
rect 369268 552 369274 604
rect 375466 552 375472 604
rect 375524 592 375530 604
rect 376386 592 376392 604
rect 375524 564 376392 592
rect 375524 552 375530 564
rect 376386 552 376392 564
rect 376444 552 376450 604
rect 379514 552 379520 604
rect 379572 592 379578 604
rect 379974 592 379980 604
rect 379572 564 379980 592
rect 379572 552 379578 564
rect 379974 552 379980 564
rect 380032 552 380038 604
rect 382458 552 382464 604
rect 382516 592 382522 604
rect 383562 592 383568 604
rect 382516 564 383568 592
rect 382516 552 382522 564
rect 383562 552 383568 564
rect 383620 552 383626 604
rect 386506 552 386512 604
rect 386564 592 386570 604
rect 387058 592 387064 604
rect 386564 564 387064 592
rect 386564 552 386570 564
rect 387058 552 387064 564
rect 387116 552 387122 604
rect 393498 552 393504 604
rect 393556 592 393562 604
rect 394234 592 394240 604
rect 393556 564 394240 592
rect 393556 552 393562 564
rect 394234 552 394240 564
rect 394292 552 394298 604
rect 397638 552 397644 604
rect 397696 592 397702 604
rect 397822 592 397828 604
rect 397696 564 397828 592
rect 397696 552 397702 564
rect 397822 552 397828 564
rect 397880 552 397886 604
rect 400398 552 400404 604
rect 400456 592 400462 604
rect 401318 592 401324 604
rect 400456 564 401324 592
rect 400456 552 400462 564
rect 401318 552 401324 564
rect 401376 552 401382 604
rect 404906 552 404912 604
rect 404964 552 404970 604
rect 411438 552 411444 604
rect 411496 592 411502 604
rect 412082 592 412088 604
rect 411496 564 412088 592
rect 411496 552 411502 564
rect 412082 552 412088 564
rect 412140 552 412146 604
rect 415486 552 415492 604
rect 415544 592 415550 604
rect 415670 592 415676 604
rect 415544 564 415676 592
rect 415544 552 415550 564
rect 415670 552 415676 564
rect 415728 552 415734 604
rect 418246 552 418252 604
rect 418304 592 418310 604
rect 419166 592 419172 604
rect 418304 564 419172 592
rect 418304 552 418310 564
rect 419166 552 419172 564
rect 419224 552 419230 604
rect 425238 552 425244 604
rect 425296 592 425302 604
rect 426342 592 426348 604
rect 425296 564 426348 592
rect 425296 552 425302 564
rect 426342 552 426348 564
rect 426400 552 426406 604
rect 433518 592 433524 604
rect 433479 564 433524 592
rect 433518 552 433524 564
rect 433576 552 433582 604
rect 445754 552 445760 604
rect 445812 592 445818 604
rect 446582 592 446588 604
rect 445812 564 446588 592
rect 445812 552 445818 564
rect 446582 552 446588 564
rect 446640 552 446646 604
rect 454126 552 454132 604
rect 454184 592 454190 604
rect 454862 592 454868 604
rect 454184 564 454868 592
rect 454184 552 454190 564
rect 454862 552 454868 564
rect 454920 552 454926 604
rect 499666 552 499672 604
rect 499724 592 499730 604
rect 500126 592 500132 604
rect 499724 564 500132 592
rect 499724 552 499730 564
rect 500126 552 500132 564
rect 500184 552 500190 604
rect 506474 552 506480 604
rect 506532 592 506538 604
rect 507210 592 507216 604
rect 506532 564 507216 592
rect 506532 552 506538 564
rect 507210 552 507216 564
rect 507268 552 507274 604
<< via1 >>
rect 154120 700952 154172 701004
rect 318800 700952 318852 701004
rect 137836 700884 137888 700936
rect 314660 700884 314712 700936
rect 252468 700816 252520 700868
rect 462320 700816 462372 700868
rect 105452 700748 105504 700800
rect 322940 700748 322992 700800
rect 256608 700680 256660 700732
rect 478512 700680 478564 700732
rect 89168 700612 89220 700664
rect 331220 700612 331272 700664
rect 72976 700544 73028 700596
rect 327080 700544 327132 700596
rect 240048 700476 240100 700528
rect 527180 700476 527232 700528
rect 40500 700408 40552 700460
rect 335360 700408 335412 700460
rect 244188 700340 244240 700392
rect 543464 700340 543516 700392
rect 24308 700272 24360 700324
rect 343640 700272 343692 700324
rect 269028 700204 269080 700256
rect 413652 700204 413704 700256
rect 170312 700136 170364 700188
rect 310520 700136 310572 700188
rect 264888 700068 264940 700120
rect 397460 700068 397512 700120
rect 202788 700000 202840 700052
rect 302240 700000 302292 700052
rect 218980 699932 219032 699984
rect 306380 699932 306432 699984
rect 281448 699864 281500 699916
rect 348792 699864 348844 699916
rect 277308 699796 277360 699848
rect 332508 699796 332560 699848
rect 267648 699728 267700 699780
rect 288440 699728 288492 699780
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 283840 699660 283892 699712
rect 293960 699660 294012 699712
rect 227628 696940 227680 696992
rect 580172 696940 580224 696992
rect 299664 688576 299716 688628
rect 300124 688576 300176 688628
rect 429384 688576 429436 688628
rect 429844 688576 429896 688628
rect 559104 688576 559156 688628
rect 559656 688576 559708 688628
rect 231768 685856 231820 685908
rect 580172 685856 580224 685908
rect 299572 684428 299624 684480
rect 429292 684428 429344 684480
rect 559012 684428 559064 684480
rect 3516 681708 3568 681760
rect 347780 681708 347832 681760
rect 364340 676175 364392 676184
rect 364340 676141 364349 676175
rect 364349 676141 364383 676175
rect 364383 676141 364392 676175
rect 364340 676132 364392 676141
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 223488 673480 223540 673532
rect 580172 673480 580224 673532
rect 3424 667904 3476 667956
rect 356060 667904 356112 667956
rect 299756 666587 299808 666596
rect 299756 666553 299765 666587
rect 299765 666553 299799 666587
rect 299799 666553 299808 666587
rect 299756 666544 299808 666553
rect 364432 666544 364484 666596
rect 429476 666587 429528 666596
rect 429476 666553 429485 666587
rect 429485 666553 429519 666587
rect 429519 666553 429528 666587
rect 429476 666544 429528 666553
rect 494152 666544 494204 666596
rect 559196 666587 559248 666596
rect 559196 666553 559205 666587
rect 559205 666553 559239 666587
rect 559239 666553 559248 666587
rect 559196 666544 559248 666553
rect 299756 659719 299808 659728
rect 299756 659685 299765 659719
rect 299765 659685 299799 659719
rect 299799 659685 299808 659719
rect 299756 659676 299808 659685
rect 299664 656956 299716 657008
rect 299572 656863 299624 656872
rect 299572 656829 299581 656863
rect 299581 656829 299615 656863
rect 299615 656829 299624 656863
rect 299572 656820 299624 656829
rect 429292 656863 429344 656872
rect 429292 656829 429301 656863
rect 429301 656829 429335 656863
rect 429335 656829 429344 656863
rect 429292 656820 429344 656829
rect 559012 656863 559064 656872
rect 559012 656829 559021 656863
rect 559021 656829 559055 656863
rect 559055 656829 559064 656863
rect 559012 656820 559064 656829
rect 364340 654100 364392 654152
rect 364524 654100 364576 654152
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 351920 652740 351972 652792
rect 215208 650020 215260 650072
rect 580172 650020 580224 650072
rect 285496 648184 285548 648236
rect 235908 648116 235960 648168
rect 298100 648116 298152 648168
rect 272892 648048 272944 648100
rect 364340 648048 364392 648100
rect 260196 647980 260248 648032
rect 247592 647912 247644 647964
rect 494060 647912 494112 647964
rect 234988 647844 235040 647896
rect 180248 647164 180300 647216
rect 386604 647164 386656 647216
rect 125508 647096 125560 647148
rect 168196 647096 168248 647148
rect 191840 647096 191892 647148
rect 407580 647096 407632 647148
rect 167644 647028 167696 647080
rect 522672 647028 522724 647080
rect 3976 646960 4028 647012
rect 365536 646960 365588 647012
rect 150808 646892 150860 646944
rect 525524 646892 525576 646944
rect 5080 646824 5132 646876
rect 382372 646824 382424 646876
rect 154948 646756 155000 646808
rect 537484 646756 537536 646808
rect 104440 646688 104492 646740
rect 140044 646688 140096 646740
rect 142344 646688 142396 646740
rect 525340 646688 525392 646740
rect 138112 646620 138164 646672
rect 525432 646620 525484 646672
rect 129740 646552 129792 646604
rect 525248 646552 525300 646604
rect 3608 646484 3660 646536
rect 432880 646484 432932 646536
rect 4988 646416 5040 646468
rect 441252 646416 441304 646468
rect 6460 646348 6512 646400
rect 445484 646348 445536 646400
rect 6276 646280 6328 646332
rect 458088 646280 458140 646332
rect 4896 646212 4948 646264
rect 466552 646212 466604 646264
rect 6184 646144 6236 646196
rect 470784 646144 470836 646196
rect 10324 646076 10376 646128
rect 483388 646076 483440 646128
rect 13084 646008 13136 646060
rect 495992 646008 496044 646060
rect 4804 645940 4856 645992
rect 491760 645940 491812 645992
rect 14464 645872 14516 645924
rect 508596 645872 508648 645924
rect 25596 645668 25648 645720
rect 378140 645668 378192 645720
rect 159180 645600 159232 645652
rect 525616 645600 525668 645652
rect 40684 645532 40736 645584
rect 416044 645532 416096 645584
rect 7932 645464 7984 645516
rect 386512 645464 386564 645516
rect 386604 645464 386656 645516
rect 580816 645464 580868 645516
rect 133972 645396 134024 645448
rect 524144 645396 524196 645448
rect 7840 645328 7892 645380
rect 399208 645328 399260 645380
rect 7748 645260 7800 645312
rect 411812 645260 411864 645312
rect 168196 645192 168248 645244
rect 580724 645192 580776 645244
rect 7656 645124 7708 645176
rect 424416 645124 424468 645176
rect 108672 645056 108724 645108
rect 523960 645056 524012 645108
rect 9220 644988 9272 645040
rect 437020 644988 437072 645040
rect 83372 644920 83424 644972
rect 522580 644920 522632 644972
rect 6368 644852 6420 644904
rect 449716 644852 449768 644904
rect 70768 644784 70820 644836
rect 522488 644784 522540 644836
rect 7564 644716 7616 644768
rect 462320 644716 462372 644768
rect 9128 644648 9180 644700
rect 474924 644648 474976 644700
rect 9036 644580 9088 644632
rect 487620 644580 487672 644632
rect 25504 644512 25556 644564
rect 512828 644512 512880 644564
rect 8944 644444 8996 644496
rect 500224 644444 500276 644496
rect 209688 644376 209740 644428
rect 523408 644376 523460 644428
rect 3884 644308 3936 644360
rect 191840 644308 191892 644360
rect 197084 644308 197136 644360
rect 523500 644308 523552 644360
rect 184480 644240 184532 644292
rect 523592 644240 523644 644292
rect 192852 644172 192904 644224
rect 531964 644172 532016 644224
rect 176016 644104 176068 644156
rect 524328 644104 524380 644156
rect 8116 644036 8168 644088
rect 361304 644036 361356 644088
rect 8024 643968 8076 644020
rect 373540 643968 373592 644020
rect 140044 643900 140096 643952
rect 580540 643900 580592 643952
rect 146944 643832 146996 643884
rect 524236 643832 524288 643884
rect 9404 643764 9456 643816
rect 402980 643764 403032 643816
rect 125784 643739 125836 643748
rect 125784 643705 125793 643739
rect 125793 643705 125827 643739
rect 125827 643705 125836 643739
rect 125784 643696 125836 643705
rect 172152 643696 172204 643748
rect 567844 643696 567896 643748
rect 117228 643671 117280 643680
rect 117228 643637 117237 643671
rect 117237 643637 117271 643671
rect 117271 643637 117280 643671
rect 117228 643628 117280 643637
rect 121368 643628 121420 643680
rect 524052 643628 524104 643680
rect 3792 643560 3844 643612
rect 419908 643560 419960 643612
rect 96344 643492 96396 643544
rect 523868 643492 523920 643544
rect 92112 643424 92164 643476
rect 525064 643424 525116 643476
rect 79600 643399 79652 643408
rect 79600 643365 79609 643399
rect 79609 643365 79643 643399
rect 79643 643365 79652 643399
rect 79600 643356 79652 643365
rect 87880 643356 87932 643408
rect 523776 643356 523828 643408
rect 45836 643288 45888 643340
rect 58440 643288 58492 643340
rect 522396 643288 522448 643340
rect 580632 643220 580684 643272
rect 522304 643152 522356 643204
rect 580448 643084 580500 643136
rect 580356 641724 580408 641776
rect 571984 640228 572036 640280
rect 580172 640228 580224 640280
rect 523408 627852 523460 627904
rect 579804 627852 579856 627904
rect 3332 624860 3384 624912
rect 8116 624860 8168 624912
rect 3332 611260 3384 611312
rect 10416 611260 10468 611312
rect 544384 593308 544436 593360
rect 579988 593308 580040 593360
rect 523500 580932 523552 580984
rect 579804 580932 579856 580984
rect 3240 568080 3292 568132
rect 8024 568080 8076 568132
rect 2780 553052 2832 553104
rect 5080 553052 5132 553104
rect 531964 546388 532016 546440
rect 579988 546388 580040 546440
rect 3056 539520 3108 539572
rect 25596 539520 25648 539572
rect 523592 534012 523644 534064
rect 579804 534012 579856 534064
rect 524328 510552 524380 510604
rect 580172 510552 580224 510604
rect 3332 509940 3384 509992
rect 7932 509940 7984 509992
rect 3332 495524 3384 495576
rect 8852 495524 8904 495576
rect 567844 487092 567896 487144
rect 579620 487092 579672 487144
rect 3332 481108 3384 481160
rect 9496 481108 9548 481160
rect 553308 462476 553360 462528
rect 560208 462476 560260 462528
rect 522672 452548 522724 452600
rect 579988 452548 580040 452600
rect 3332 452480 3384 452532
rect 7840 452480 7892 452532
rect 525616 440172 525668 440224
rect 579620 440172 579672 440224
rect 3332 424056 3384 424108
rect 9404 424056 9456 424108
rect 525524 416712 525576 416764
rect 580172 416712 580224 416764
rect 537484 405628 537536 405680
rect 579988 405628 580040 405680
rect 3056 395224 3108 395276
rect 7748 395224 7800 395276
rect 524236 393252 524288 393304
rect 579620 393252 579672 393304
rect 525432 369792 525484 369844
rect 580172 369792 580224 369844
rect 3148 367004 3200 367056
rect 40684 367004 40736 367056
rect 525340 358708 525392 358760
rect 579988 358708 580040 358760
rect 524144 346332 524196 346384
rect 579620 346332 579672 346384
rect 3148 337764 3200 337816
rect 7656 337764 7708 337816
rect 525248 311788 525300 311840
rect 580172 311788 580224 311840
rect 3332 308796 3384 308848
rect 9312 308796 9364 308848
rect 524052 299412 524104 299464
rect 580172 299412 580224 299464
rect 3608 294924 3660 294976
rect 9220 294924 9272 294976
rect 3240 280100 3292 280152
rect 6460 280100 6512 280152
rect 553308 274796 553360 274848
rect 560208 274796 560260 274848
rect 2780 266160 2832 266212
rect 4988 266160 5040 266212
rect 523960 252492 524012 252544
rect 579712 252492 579764 252544
rect 3148 251268 3200 251320
rect 6368 251268 6420 251320
rect 3148 237056 3200 237108
rect 6276 237056 6328 237108
rect 525156 229032 525208 229084
rect 580172 229032 580224 229084
rect 3332 208156 3384 208208
rect 7564 208156 7616 208208
rect 523868 205572 523920 205624
rect 580172 205572 580224 205624
rect 3056 193944 3108 193996
rect 6184 193944 6236 193996
rect 523776 182112 523828 182164
rect 580172 182112 580224 182164
rect 2780 179460 2832 179512
rect 4896 179460 4948 179512
rect 525064 171028 525116 171080
rect 580172 171028 580224 171080
rect 3148 165180 3200 165232
rect 9128 165180 9180 165232
rect 522580 158652 522632 158704
rect 580172 158652 580224 158704
rect 3332 151716 3384 151768
rect 10324 151716 10376 151768
rect 523684 135192 523736 135244
rect 580172 135192 580224 135244
rect 2964 122748 3016 122800
rect 9036 122748 9088 122800
rect 522488 111732 522540 111784
rect 579620 111732 579672 111784
rect 3240 108944 3292 108996
rect 13084 108944 13136 108996
rect 2780 93236 2832 93288
rect 4804 93236 4856 93288
rect 553308 87116 553360 87168
rect 560208 87116 560260 87168
rect 3056 79840 3108 79892
rect 8944 79840 8996 79892
rect 3332 64812 3384 64864
rect 14464 64812 14516 64864
rect 522488 64812 522540 64864
rect 580172 64812 580224 64864
rect 21916 42712 21968 42764
rect 60556 42712 60608 42764
rect 67456 42712 67508 42764
rect 69020 42780 69072 42832
rect 68928 42712 68980 42764
rect 98828 42712 98880 42764
rect 107568 42712 107620 42764
rect 131212 42712 131264 42764
rect 23388 42644 23440 42696
rect 62580 42644 62632 42696
rect 64788 42644 64840 42696
rect 19248 42576 19300 42628
rect 58624 42576 58676 42628
rect 60648 42576 60700 42628
rect 20628 42508 20680 42560
rect 59636 42508 59688 42560
rect 66168 42508 66220 42560
rect 72332 42576 72384 42628
rect 95884 42644 95936 42696
rect 99288 42644 99340 42696
rect 125232 42644 125284 42696
rect 129648 42644 129700 42696
rect 133788 42712 133840 42764
rect 153660 42712 153712 42764
rect 154488 42712 154540 42764
rect 170312 42712 170364 42764
rect 173808 42712 173860 42764
rect 185952 42712 186004 42764
rect 190368 42712 190420 42764
rect 199660 42712 199712 42764
rect 237288 42712 237340 42764
rect 238852 42712 238904 42764
rect 240048 42712 240100 42764
rect 240876 42712 240928 42764
rect 251640 42712 251692 42764
rect 252468 42712 252520 42764
rect 382832 42712 382884 42764
rect 411444 42712 411496 42764
rect 414204 42712 414256 42764
rect 422944 42712 422996 42764
rect 455328 42712 455380 42764
rect 499672 42712 499724 42764
rect 502340 42712 502392 42764
rect 543004 42712 543056 42764
rect 99748 42576 99800 42628
rect 107476 42576 107528 42628
rect 131120 42576 131172 42628
rect 134064 42644 134116 42696
rect 149704 42644 149756 42696
rect 151636 42644 151688 42696
rect 167368 42644 167420 42696
rect 169668 42644 169720 42696
rect 183008 42644 183060 42696
rect 183468 42644 183520 42696
rect 193772 42644 193824 42696
rect 399484 42644 399536 42696
rect 402244 42644 402296 42696
rect 403440 42644 403492 42696
rect 404268 42644 404320 42696
rect 404452 42644 404504 42696
rect 405648 42644 405700 42696
rect 154672 42576 154724 42628
rect 155868 42576 155920 42628
rect 171324 42576 171376 42628
rect 172428 42576 172480 42628
rect 185032 42576 185084 42628
rect 186228 42576 186280 42628
rect 196716 42576 196768 42628
rect 197268 42576 197320 42628
rect 205548 42576 205600 42628
rect 365260 42576 365312 42628
rect 390652 42576 390704 42628
rect 405372 42576 405424 42628
rect 417424 42644 417476 42696
rect 461216 42644 461268 42696
rect 506480 42644 506532 42696
rect 508228 42644 508280 42696
rect 544384 42644 544436 42696
rect 92940 42508 92992 42560
rect 96528 42508 96580 42560
rect 122288 42508 122340 42560
rect 9588 42440 9640 42492
rect 50804 42440 50856 42492
rect 50988 42440 51040 42492
rect 91008 42440 91060 42492
rect 92388 42440 92440 42492
rect 119344 42440 119396 42492
rect 13636 42372 13688 42424
rect 54760 42372 54812 42424
rect 55128 42372 55180 42424
rect 88064 42372 88116 42424
rect 89628 42372 89680 42424
rect 116400 42372 116452 42424
rect 121368 42440 121420 42492
rect 142896 42508 142948 42560
rect 144644 42508 144696 42560
rect 162492 42508 162544 42560
rect 168288 42508 168340 42560
rect 181076 42508 181128 42560
rect 182180 42508 182232 42560
rect 192852 42508 192904 42560
rect 347596 42508 347648 42560
rect 368572 42508 368624 42560
rect 374092 42508 374144 42560
rect 400404 42508 400456 42560
rect 138940 42440 138992 42492
rect 139308 42440 139360 42492
rect 157616 42440 157668 42492
rect 158628 42440 158680 42492
rect 173256 42440 173308 42492
rect 175188 42440 175240 42492
rect 186964 42440 187016 42492
rect 187608 42440 187660 42492
rect 197728 42440 197780 42492
rect 198648 42440 198700 42492
rect 206560 42440 206612 42492
rect 359372 42440 359424 42492
rect 382464 42440 382516 42492
rect 402428 42440 402480 42492
rect 433984 42576 434036 42628
rect 452384 42576 452436 42628
rect 494704 42576 494756 42628
rect 496452 42576 496504 42628
rect 541624 42576 541676 42628
rect 411260 42508 411312 42560
rect 445760 42508 445812 42560
rect 471980 42508 472032 42560
rect 483664 42508 483716 42560
rect 486700 42508 486752 42560
rect 531964 42508 532016 42560
rect 417148 42440 417200 42492
rect 451924 42440 451976 42492
rect 467104 42440 467156 42492
rect 512644 42440 512696 42492
rect 514116 42440 514168 42492
rect 545764 42440 545816 42492
rect 119988 42372 120040 42424
rect 141884 42372 141936 42424
rect 141976 42372 142028 42424
rect 159548 42372 159600 42424
rect 159916 42372 159968 42424
rect 174268 42372 174320 42424
rect 176476 42372 176528 42424
rect 187976 42372 188028 42424
rect 191748 42372 191800 42424
rect 200672 42372 200724 42424
rect 219348 42372 219400 42424
rect 223212 42372 223264 42424
rect 353484 42372 353536 42424
rect 375472 42372 375524 42424
rect 379888 42372 379940 42424
rect 408592 42372 408644 42424
rect 418160 42372 418212 42424
rect 454132 42372 454184 42424
rect 483756 42372 483808 42424
rect 530584 42372 530636 42424
rect 16488 42304 16540 42356
rect 56692 42304 56744 42356
rect 57888 42304 57940 42356
rect 62028 42304 62080 42356
rect 93860 42304 93912 42356
rect 97908 42304 97960 42356
rect 123300 42304 123352 42356
rect 125416 42304 125468 42356
rect 145840 42304 145892 42356
rect 151728 42304 151780 42356
rect 168380 42304 168432 42356
rect 171048 42304 171100 42356
rect 184020 42304 184072 42356
rect 188988 42304 189040 42356
rect 198740 42304 198792 42356
rect 200028 42304 200080 42356
rect 207572 42304 207624 42356
rect 208308 42304 208360 42356
rect 214380 42304 214432 42356
rect 356428 42304 356480 42356
rect 379520 42304 379572 42356
rect 385776 42304 385828 42356
rect 415492 42304 415544 42356
rect 428924 42304 428976 42356
rect 464344 42304 464396 42356
rect 472992 42304 473044 42356
rect 520464 42304 520516 42356
rect 522948 42304 523000 42356
rect 547236 42304 547288 42356
rect 12348 42236 12400 42288
rect 52736 42236 52788 42288
rect 56508 42236 56560 42288
rect 89996 42236 90048 42288
rect 93768 42236 93820 42288
rect 120356 42236 120408 42288
rect 122748 42236 122800 42288
rect 143816 42236 143868 42288
rect 146208 42236 146260 42288
rect 163412 42236 163464 42288
rect 165528 42236 165580 42288
rect 179144 42236 179196 42288
rect 180708 42236 180760 42288
rect 191840 42236 191892 42288
rect 209688 42236 209740 42288
rect 215392 42236 215444 42288
rect 362316 42236 362368 42288
rect 386512 42236 386564 42288
rect 388720 42236 388772 42288
rect 418252 42236 418304 42288
rect 423036 42236 423088 42288
rect 459652 42236 459704 42288
rect 469036 42236 469088 42288
rect 478144 42236 478196 42288
rect 478880 42236 478932 42288
rect 528560 42236 528612 42288
rect 10968 42168 11020 42220
rect 51816 42168 51868 42220
rect 53748 42168 53800 42220
rect 87052 42168 87104 42220
rect 91008 42168 91060 42220
rect 117412 42168 117464 42220
rect 4068 42100 4120 42152
rect 46848 42100 46900 42152
rect 46940 42100 46992 42152
rect 81164 42100 81216 42152
rect 82728 42100 82780 42152
rect 110512 42100 110564 42152
rect 117136 42100 117188 42152
rect 118608 42100 118660 42152
rect 5448 42032 5500 42084
rect 47860 42032 47912 42084
rect 49608 42032 49660 42084
rect 59912 42032 59964 42084
rect 85120 42032 85172 42084
rect 85488 42032 85540 42084
rect 113456 42032 113508 42084
rect 117228 42032 117280 42084
rect 125692 42168 125744 42220
rect 146760 42168 146812 42220
rect 147588 42168 147640 42220
rect 164424 42168 164476 42220
rect 168196 42168 168248 42220
rect 182088 42168 182140 42220
rect 184756 42168 184808 42220
rect 195796 42168 195848 42220
rect 195888 42168 195940 42220
rect 204628 42168 204680 42220
rect 206928 42168 206980 42220
rect 213368 42168 213420 42220
rect 213828 42168 213880 42220
rect 219256 42168 219308 42220
rect 368204 42168 368256 42220
rect 393504 42168 393556 42220
rect 407396 42168 407448 42220
rect 408408 42168 408460 42220
rect 425980 42168 426032 42220
rect 462964 42168 463016 42220
rect 477868 42168 477920 42220
rect 527180 42168 527232 42220
rect 140964 42100 141016 42152
rect 143448 42100 143500 42152
rect 161480 42100 161532 42152
rect 164148 42100 164200 42152
rect 178132 42100 178184 42152
rect 179328 42100 179380 42152
rect 190920 42100 190972 42152
rect 193128 42100 193180 42152
rect 201684 42100 201736 42152
rect 202788 42100 202840 42152
rect 210424 42100 210476 42152
rect 217968 42100 218020 42152
rect 222200 42100 222252 42152
rect 344652 42100 344704 42152
rect 365812 42100 365864 42152
rect 371148 42100 371200 42152
rect 397644 42100 397696 42152
rect 400496 42100 400548 42152
rect 433432 42100 433484 42152
rect 443552 42100 443604 42152
rect 485780 42100 485832 42152
rect 490656 42100 490708 42152
rect 540244 42100 540296 42152
rect 139952 42032 140004 42084
rect 142068 42032 142120 42084
rect 160468 42032 160520 42084
rect 162768 42032 162820 42084
rect 177120 42032 177172 42084
rect 177948 42032 178000 42084
rect 189908 42032 189960 42084
rect 194416 42032 194468 42084
rect 203616 42032 203668 42084
rect 219256 42032 219308 42084
rect 224224 42032 224276 42084
rect 229008 42032 229060 42084
rect 232044 42032 232096 42084
rect 350540 42032 350592 42084
rect 372712 42032 372764 42084
rect 376944 42032 376996 42084
rect 404544 42032 404596 42084
rect 408316 42032 408368 42084
rect 443000 42032 443052 42084
rect 445576 42032 445628 42084
rect 483756 42032 483808 42084
rect 484768 42032 484820 42084
rect 535460 42032 535512 42084
rect 31668 41964 31720 42016
rect 75828 41964 75880 42016
rect 105636 41964 105688 42016
rect 133052 41964 133104 42016
rect 133696 41964 133748 42016
rect 152648 41964 152700 42016
rect 153108 41964 153160 42016
rect 169300 41964 169352 42016
rect 176568 41964 176620 42016
rect 188896 41964 188948 42016
rect 394608 41964 394660 42016
rect 425244 41964 425296 42016
rect 464160 41964 464212 42016
rect 508504 41964 508556 42016
rect 520004 41964 520056 42016
rect 547144 41964 547196 42016
rect 28908 41896 28960 41948
rect 59912 41896 59964 41948
rect 96804 41896 96856 41948
rect 104808 41896 104860 41948
rect 129188 41896 129240 41948
rect 131028 41896 131080 41948
rect 150716 41896 150768 41948
rect 160008 41896 160060 41948
rect 174820 41896 174872 41948
rect 184848 41896 184900 41948
rect 194784 41896 194836 41948
rect 458272 41896 458324 41948
rect 502432 41896 502484 41948
rect 507308 41896 507360 41948
rect 537484 41896 537536 41948
rect 38476 41828 38528 41880
rect 75276 41828 75328 41880
rect 77208 41828 77260 41880
rect 78588 41828 78640 41880
rect 107660 41828 107712 41880
rect 110328 41828 110380 41880
rect 127532 41828 127584 41880
rect 135076 41828 135128 41880
rect 135168 41828 135220 41880
rect 137928 41828 137980 41880
rect 156604 41828 156656 41880
rect 157248 41828 157300 41880
rect 172244 41828 172296 41880
rect 446496 41828 446548 41880
rect 486424 41828 486476 41880
rect 495532 41828 495584 41880
rect 533344 41828 533396 41880
rect 35808 41760 35860 41812
rect 66904 41760 66956 41812
rect 74448 41760 74500 41812
rect 104716 41760 104768 41812
rect 106188 41760 106240 41812
rect 124128 41760 124180 41812
rect 144828 41760 144880 41812
rect 148968 41760 149020 41812
rect 165436 41760 165488 41812
rect 166908 41760 166960 41812
rect 180064 41760 180116 41812
rect 463148 41760 463200 41812
rect 501604 41760 501656 41812
rect 513104 41760 513156 41812
rect 537576 41760 537628 41812
rect 42708 41692 42760 41744
rect 78220 41692 78272 41744
rect 79968 41692 80020 41744
rect 108580 41692 108632 41744
rect 115848 41692 115900 41744
rect 138020 41692 138072 41744
rect 140688 41692 140740 41744
rect 158536 41692 158588 41744
rect 161388 41692 161440 41744
rect 176200 41692 176252 41744
rect 211068 41692 211120 41744
rect 217324 41692 217376 41744
rect 434812 41692 434864 41744
rect 467104 41692 467156 41744
rect 475936 41692 475988 41744
rect 496084 41692 496136 41744
rect 501420 41692 501472 41744
rect 534724 41692 534776 41744
rect 45468 41624 45520 41676
rect 80152 41624 80204 41676
rect 83372 41624 83424 41676
rect 83464 41624 83516 41676
rect 111524 41624 111576 41676
rect 111708 41624 111760 41676
rect 41328 41556 41380 41608
rect 68284 41556 68336 41608
rect 73344 41556 73396 41608
rect 73804 41556 73856 41608
rect 102692 41556 102744 41608
rect 103428 41556 103480 41608
rect 130108 41624 130160 41676
rect 132408 41624 132460 41676
rect 151452 41624 151504 41676
rect 201408 41624 201460 41676
rect 208492 41624 208544 41676
rect 212540 41624 212592 41676
rect 218336 41624 218388 41676
rect 220728 41624 220780 41676
rect 225144 41624 225196 41676
rect 440700 41624 440752 41676
rect 468484 41624 468536 41676
rect 518992 41624 519044 41676
rect 538864 41624 538916 41676
rect 128268 41556 128320 41608
rect 148784 41556 148836 41608
rect 150348 41556 150400 41608
rect 166356 41556 166408 41608
rect 202696 41556 202748 41608
rect 209504 41556 209556 41608
rect 210976 41556 211028 41608
rect 216312 41556 216364 41608
rect 224868 41556 224920 41608
rect 228088 41556 228140 41608
rect 521016 41556 521068 41608
rect 529204 41556 529256 41608
rect 46204 41488 46256 41540
rect 48872 41488 48924 41540
rect 50344 41488 50396 41540
rect 55680 41488 55732 41540
rect 57244 41488 57296 41540
rect 64512 41488 64564 41540
rect 80704 41488 80756 41540
rect 82176 41488 82228 41540
rect 86868 41488 86920 41540
rect 114100 41488 114152 41540
rect 114468 41488 114520 41540
rect 137008 41488 137060 41540
rect 204168 41488 204220 41540
rect 211436 41488 211488 41540
rect 215208 41488 215260 41540
rect 220268 41488 220320 41540
rect 222108 41488 222160 41540
rect 226156 41488 226208 41540
rect 226248 41488 226300 41540
rect 229100 41488 229152 41540
rect 230388 41488 230440 41540
rect 232964 41488 233016 41540
rect 233148 41488 233200 41540
rect 234988 41488 235040 41540
rect 257528 41488 257580 41540
rect 258724 41488 258776 41540
rect 264336 41488 264388 41540
rect 267004 41488 267056 41540
rect 271236 41488 271288 41540
rect 272524 41488 272576 41540
rect 396540 41488 396592 41540
rect 39304 41420 39356 41472
rect 60004 41420 60056 41472
rect 63500 41420 63552 41472
rect 67548 41420 67600 41472
rect 71688 41420 71740 41472
rect 101772 41420 101824 41472
rect 113088 41420 113140 41472
rect 135996 41420 136048 41472
rect 136548 41420 136600 41472
rect 155592 41420 155644 41472
rect 194508 41420 194560 41472
rect 202604 41420 202656 41472
rect 205548 41420 205600 41472
rect 212448 41420 212500 41472
rect 216588 41420 216640 41472
rect 221280 41420 221332 41472
rect 223488 41420 223540 41472
rect 227076 41420 227128 41472
rect 227628 41420 227680 41472
rect 230020 41420 230072 41472
rect 231768 41420 231820 41472
rect 233976 41420 234028 41472
rect 234528 41420 234580 41472
rect 235908 41420 235960 41472
rect 255504 41420 255556 41472
rect 256700 41420 256752 41472
rect 258448 41420 258500 41472
rect 259368 41420 259420 41472
rect 259460 41420 259512 41472
rect 261484 41420 261536 41472
rect 262404 41420 262456 41472
rect 263416 41420 263468 41472
rect 265348 41420 265400 41472
rect 266176 41420 266228 41472
rect 268292 41420 268344 41472
rect 269028 41420 269080 41472
rect 269212 41420 269264 41472
rect 270408 41420 270460 41472
rect 272156 41420 272208 41472
rect 273076 41420 273128 41472
rect 275100 41420 275152 41472
rect 275928 41420 275980 41472
rect 276112 41420 276164 41472
rect 277308 41420 277360 41472
rect 279056 41420 279108 41472
rect 280068 41420 280120 41472
rect 282000 41420 282052 41472
rect 282828 41420 282880 41472
rect 282920 41420 282972 41472
rect 284116 41420 284168 41472
rect 285864 41420 285916 41472
rect 286876 41420 286928 41472
rect 288808 41420 288860 41472
rect 289728 41420 289780 41472
rect 289820 41420 289872 41472
rect 291108 41420 291160 41472
rect 292764 41420 292816 41472
rect 293776 41420 293828 41472
rect 295708 41420 295760 41472
rect 296536 41420 296588 41472
rect 298652 41420 298704 41472
rect 299388 41420 299440 41472
rect 299572 41420 299624 41472
rect 300768 41420 300820 41472
rect 302516 41420 302568 41472
rect 303528 41420 303580 41472
rect 305460 41420 305512 41472
rect 306288 41420 306340 41472
rect 306472 41420 306524 41472
rect 307576 41420 307628 41472
rect 309416 41420 309468 41472
rect 310336 41420 310388 41472
rect 312360 41420 312412 41472
rect 313188 41420 313240 41472
rect 313280 41420 313332 41472
rect 314568 41420 314620 41472
rect 316224 41420 316276 41472
rect 317236 41420 317288 41472
rect 319168 41420 319220 41472
rect 320088 41420 320140 41472
rect 320180 41420 320232 41472
rect 321468 41420 321520 41472
rect 323124 41420 323176 41472
rect 324228 41420 324280 41472
rect 326068 41420 326120 41472
rect 326896 41420 326948 41472
rect 329012 41420 329064 41472
rect 329748 41420 329800 41472
rect 329932 41420 329984 41472
rect 331036 41420 331088 41472
rect 332876 41420 332928 41472
rect 333796 41420 333848 41472
rect 335820 41420 335872 41472
rect 336648 41420 336700 41472
rect 336832 41420 336884 41472
rect 338028 41420 338080 41472
rect 339776 41420 339828 41472
rect 340788 41420 340840 41472
rect 342720 41420 342772 41472
rect 343548 41420 343600 41472
rect 343640 41420 343692 41472
rect 344928 41420 344980 41472
rect 346584 41420 346636 41472
rect 347688 41420 347740 41472
rect 349528 41420 349580 41472
rect 350448 41420 350500 41472
rect 357440 41420 357492 41472
rect 358728 41420 358780 41472
rect 360292 41420 360344 41472
rect 361488 41420 361540 41472
rect 363236 41420 363288 41472
rect 364248 41420 364300 41472
rect 366180 41420 366232 41472
rect 367008 41420 367060 41472
rect 367192 41420 367244 41472
rect 368388 41420 368440 41472
rect 370136 41420 370188 41472
rect 371148 41420 371200 41472
rect 373080 41420 373132 41472
rect 373908 41420 373960 41472
rect 380900 41420 380952 41472
rect 382188 41420 382240 41472
rect 383844 41420 383896 41472
rect 384948 41420 385000 41472
rect 386788 41420 386840 41472
rect 387708 41420 387760 41472
rect 387800 41420 387852 41472
rect 389088 41420 389140 41472
rect 389732 41420 389784 41472
rect 390468 41420 390520 41472
rect 390744 41420 390796 41472
rect 391848 41420 391900 41472
rect 393596 41420 393648 41472
rect 394608 41420 394660 41472
rect 397552 41420 397604 41472
rect 398656 41420 398708 41472
rect 436744 41488 436796 41540
rect 443644 41488 443696 41540
rect 410248 41420 410300 41472
rect 411168 41420 411220 41472
rect 420092 41420 420144 41472
rect 420828 41420 420880 41472
rect 421104 41420 421156 41472
rect 422116 41420 422168 41472
rect 424048 41420 424100 41472
rect 424876 41420 424928 41472
rect 426900 41420 426952 41472
rect 427728 41420 427780 41472
rect 427912 41420 427964 41472
rect 429108 41420 429160 41472
rect 430856 41420 430908 41472
rect 431868 41420 431920 41472
rect 433800 41420 433852 41472
rect 434628 41420 434680 41472
rect 437756 41420 437808 41472
rect 438768 41420 438820 41472
rect 441620 41420 441672 41472
rect 442816 41420 442868 41472
rect 444564 41420 444616 41472
rect 445668 41420 445720 41472
rect 447508 41420 447560 41472
rect 448428 41420 448480 41472
rect 448520 41420 448572 41472
rect 449716 41420 449768 41472
rect 450452 41420 450504 41472
rect 451188 41420 451240 41472
rect 451464 41420 451516 41472
rect 452568 41420 452620 41472
rect 454408 41420 454460 41472
rect 455328 41420 455380 41472
rect 465172 41420 465224 41472
rect 466276 41420 466328 41472
rect 468116 41420 468168 41472
rect 469128 41420 469180 41472
rect 471060 41420 471112 41472
rect 471888 41420 471940 41472
rect 474924 41420 474976 41472
rect 476028 41420 476080 41472
rect 480812 41420 480864 41472
rect 481548 41420 481600 41472
rect 481824 41420 481876 41472
rect 482928 41420 482980 41472
rect 488632 41420 488684 41472
rect 489736 41420 489788 41472
rect 491576 41420 491628 41472
rect 492496 41420 492548 41472
rect 494520 41420 494572 41472
rect 495348 41420 495400 41472
rect 498476 41420 498528 41472
rect 499488 41420 499540 41472
rect 505284 41420 505336 41472
rect 506388 41420 506440 41472
rect 509240 41420 509292 41472
rect 510436 41420 510488 41472
rect 511172 41420 511224 41472
rect 511908 41420 511960 41472
rect 512184 41420 512236 41472
rect 513288 41420 513340 41472
rect 515128 41420 515180 41472
rect 515956 41420 516008 41472
rect 521936 41420 521988 41472
rect 522948 41420 523000 41472
rect 399484 41284 399536 41336
rect 238852 39992 238904 40044
rect 239588 39992 239640 40044
rect 108948 38675 109000 38684
rect 108948 38641 108957 38675
rect 108957 38641 108991 38675
rect 108991 38641 109000 38675
rect 108948 38632 109000 38641
rect 31668 38607 31720 38616
rect 31668 38573 31677 38607
rect 31677 38573 31711 38607
rect 31711 38573 31720 38607
rect 31668 38564 31720 38573
rect 53380 38564 53432 38616
rect 73528 38607 73580 38616
rect 73528 38573 73537 38607
rect 73537 38573 73571 38607
rect 73571 38573 73580 38607
rect 73528 38564 73580 38573
rect 75736 38564 75788 38616
rect 75828 38564 75880 38616
rect 244280 38564 244332 38616
rect 244372 38564 244424 38616
rect 246028 38564 246080 38616
rect 108948 38539 109000 38548
rect 108948 38505 108957 38539
rect 108957 38505 108991 38539
rect 108991 38505 109000 38539
rect 108948 38496 109000 38505
rect 75736 37247 75788 37256
rect 75736 37213 75745 37247
rect 75745 37213 75779 37247
rect 75779 37213 75788 37247
rect 244372 37247 244424 37256
rect 75736 37204 75788 37213
rect 244372 37213 244381 37247
rect 244381 37213 244415 37247
rect 244415 37213 244424 37247
rect 244372 37204 244424 37213
rect 433432 37247 433484 37256
rect 433432 37213 433441 37247
rect 433441 37213 433475 37247
rect 433475 37213 433484 37247
rect 433432 37204 433484 37213
rect 241612 35912 241664 35964
rect 242532 35912 242584 35964
rect 3424 35844 3476 35896
rect 25504 35844 25556 35896
rect 175188 35844 175240 35896
rect 56876 31764 56928 31816
rect 57428 31764 57480 31816
rect 31668 29019 31720 29028
rect 31668 28985 31677 29019
rect 31677 28985 31711 29019
rect 31711 28985 31720 29019
rect 31668 28976 31720 28985
rect 53288 29019 53340 29028
rect 53288 28985 53297 29019
rect 53297 28985 53331 29019
rect 53331 28985 53340 29019
rect 53288 28976 53340 28985
rect 73620 28976 73672 29028
rect 96620 28976 96672 29028
rect 97540 28976 97592 29028
rect 108948 29019 109000 29028
rect 108948 28985 108957 29019
rect 108957 28985 108991 29019
rect 108991 28985 109000 29019
rect 108948 28976 109000 28985
rect 175004 29019 175056 29028
rect 175004 28985 175013 29019
rect 175013 28985 175047 29019
rect 175047 28985 175056 29019
rect 175004 28976 175056 28985
rect 245936 29019 245988 29028
rect 245936 28985 245945 29019
rect 245945 28985 245979 29019
rect 245979 28985 245988 29019
rect 245936 28976 245988 28985
rect 75828 27616 75880 27668
rect 244280 27616 244332 27668
rect 433432 27659 433484 27668
rect 433432 27625 433441 27659
rect 433441 27625 433475 27659
rect 433475 27625 433484 27659
rect 433432 27616 433484 27625
rect 117412 27548 117464 27600
rect 120172 27548 120224 27600
rect 244280 22763 244332 22772
rect 244280 22729 244289 22763
rect 244289 22729 244323 22763
rect 244323 22729 244332 22763
rect 244280 22720 244332 22729
rect 52552 22108 52604 22160
rect 53288 22108 53340 22160
rect 175004 22108 175056 22160
rect 174820 22040 174872 22092
rect 245844 22040 245896 22092
rect 246028 22040 246080 22092
rect 75828 20952 75880 21004
rect 100668 19524 100720 19576
rect 100668 19388 100720 19440
rect 96620 19320 96672 19372
rect 96712 19320 96764 19372
rect 31484 19252 31536 19304
rect 31668 19252 31720 19304
rect 108764 19252 108816 19304
rect 108948 19252 109000 19304
rect 246028 19295 246080 19304
rect 246028 19261 246037 19295
rect 246037 19261 246071 19295
rect 246071 19261 246080 19295
rect 246028 19252 246080 19261
rect 404728 19252 404780 19304
rect 433432 17935 433484 17944
rect 433432 17901 433441 17935
rect 433441 17901 433475 17935
rect 433475 17901 433484 17935
rect 433432 17892 433484 17901
rect 522304 17892 522356 17944
rect 579804 17892 579856 17944
rect 120448 12427 120500 12436
rect 120448 12393 120457 12427
rect 120457 12393 120491 12427
rect 120491 12393 120500 12427
rect 120448 12384 120500 12393
rect 125324 12384 125376 12436
rect 125508 12384 125560 12436
rect 252284 12384 252336 12436
rect 252468 12384 252520 12436
rect 75460 9707 75512 9716
rect 75460 9673 75469 9707
rect 75469 9673 75503 9707
rect 75503 9673 75512 9707
rect 75460 9664 75512 9673
rect 117688 9707 117740 9716
rect 117688 9673 117697 9707
rect 117697 9673 117731 9707
rect 117731 9673 117740 9707
rect 117688 9664 117740 9673
rect 244372 9664 244424 9716
rect 246028 9707 246080 9716
rect 246028 9673 246037 9707
rect 246037 9673 246071 9707
rect 246071 9673 246080 9707
rect 246028 9664 246080 9673
rect 404452 9707 404504 9716
rect 404452 9673 404461 9707
rect 404461 9673 404495 9707
rect 404495 9673 404504 9707
rect 404452 9664 404504 9673
rect 31668 9596 31720 9648
rect 100668 9596 100720 9648
rect 108948 9596 109000 9648
rect 433432 8415 433484 8424
rect 433432 8381 433441 8415
rect 433441 8381 433475 8415
rect 433475 8381 433484 8415
rect 433432 8372 433484 8381
rect 433432 8236 433484 8288
rect 471888 6536 471940 6588
rect 519084 6536 519136 6588
rect 474648 6468 474700 6520
rect 522672 6468 522724 6520
rect 477408 6400 477460 6452
rect 526260 6400 526312 6452
rect 513288 6332 513340 6384
rect 569040 6332 569092 6384
rect 515956 6264 516008 6316
rect 572628 6264 572680 6316
rect 506296 6196 506348 6248
rect 561956 6196 562008 6248
rect 469128 6128 469180 6180
rect 515588 6128 515640 6180
rect 518808 6128 518860 6180
rect 576216 6128 576268 6180
rect 466276 5448 466328 5500
rect 512000 5448 512052 5500
rect 340512 5312 340564 5364
rect 340788 5312 340840 5364
rect 422116 5312 422168 5364
rect 480168 5380 480220 5432
rect 529848 5380 529900 5432
rect 489736 5312 489788 5364
rect 540520 5312 540572 5364
rect 37372 5244 37424 5296
rect 73252 5244 73304 5296
rect 456708 5244 456760 5296
rect 482836 5244 482888 5296
rect 533436 5244 533488 5296
rect 33876 5176 33928 5228
rect 70492 5176 70544 5228
rect 398656 5176 398708 5228
rect 429936 5176 429988 5228
rect 445668 5176 445720 5228
rect 486976 5176 487028 5228
rect 495348 5176 495400 5228
rect 547696 5176 547748 5228
rect 30288 5108 30340 5160
rect 67640 5108 67692 5160
rect 404268 5108 404320 5160
rect 437020 5108 437072 5160
rect 442816 5108 442868 5160
rect 483480 5108 483532 5160
rect 485688 5108 485740 5160
rect 536932 5108 536984 5160
rect 26700 5040 26752 5092
rect 64880 5040 64932 5092
rect 407028 5040 407080 5092
rect 440608 5040 440660 5092
rect 448428 5040 448480 5092
rect 490564 5040 490616 5092
rect 492496 5040 492548 5092
rect 544108 5040 544160 5092
rect 22008 4972 22060 5024
rect 60740 4972 60792 5024
rect 409788 4972 409840 5024
rect 444196 4972 444248 5024
rect 453948 4972 454000 5024
rect 497740 4972 497792 5024
rect 498108 4972 498160 5024
rect 551192 4972 551244 5024
rect 17224 4904 17276 4956
rect 56692 4904 56744 4956
rect 415308 4904 415360 4956
rect 451280 4904 451332 4956
rect 458456 4904 458508 4956
rect 501236 4904 501288 4956
rect 503628 4904 503680 4956
rect 558368 4904 558420 4956
rect 12440 4836 12492 4888
rect 52644 4836 52696 4888
rect 412548 4836 412600 4888
rect 447784 4836 447836 4888
rect 451188 4836 451240 4888
rect 494152 4836 494204 4888
rect 500868 4836 500920 4888
rect 554780 4836 554832 4888
rect 7656 4768 7708 4820
rect 49792 4768 49844 4820
rect 73068 4768 73120 4820
rect 103612 4768 103664 4820
rect 391756 4768 391808 4820
rect 422760 4768 422812 4820
rect 424876 4768 424928 4820
rect 462044 4768 462096 4820
rect 462228 4768 462280 4820
rect 508412 4768 508464 4820
rect 510436 4768 510488 4820
rect 565544 4768 565596 4820
rect 459468 4700 459520 4752
rect 504824 4700 504876 4752
rect 120448 4360 120500 4412
rect 16028 4088 16080 4140
rect 16488 4088 16540 4140
rect 18328 4088 18380 4140
rect 19248 4088 19300 4140
rect 19524 4088 19576 4140
rect 20628 4088 20680 4140
rect 20720 4088 20772 4140
rect 21916 4088 21968 4140
rect 36176 4088 36228 4140
rect 29092 4020 29144 4072
rect 39304 4020 39356 4072
rect 54024 4088 54076 4140
rect 55128 4088 55180 4140
rect 60004 4088 60056 4140
rect 60648 4088 60700 4140
rect 71872 4088 71924 4140
rect 73804 4088 73856 4140
rect 80704 4088 80756 4140
rect 84936 4088 84988 4140
rect 85488 4088 85540 4140
rect 86132 4088 86184 4140
rect 86868 4088 86920 4140
rect 93308 4088 93360 4140
rect 93768 4088 93820 4140
rect 96896 4088 96948 4140
rect 97908 4088 97960 4140
rect 102784 4088 102836 4140
rect 103428 4088 103480 4140
rect 106372 4088 106424 4140
rect 107476 4088 107528 4140
rect 111156 4088 111208 4140
rect 111708 4088 111760 4140
rect 112352 4088 112404 4140
rect 113088 4088 113140 4140
rect 113548 4088 113600 4140
rect 114468 4088 114520 4140
rect 115940 4088 115992 4140
rect 117228 4088 117280 4140
rect 119436 4088 119488 4140
rect 119988 4088 120040 4140
rect 127808 4088 127860 4140
rect 128268 4088 128320 4140
rect 170588 4088 170640 4140
rect 171048 4088 171100 4140
rect 171784 4088 171836 4140
rect 172428 4088 172480 4140
rect 238392 4088 238444 4140
rect 238852 4088 238904 4140
rect 240784 4088 240836 4140
rect 241428 4088 241480 4140
rect 246028 4088 246080 4140
rect 246764 4088 246816 4140
rect 247040 4088 247092 4140
rect 247960 4088 248012 4140
rect 248512 4088 248564 4140
rect 249156 4088 249208 4140
rect 249708 4088 249760 4140
rect 250352 4088 250404 4140
rect 252560 4088 252612 4140
rect 253848 4088 253900 4140
rect 267004 4088 267056 4140
rect 268108 4088 268160 4140
rect 303528 4088 303580 4140
rect 314384 4088 314436 4140
rect 314568 4088 314620 4140
rect 327632 4088 327684 4140
rect 328368 4088 328420 4140
rect 345480 4088 345532 4140
rect 346308 4088 346360 4140
rect 366916 4088 366968 4140
rect 368388 4088 368440 4140
rect 393044 4088 393096 4140
rect 394608 4088 394660 4140
rect 425152 4088 425204 4140
rect 427728 4088 427780 4140
rect 68284 4020 68336 4072
rect 69480 4020 69532 4072
rect 100852 4020 100904 4072
rect 252284 4020 252336 4072
rect 252652 4020 252704 4072
rect 289728 4020 289780 4072
rect 297916 4020 297968 4072
rect 310336 4020 310388 4072
rect 322756 4020 322808 4072
rect 325608 4020 325660 4072
rect 341892 4020 341944 4072
rect 344928 4020 344980 4072
rect 364524 4020 364576 4072
rect 371148 4020 371200 4072
rect 396632 4020 396684 4072
rect 398748 4020 398800 4072
rect 431132 4020 431184 4072
rect 433984 4088 434036 4140
rect 435824 4088 435876 4140
rect 436008 4088 436060 4140
rect 476304 4088 476356 4140
rect 499488 4088 499540 4140
rect 552388 4088 552440 4140
rect 440148 4020 440200 4072
rect 481088 4020 481140 4072
rect 492588 4020 492640 4072
rect 545304 4020 545356 4072
rect 545764 4020 545816 4072
rect 571432 4020 571484 4072
rect 25504 3952 25556 4004
rect 57244 3952 57296 4004
rect 65984 3952 66036 4004
rect 96804 3952 96856 4004
rect 295248 3952 295300 4004
rect 305000 3952 305052 4004
rect 307576 3952 307628 4004
rect 319260 3952 319312 4004
rect 326988 3952 327040 4004
rect 344284 3952 344336 4004
rect 350448 3952 350500 4004
rect 371608 3952 371660 4004
rect 373908 3952 373960 4004
rect 395988 3952 396040 4004
rect 401508 3952 401560 4004
rect 429108 3952 429160 4004
rect 433248 3952 433300 4004
rect 438676 3952 438728 4004
rect 479892 3952 479944 4004
rect 493968 3952 494020 4004
rect 546500 3952 546552 4004
rect 547144 3952 547196 4004
rect 578608 3952 578660 4004
rect 24308 3884 24360 3936
rect 59912 3884 59964 3936
rect 62396 3884 62448 3936
rect 93952 3884 94004 3936
rect 98092 3884 98144 3936
rect 124312 3884 124364 3936
rect 293868 3884 293920 3936
rect 303804 3884 303856 3936
rect 313188 3884 313240 3936
rect 326436 3884 326488 3936
rect 331036 3884 331088 3936
rect 347872 3884 347924 3936
rect 349068 3884 349120 3936
rect 370412 3884 370464 3936
rect 372528 3884 372580 3936
rect 399024 3884 399076 3936
rect 402244 3884 402296 3936
rect 402796 3884 402848 3936
rect 14832 3816 14884 3868
rect 50344 3816 50396 3868
rect 55220 3816 55272 3868
rect 82636 3816 82688 3868
rect 83464 3816 83516 3868
rect 101588 3816 101640 3868
rect 127072 3816 127124 3868
rect 273168 3816 273220 3868
rect 278872 3816 278924 3868
rect 285588 3816 285640 3868
rect 293132 3816 293184 3868
rect 293776 3816 293828 3868
rect 302608 3816 302660 3868
rect 303436 3816 303488 3868
rect 315764 3816 315816 3868
rect 315948 3816 316000 3868
rect 330024 3816 330076 3868
rect 336648 3816 336700 3868
rect 354956 3816 355008 3868
rect 355968 3816 356020 3868
rect 378784 3816 378836 3868
rect 379428 3816 379480 3868
rect 407304 3816 407356 3868
rect 6460 3612 6512 3664
rect 2872 3544 2924 3596
rect 39764 3748 39816 3800
rect 76104 3748 76156 3800
rect 79048 3748 79100 3800
rect 79968 3748 80020 3800
rect 80244 3748 80296 3800
rect 109040 3748 109092 3800
rect 277308 3748 277360 3800
rect 282460 3748 282512 3800
rect 284208 3748 284260 3800
rect 291936 3748 291988 3800
rect 292488 3748 292540 3800
rect 301412 3748 301464 3800
rect 302148 3748 302200 3800
rect 313372 3748 313424 3800
rect 314476 3748 314528 3800
rect 328828 3748 328880 3800
rect 335268 3748 335320 3800
rect 353760 3748 353812 3800
rect 354588 3748 354640 3800
rect 377588 3748 377640 3800
rect 378048 3748 378100 3800
rect 406108 3748 406160 3800
rect 408408 3748 408460 3800
rect 441804 3884 441856 3936
rect 443644 3884 443696 3936
rect 449808 3884 449860 3936
rect 451924 3884 451976 3936
rect 453672 3884 453724 3936
rect 457260 3884 457312 3936
rect 495348 3884 495400 3936
rect 508504 3884 508556 3936
rect 510804 3884 510856 3936
rect 559564 3884 559616 3936
rect 411168 3816 411220 3868
rect 445392 3816 445444 3868
rect 452476 3816 452528 3868
rect 416688 3748 416740 3800
rect 449716 3748 449768 3800
rect 491760 3816 491812 3868
rect 501604 3816 501656 3868
rect 27896 3680 27948 3732
rect 28908 3680 28960 3732
rect 32680 3680 32732 3732
rect 70400 3680 70452 3732
rect 76656 3680 76708 3732
rect 106280 3680 106332 3732
rect 45652 3612 45704 3664
rect 56508 3612 56560 3664
rect 58808 3612 58860 3664
rect 91100 3612 91152 3664
rect 94504 3612 94556 3664
rect 121828 3680 121880 3732
rect 122748 3680 122800 3732
rect 227720 3680 227772 3732
rect 230572 3680 230624 3732
rect 267648 3680 267700 3732
rect 271696 3680 271748 3732
rect 300676 3680 300728 3732
rect 312176 3680 312228 3732
rect 317236 3680 317288 3732
rect 331220 3680 331272 3732
rect 333888 3680 333940 3732
rect 352564 3680 352616 3732
rect 358728 3680 358780 3732
rect 381176 3680 381228 3732
rect 382096 3680 382148 3732
rect 410892 3680 410944 3732
rect 413928 3680 413980 3732
rect 448980 3680 449032 3732
rect 123024 3612 123076 3664
rect 124128 3612 124180 3664
rect 275928 3612 275980 3664
rect 281264 3612 281316 3664
rect 284116 3612 284168 3664
rect 290740 3612 290792 3664
rect 291016 3612 291068 3664
rect 300308 3612 300360 3664
rect 300768 3612 300820 3664
rect 310980 3612 311032 3664
rect 311808 3612 311860 3664
rect 325240 3612 325292 3664
rect 326896 3612 326948 3664
rect 343088 3612 343140 3664
rect 343548 3612 343600 3664
rect 363328 3612 363380 3664
rect 364248 3612 364300 3664
rect 388260 3612 388312 3664
rect 390468 3612 390520 3664
rect 420368 3612 420420 3664
rect 420828 3612 420880 3664
rect 455328 3748 455380 3800
rect 498936 3748 498988 3800
rect 499396 3748 499448 3800
rect 492956 3680 493008 3732
rect 494704 3680 494756 3732
rect 496544 3680 496596 3732
rect 502432 3680 502484 3732
rect 503628 3680 503680 3732
rect 505008 3680 505060 3732
rect 506388 3816 506440 3868
rect 560760 3816 560812 3868
rect 553584 3748 553636 3800
rect 459560 3612 459612 3664
rect 572 3476 624 3528
rect 1676 3408 1728 3460
rect 46204 3544 46256 3596
rect 46940 3544 46992 3596
rect 43352 3476 43404 3528
rect 44088 3476 44140 3528
rect 44548 3476 44600 3528
rect 45468 3476 45520 3528
rect 45744 3476 45796 3528
rect 46848 3476 46900 3528
rect 50528 3476 50580 3528
rect 50988 3476 51040 3528
rect 51632 3476 51684 3528
rect 88340 3544 88392 3596
rect 89720 3544 89772 3596
rect 91008 3544 91060 3596
rect 90916 3476 90968 3528
rect 117688 3544 117740 3596
rect 150440 3544 150492 3596
rect 151636 3544 151688 3596
rect 158720 3544 158772 3596
rect 159916 3544 159968 3596
rect 183744 3544 183796 3596
rect 184848 3544 184900 3596
rect 201500 3544 201552 3596
rect 202696 3544 202748 3596
rect 236000 3544 236052 3596
rect 237380 3544 237432 3596
rect 263508 3544 263560 3596
rect 267004 3544 267056 3596
rect 270408 3544 270460 3596
rect 274088 3544 274140 3596
rect 279976 3544 280028 3596
rect 8852 3340 8904 3392
rect 9588 3340 9640 3392
rect 10048 3340 10100 3392
rect 10968 3340 11020 3392
rect 11244 3340 11296 3392
rect 12348 3340 12400 3392
rect 34980 3340 35032 3392
rect 35808 3340 35860 3392
rect 42892 3408 42944 3460
rect 52828 3408 52880 3460
rect 53748 3408 53800 3460
rect 61200 3408 61252 3460
rect 62028 3408 62080 3460
rect 63592 3408 63644 3460
rect 64788 3408 64840 3460
rect 68284 3408 68336 3460
rect 68928 3408 68980 3460
rect 81440 3408 81492 3460
rect 82728 3408 82780 3460
rect 114652 3476 114704 3528
rect 114744 3476 114796 3528
rect 115848 3476 115900 3528
rect 130200 3476 130252 3528
rect 131028 3476 131080 3528
rect 131396 3476 131448 3528
rect 132408 3476 132460 3528
rect 132592 3476 132644 3528
rect 133696 3476 133748 3528
rect 137284 3476 137336 3528
rect 137928 3476 137980 3528
rect 138480 3476 138532 3528
rect 139308 3476 139360 3528
rect 139676 3476 139728 3528
rect 140688 3476 140740 3528
rect 140872 3476 140924 3528
rect 141976 3476 142028 3528
rect 145656 3476 145708 3528
rect 146208 3476 146260 3528
rect 146852 3476 146904 3528
rect 147588 3476 147640 3528
rect 148048 3476 148100 3528
rect 148968 3476 149020 3528
rect 149244 3476 149296 3528
rect 150348 3476 150400 3528
rect 153936 3476 153988 3528
rect 154488 3476 154540 3528
rect 155132 3476 155184 3528
rect 155868 3476 155920 3528
rect 156328 3476 156380 3528
rect 157248 3476 157300 3528
rect 162308 3476 162360 3528
rect 162768 3476 162820 3528
rect 163504 3476 163556 3528
rect 164148 3476 164200 3528
rect 165896 3476 165948 3528
rect 166908 3476 166960 3528
rect 172980 3476 173032 3528
rect 173808 3476 173860 3528
rect 180156 3476 180208 3528
rect 180708 3476 180760 3528
rect 182548 3476 182600 3528
rect 183468 3476 183520 3528
rect 188436 3476 188488 3528
rect 188988 3476 189040 3528
rect 189632 3476 189684 3528
rect 190368 3476 190420 3528
rect 192024 3476 192076 3528
rect 193128 3476 193180 3528
rect 193220 3476 193272 3528
rect 194508 3476 194560 3528
rect 196808 3476 196860 3528
rect 197268 3476 197320 3528
rect 198004 3476 198056 3528
rect 198648 3476 198700 3528
rect 199200 3476 199252 3528
rect 200028 3476 200080 3528
rect 200396 3476 200448 3528
rect 201408 3476 201460 3528
rect 205088 3476 205140 3528
rect 205548 3476 205600 3528
rect 207480 3476 207532 3528
rect 208308 3476 208360 3528
rect 208676 3476 208728 3528
rect 209688 3476 209740 3528
rect 209872 3476 209924 3528
rect 210976 3476 211028 3528
rect 214656 3476 214708 3528
rect 215208 3476 215260 3528
rect 215852 3476 215904 3528
rect 216588 3476 216640 3528
rect 217048 3476 217100 3528
rect 217968 3476 218020 3528
rect 222936 3476 222988 3528
rect 223488 3476 223540 3528
rect 224132 3476 224184 3528
rect 224868 3476 224920 3528
rect 225328 3476 225380 3528
rect 226248 3476 226300 3528
rect 231308 3476 231360 3528
rect 231768 3476 231820 3528
rect 232504 3476 232556 3528
rect 233148 3476 233200 3528
rect 233700 3476 233752 3528
rect 234528 3476 234580 3528
rect 234804 3476 234856 3528
rect 236184 3476 236236 3528
rect 239588 3476 239640 3528
rect 240048 3476 240100 3528
rect 255228 3476 255280 3528
rect 256240 3476 256292 3528
rect 258724 3476 258776 3528
rect 259828 3476 259880 3528
rect 261484 3476 261536 3528
rect 262220 3476 262272 3528
rect 263416 3476 263468 3528
rect 265808 3476 265860 3528
rect 266268 3476 266320 3528
rect 270500 3476 270552 3528
rect 280068 3476 280120 3528
rect 285956 3476 286008 3528
rect 286876 3544 286928 3596
rect 294328 3544 294380 3596
rect 298008 3544 298060 3596
rect 308588 3544 308640 3596
rect 309048 3544 309100 3596
rect 321652 3544 321704 3596
rect 322848 3544 322900 3596
rect 338304 3544 338356 3596
rect 339408 3544 339460 3596
rect 358544 3544 358596 3596
rect 361396 3544 361448 3596
rect 385868 3544 385920 3596
rect 387708 3544 387760 3596
rect 416872 3544 416924 3596
rect 419448 3544 419500 3596
rect 456064 3544 456116 3596
rect 458088 3544 458140 3596
rect 502340 3612 502392 3664
rect 460848 3544 460900 3596
rect 506020 3612 506072 3664
rect 509608 3680 509660 3732
rect 511908 3680 511960 3732
rect 516048 3612 516100 3664
rect 566740 3680 566792 3732
rect 517888 3544 517940 3596
rect 567844 3612 567896 3664
rect 573824 3544 573876 3596
rect 287152 3476 287204 3528
rect 288348 3476 288400 3528
rect 296720 3476 296772 3528
rect 299388 3476 299440 3528
rect 309784 3476 309836 3528
rect 310428 3476 310480 3528
rect 324044 3476 324096 3528
rect 324136 3476 324188 3528
rect 340696 3476 340748 3528
rect 340788 3476 340840 3528
rect 360936 3476 360988 3528
rect 364156 3476 364208 3528
rect 389456 3476 389508 3528
rect 393228 3476 393280 3528
rect 423956 3476 424008 3528
rect 424968 3476 425020 3528
rect 48136 3340 48188 3392
rect 83004 3340 83056 3392
rect 42156 3272 42208 3324
rect 42708 3272 42760 3324
rect 85672 3340 85724 3392
rect 87328 3340 87380 3392
rect 83832 3272 83884 3324
rect 105176 3408 105228 3460
rect 106188 3408 106240 3460
rect 126612 3408 126664 3460
rect 147772 3408 147824 3460
rect 164700 3408 164752 3460
rect 165528 3408 165580 3460
rect 259368 3408 259420 3460
rect 261024 3408 261076 3460
rect 266176 3408 266228 3460
rect 269304 3408 269356 3460
rect 270316 3408 270368 3460
rect 275284 3408 275336 3460
rect 277216 3408 277268 3460
rect 283656 3408 283708 3460
rect 286968 3408 287020 3460
rect 295524 3408 295576 3460
rect 296628 3408 296680 3460
rect 307392 3408 307444 3460
rect 307668 3408 307720 3460
rect 320456 3408 320508 3460
rect 321376 3408 321428 3460
rect 337108 3408 337160 3460
rect 337936 3408 337988 3460
rect 357348 3408 357400 3460
rect 358636 3408 358688 3460
rect 382372 3408 382424 3460
rect 384856 3408 384908 3460
rect 414480 3408 414532 3460
rect 422208 3408 422260 3460
rect 452568 3408 452620 3460
rect 459652 3408 459704 3460
rect 460848 3408 460900 3460
rect 462964 3476 463016 3528
rect 464436 3476 464488 3528
rect 466368 3476 466420 3528
rect 463240 3408 463292 3460
rect 464344 3408 464396 3460
rect 467932 3408 467984 3460
rect 468484 3408 468536 3460
rect 470508 3408 470560 3460
rect 512644 3476 512696 3528
rect 514392 3476 514444 3528
rect 517428 3476 517480 3528
rect 575020 3476 575072 3528
rect 513196 3408 513248 3460
rect 522948 3408 523000 3460
rect 581000 3408 581052 3460
rect 111892 3340 111944 3392
rect 120632 3340 120684 3392
rect 121368 3340 121420 3392
rect 260748 3340 260800 3392
rect 263416 3340 263468 3392
rect 281448 3340 281500 3392
rect 288348 3340 288400 3392
rect 296536 3340 296588 3392
rect 306196 3340 306248 3392
rect 306288 3340 306340 3392
rect 318064 3340 318116 3392
rect 329748 3340 329800 3392
rect 346676 3340 346728 3392
rect 347688 3340 347740 3392
rect 368020 3340 368072 3392
rect 369768 3340 369820 3392
rect 395436 3340 395488 3392
rect 400220 3340 400272 3392
rect 427544 3340 427596 3392
rect 434628 3340 434680 3392
rect 471520 3340 471572 3392
rect 486424 3340 486476 3392
rect 489368 3340 489420 3392
rect 489828 3340 489880 3392
rect 540244 3340 540296 3392
rect 542912 3340 542964 3392
rect 544384 3340 544436 3392
rect 564348 3340 564400 3392
rect 157524 3272 157576 3324
rect 158628 3272 158680 3324
rect 175372 3272 175424 3324
rect 176476 3272 176528 3324
rect 226524 3272 226576 3324
rect 227628 3272 227680 3324
rect 256608 3272 256660 3324
rect 258632 3272 258684 3324
rect 272524 3272 272576 3324
rect 276480 3272 276532 3324
rect 278688 3272 278740 3324
rect 284760 3272 284812 3324
rect 304908 3272 304960 3324
rect 316960 3272 317012 3324
rect 317328 3272 317380 3324
rect 332416 3272 332468 3324
rect 333796 3272 333848 3324
rect 351368 3272 351420 3324
rect 351828 3272 351880 3324
rect 374000 3272 374052 3324
rect 375288 3272 375340 3324
rect 402520 3272 402572 3324
rect 402796 3272 402848 3324
rect 432328 3272 432380 3324
rect 438768 3272 438820 3324
rect 442264 3272 442316 3324
rect 473912 3272 473964 3324
rect 476028 3272 476080 3324
rect 523868 3272 523920 3324
rect 530584 3272 530636 3324
rect 534540 3272 534592 3324
rect 579804 3272 579856 3324
rect 44272 3204 44324 3256
rect 70676 3204 70728 3256
rect 71688 3204 71740 3256
rect 95700 3204 95752 3256
rect 96528 3204 96580 3256
rect 324228 3204 324280 3256
rect 339500 3204 339552 3256
rect 342168 3204 342220 3256
rect 362132 3204 362184 3256
rect 376668 3204 376720 3256
rect 403716 3204 403768 3256
rect 405648 3204 405700 3256
rect 438216 3204 438268 3256
rect 77852 3136 77904 3188
rect 78588 3136 78640 3188
rect 88524 3136 88576 3188
rect 89628 3136 89680 3188
rect 103980 3136 104032 3188
rect 104808 3136 104860 3188
rect 124220 3136 124272 3188
rect 125416 3136 125468 3188
rect 269028 3136 269080 3188
rect 272892 3136 272944 3188
rect 318708 3136 318760 3188
rect 333612 3136 333664 3188
rect 338028 3136 338080 3188
rect 356152 3136 356204 3188
rect 367008 3136 367060 3188
rect 391848 3136 391900 3188
rect 64788 3068 64840 3120
rect 66904 3068 66956 3120
rect 167092 3068 167144 3120
rect 168288 3068 168340 3120
rect 181352 3068 181404 3120
rect 182088 3068 182140 3120
rect 262128 3068 262180 3120
rect 264612 3068 264664 3120
rect 273076 3068 273128 3120
rect 277676 3068 277728 3120
rect 320088 3068 320140 3120
rect 334716 3068 334768 3120
rect 340512 3068 340564 3120
rect 359740 3068 359792 3120
rect 361488 3068 361540 3120
rect 384672 3068 384724 3120
rect 391756 3068 391808 3120
rect 421564 3136 421616 3188
rect 434536 3136 434588 3188
rect 442264 3136 442316 3188
rect 478696 3204 478748 3256
rect 483756 3204 483808 3256
rect 488172 3204 488224 3256
rect 488448 3204 488500 3256
rect 539324 3204 539376 3256
rect 541716 3204 541768 3256
rect 472716 3136 472768 3188
rect 482928 3136 482980 3188
rect 532240 3136 532292 3188
rect 399576 3068 399628 3120
rect 428740 3068 428792 3120
rect 431776 3068 431828 3120
rect 466828 3068 466880 3120
rect 467104 3068 467156 3120
rect 475108 3068 475160 3120
rect 481548 3068 481600 3120
rect 531044 3068 531096 3120
rect 537576 3068 537628 3120
rect 538864 3068 538916 3120
rect 577412 3204 577464 3256
rect 570236 3136 570288 3188
rect 129004 3000 129056 3052
rect 129648 3000 129700 3052
rect 174176 3000 174228 3052
rect 174820 3000 174872 3052
rect 190828 3000 190880 3052
rect 191748 3000 191800 3052
rect 206284 3000 206336 3052
rect 206928 3000 206980 3052
rect 218152 3000 218204 3052
rect 219348 3000 219400 3052
rect 282828 3000 282880 3052
rect 289544 3000 289596 3052
rect 332508 3000 332560 3052
rect 350264 3000 350316 3052
rect 353208 3000 353260 3052
rect 375196 3000 375248 3052
rect 389088 3000 389140 3052
rect 417976 3000 418028 3052
rect 430488 3000 430540 3052
rect 441436 3000 441488 3052
rect 470324 3000 470376 3052
rect 478144 3000 478196 3052
rect 516784 3000 516836 3052
rect 529204 3000 529256 3052
rect 537484 3000 537536 3052
rect 563152 3068 563204 3120
rect 555976 3000 556028 3052
rect 274548 2932 274600 2984
rect 280068 2932 280120 2984
rect 291108 2932 291160 2984
rect 299112 2932 299164 2984
rect 331128 2932 331180 2984
rect 349068 2932 349120 2984
rect 384948 2932 385000 2984
rect 413284 2932 413336 2984
rect 422944 2932 422996 2984
rect 431868 2932 431920 2984
rect 447048 2932 447100 2984
rect 469128 2932 469180 2984
rect 482284 2932 482336 2984
rect 483664 2932 483716 2984
rect 520280 2932 520332 2984
rect 531964 2932 532016 2984
rect 538128 2932 538180 2984
rect 541624 2932 541676 2984
rect 136088 2864 136140 2916
rect 136548 2864 136600 2916
rect 321468 2864 321520 2916
rect 335912 2864 335964 2916
rect 382188 2864 382240 2916
rect 409696 2864 409748 2916
rect 465632 2864 465684 2916
rect 496084 2864 496136 2916
rect 525064 2864 525116 2916
rect 534724 2864 534776 2916
rect 23112 2796 23164 2848
rect 23388 2796 23440 2848
rect 57888 2796 57940 2848
rect 92112 2796 92164 2848
rect 92388 2796 92440 2848
rect 109960 2796 110012 2848
rect 110328 2796 110380 2848
rect 118240 2796 118292 2848
rect 118608 2796 118660 2848
rect 169392 2796 169444 2848
rect 169668 2796 169720 2848
rect 417424 2796 417476 2848
rect 450176 2796 450228 2848
rect 477500 2796 477552 2848
rect 510528 2796 510580 2848
rect 533344 2796 533396 2848
rect 548892 2932 548944 2984
rect 543188 2864 543240 2916
rect 557172 2864 557224 2916
rect 550088 2796 550140 2848
rect 439412 2252 439464 2304
rect 404452 620 404504 672
rect 31484 595 31536 604
rect 31484 561 31493 595
rect 31493 561 31527 595
rect 31527 561 31536 595
rect 31484 552 31536 561
rect 40960 552 41012 604
rect 41328 552 41380 604
rect 56416 595 56468 604
rect 56416 561 56425 595
rect 56425 561 56459 595
rect 56459 561 56468 595
rect 56416 552 56468 561
rect 57612 595 57664 604
rect 57612 561 57621 595
rect 57621 561 57655 595
rect 57655 561 57664 595
rect 57612 552 57664 561
rect 74264 552 74316 604
rect 74448 552 74500 604
rect 100484 595 100536 604
rect 100484 561 100493 595
rect 100493 561 100527 595
rect 100527 561 100536 595
rect 100484 552 100536 561
rect 108764 595 108816 604
rect 108764 561 108773 595
rect 108773 561 108807 595
rect 108807 561 108816 595
rect 108764 552 108816 561
rect 254032 552 254084 604
rect 255044 552 255096 604
rect 256700 552 256752 604
rect 257436 552 257488 604
rect 368572 552 368624 604
rect 369216 552 369268 604
rect 375472 552 375524 604
rect 376392 552 376444 604
rect 379520 552 379572 604
rect 379980 552 380032 604
rect 382464 552 382516 604
rect 383568 552 383620 604
rect 386512 552 386564 604
rect 387064 552 387116 604
rect 393504 552 393556 604
rect 394240 552 394292 604
rect 397644 552 397696 604
rect 397828 552 397880 604
rect 400404 552 400456 604
rect 401324 552 401376 604
rect 404912 552 404964 604
rect 411444 552 411496 604
rect 412088 552 412140 604
rect 415492 552 415544 604
rect 415676 552 415728 604
rect 418252 552 418304 604
rect 419172 552 419224 604
rect 425244 552 425296 604
rect 426348 552 426400 604
rect 433524 595 433576 604
rect 433524 561 433533 595
rect 433533 561 433567 595
rect 433567 561 433576 595
rect 433524 552 433576 561
rect 445760 552 445812 604
rect 446588 552 446640 604
rect 454132 552 454184 604
rect 454868 552 454920 604
rect 499672 552 499724 604
rect 500132 552 500184 604
rect 506480 552 506532 604
rect 507216 552 507268 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700369 8156 703520
rect 8114 700360 8170 700369
rect 24320 700330 24348 703520
rect 40512 700466 40540 703520
rect 72988 700602 73016 703520
rect 89180 700670 89208 703520
rect 105464 700806 105492 703520
rect 137848 700942 137876 703520
rect 154132 701010 154160 703520
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 137836 700936 137888 700942
rect 137836 700878 137888 700884
rect 105452 700800 105504 700806
rect 105452 700742 105504 700748
rect 89168 700664 89220 700670
rect 89168 700606 89220 700612
rect 72976 700596 73028 700602
rect 72976 700538 73028 700544
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 8114 700295 8170 700304
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 170324 700194 170352 703520
rect 170312 700188 170364 700194
rect 170312 700130 170364 700136
rect 202800 700058 202828 703520
rect 202788 700052 202840 700058
rect 202788 699994 202840 700000
rect 218992 699990 219020 703520
rect 218980 699984 219032 699990
rect 218980 699926 219032 699932
rect 235184 699718 235212 703520
rect 252468 700868 252520 700874
rect 252468 700810 252520 700816
rect 240048 700528 240100 700534
rect 240048 700470 240100 700476
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 227628 696992 227680 696998
rect 227628 696934 227680 696940
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 223488 673532 223540 673538
rect 223488 673474 223540 673480
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 215208 650072 215260 650078
rect 215208 650014 215260 650020
rect 180248 647216 180300 647222
rect 180248 647158 180300 647164
rect 125508 647148 125560 647154
rect 125508 647090 125560 647096
rect 168196 647148 168248 647154
rect 168196 647090 168248 647096
rect 3976 647012 4028 647018
rect 3976 646954 4028 646960
rect 3608 646536 3660 646542
rect 3608 646478 3660 646484
rect 3422 646096 3478 646105
rect 3422 646031 3478 646040
rect 3332 624912 3384 624918
rect 3330 624880 3332 624889
rect 3384 624880 3386 624889
rect 3330 624815 3386 624824
rect 3332 611312 3384 611318
rect 3332 611254 3384 611260
rect 3344 610473 3372 611254
rect 3330 610464 3386 610473
rect 3330 610399 3386 610408
rect 3240 568132 3292 568138
rect 3240 568074 3292 568080
rect 3252 567361 3280 568074
rect 3238 567352 3294 567361
rect 3238 567287 3294 567296
rect 2780 553104 2832 553110
rect 2778 553072 2780 553081
rect 2832 553072 2834 553081
rect 2778 553007 2834 553016
rect 3056 539572 3108 539578
rect 3056 539514 3108 539520
rect 3068 538665 3096 539514
rect 3054 538656 3110 538665
rect 3054 538591 3110 538600
rect 3332 509992 3384 509998
rect 3330 509960 3332 509969
rect 3384 509960 3386 509969
rect 3330 509895 3386 509904
rect 3332 495576 3384 495582
rect 3330 495544 3332 495553
rect 3384 495544 3386 495553
rect 3330 495479 3386 495488
rect 3332 481160 3384 481166
rect 3330 481128 3332 481137
rect 3384 481128 3386 481137
rect 3330 481063 3386 481072
rect 3332 452532 3384 452538
rect 3332 452474 3384 452480
rect 3344 452441 3372 452474
rect 3330 452432 3386 452441
rect 3330 452367 3386 452376
rect 3332 424108 3384 424114
rect 3332 424050 3384 424056
rect 3344 423745 3372 424050
rect 3330 423736 3386 423745
rect 3330 423671 3386 423680
rect 3056 395276 3108 395282
rect 3056 395218 3108 395224
rect 3068 395049 3096 395218
rect 3054 395040 3110 395049
rect 3054 394975 3110 394984
rect 3148 367056 3200 367062
rect 3148 366998 3200 367004
rect 3160 366217 3188 366998
rect 3146 366208 3202 366217
rect 3146 366143 3202 366152
rect 3148 337816 3200 337822
rect 3148 337758 3200 337764
rect 3160 337521 3188 337758
rect 3146 337512 3202 337521
rect 3146 337447 3202 337456
rect 3332 308848 3384 308854
rect 3330 308816 3332 308825
rect 3384 308816 3386 308825
rect 3330 308751 3386 308760
rect 3240 280152 3292 280158
rect 3238 280120 3240 280129
rect 3292 280120 3294 280129
rect 3238 280055 3294 280064
rect 2780 266212 2832 266218
rect 2780 266154 2832 266160
rect 2792 265713 2820 266154
rect 2778 265704 2834 265713
rect 2778 265639 2834 265648
rect 3148 251320 3200 251326
rect 3146 251288 3148 251297
rect 3200 251288 3202 251297
rect 3146 251223 3202 251232
rect 3148 237108 3200 237114
rect 3148 237050 3200 237056
rect 3160 237017 3188 237050
rect 3146 237008 3202 237017
rect 3146 236943 3202 236952
rect 3332 208208 3384 208214
rect 3330 208176 3332 208185
rect 3384 208176 3386 208185
rect 3330 208111 3386 208120
rect 3056 193996 3108 194002
rect 3056 193938 3108 193944
rect 3068 193905 3096 193938
rect 3054 193896 3110 193905
rect 3054 193831 3110 193840
rect 2780 179512 2832 179518
rect 2778 179480 2780 179489
rect 2832 179480 2834 179489
rect 2778 179415 2834 179424
rect 3148 165232 3200 165238
rect 3148 165174 3200 165180
rect 3160 165073 3188 165174
rect 3146 165064 3202 165073
rect 3146 164999 3202 165008
rect 3332 151768 3384 151774
rect 3332 151710 3384 151716
rect 3344 150793 3372 151710
rect 3330 150784 3386 150793
rect 3330 150719 3386 150728
rect 2964 122800 3016 122806
rect 2964 122742 3016 122748
rect 2976 122097 3004 122742
rect 2962 122088 3018 122097
rect 2962 122023 3018 122032
rect 3240 108996 3292 109002
rect 3240 108938 3292 108944
rect 3252 107681 3280 108938
rect 3238 107672 3294 107681
rect 3238 107607 3294 107616
rect 2780 93288 2832 93294
rect 2778 93256 2780 93265
rect 2832 93256 2834 93265
rect 2778 93191 2834 93200
rect 3056 79892 3108 79898
rect 3056 79834 3108 79840
rect 3068 78985 3096 79834
rect 3054 78976 3110 78985
rect 3054 78911 3110 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3436 50153 3464 646031
rect 3514 642424 3570 642433
rect 3514 642359 3570 642368
rect 3528 136377 3556 642359
rect 3620 323105 3648 646478
rect 3884 644360 3936 644366
rect 3884 644302 3936 644308
rect 3792 643612 3844 643618
rect 3792 643554 3844 643560
rect 3698 642560 3754 642569
rect 3698 642495 3754 642504
rect 3606 323096 3662 323105
rect 3606 323031 3662 323040
rect 3608 294976 3660 294982
rect 3608 294918 3660 294924
rect 3620 294409 3648 294918
rect 3606 294400 3662 294409
rect 3606 294335 3662 294344
rect 3712 222601 3740 642495
rect 3804 380633 3832 643554
rect 3896 438025 3924 644302
rect 3988 596057 4016 646954
rect 53930 646912 53986 646921
rect 5080 646876 5132 646882
rect 53930 646847 53986 646856
rect 5080 646818 5132 646824
rect 4988 646468 5040 646474
rect 4988 646410 5040 646416
rect 4896 646264 4948 646270
rect 4896 646206 4948 646212
rect 4804 645992 4856 645998
rect 4804 645934 4856 645940
rect 3974 596048 4030 596057
rect 3974 595983 4030 595992
rect 3882 438016 3938 438025
rect 3882 437951 3938 437960
rect 3790 380624 3846 380633
rect 3790 380559 3846 380568
rect 3698 222592 3754 222601
rect 3698 222527 3754 222536
rect 3514 136368 3570 136377
rect 3514 136303 3570 136312
rect 4816 93294 4844 645934
rect 4908 179518 4936 646206
rect 5000 266218 5028 646410
rect 5092 553110 5120 646818
rect 6460 646400 6512 646406
rect 6460 646342 6512 646348
rect 6276 646332 6328 646338
rect 6276 646274 6328 646280
rect 6184 646196 6236 646202
rect 6184 646138 6236 646144
rect 5080 553104 5132 553110
rect 5080 553046 5132 553052
rect 4988 266212 5040 266218
rect 4988 266154 5040 266160
rect 6196 194002 6224 646138
rect 6288 237114 6316 646274
rect 6368 644904 6420 644910
rect 6368 644846 6420 644852
rect 6380 251326 6408 644846
rect 6472 280158 6500 646342
rect 10324 646128 10376 646134
rect 10324 646070 10376 646076
rect 7932 645516 7984 645522
rect 7932 645458 7984 645464
rect 7840 645380 7892 645386
rect 7840 645322 7892 645328
rect 7748 645312 7800 645318
rect 7748 645254 7800 645260
rect 7656 645176 7708 645182
rect 7656 645118 7708 645124
rect 7564 644768 7616 644774
rect 7564 644710 7616 644716
rect 6460 280152 6512 280158
rect 6460 280094 6512 280100
rect 6368 251320 6420 251326
rect 6368 251262 6420 251268
rect 6276 237108 6328 237114
rect 6276 237050 6328 237056
rect 7576 208214 7604 644710
rect 7668 337822 7696 645118
rect 7760 395282 7788 645254
rect 7852 452538 7880 645322
rect 7944 509998 7972 645458
rect 9220 645040 9272 645046
rect 9220 644982 9272 644988
rect 9128 644700 9180 644706
rect 9128 644642 9180 644648
rect 9036 644632 9088 644638
rect 9036 644574 9088 644580
rect 8944 644496 8996 644502
rect 8944 644438 8996 644444
rect 8116 644088 8168 644094
rect 8116 644030 8168 644036
rect 8024 644020 8076 644026
rect 8024 643962 8076 643968
rect 8036 568138 8064 643962
rect 8128 624918 8156 644030
rect 8850 641744 8906 641753
rect 8850 641679 8906 641688
rect 8116 624912 8168 624918
rect 8116 624854 8168 624860
rect 8024 568132 8076 568138
rect 8024 568074 8076 568080
rect 7932 509992 7984 509998
rect 7932 509934 7984 509940
rect 8864 495582 8892 641679
rect 8852 495576 8904 495582
rect 8852 495518 8904 495524
rect 7840 452532 7892 452538
rect 7840 452474 7892 452480
rect 7748 395276 7800 395282
rect 7748 395218 7800 395224
rect 7656 337816 7708 337822
rect 7656 337758 7708 337764
rect 7564 208208 7616 208214
rect 7564 208150 7616 208156
rect 6184 193996 6236 194002
rect 6184 193938 6236 193944
rect 4896 179512 4948 179518
rect 4896 179454 4948 179460
rect 4804 93288 4856 93294
rect 4804 93230 4856 93236
rect 8956 79898 8984 644438
rect 9048 122806 9076 644574
rect 9140 165238 9168 644642
rect 9232 294982 9260 644982
rect 9404 643816 9456 643822
rect 9404 643758 9456 643764
rect 9310 642968 9366 642977
rect 9310 642903 9366 642912
rect 9324 308854 9352 642903
rect 9416 424114 9444 643758
rect 9494 642288 9550 642297
rect 9494 642223 9550 642232
rect 9508 481166 9536 642223
rect 9496 481160 9548 481166
rect 9496 481102 9548 481108
rect 9404 424108 9456 424114
rect 9404 424050 9456 424056
rect 9312 308848 9364 308854
rect 9312 308790 9364 308796
rect 9220 294976 9272 294982
rect 9220 294918 9272 294924
rect 9128 165232 9180 165238
rect 9128 165174 9180 165180
rect 10336 151774 10364 646070
rect 13084 646060 13136 646066
rect 13084 646002 13136 646008
rect 10414 642152 10470 642161
rect 10414 642087 10470 642096
rect 10428 611318 10456 642087
rect 10416 611312 10468 611318
rect 10416 611254 10468 611260
rect 10324 151768 10376 151774
rect 10324 151710 10376 151716
rect 9036 122800 9088 122806
rect 9036 122742 9088 122748
rect 13096 109002 13124 646002
rect 14464 645924 14516 645930
rect 14464 645866 14516 645872
rect 13084 108996 13136 109002
rect 13084 108938 13136 108944
rect 8944 79892 8996 79898
rect 8944 79834 8996 79840
rect 14476 64870 14504 645866
rect 25596 645720 25648 645726
rect 25596 645662 25648 645668
rect 25504 644564 25556 644570
rect 25504 644506 25556 644512
rect 14464 64864 14516 64870
rect 14464 64806 14516 64812
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 21916 42764 21968 42770
rect 21916 42706 21968 42712
rect 19248 42628 19300 42634
rect 19248 42570 19300 42576
rect 9588 42492 9640 42498
rect 9588 42434 9640 42440
rect 4068 42152 4120 42158
rect 4068 42094 4120 42100
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 3476 35864 3478 35873
rect 3422 35799 3478 35808
rect 3422 8256 3478 8265
rect 3422 8191 3478 8200
rect 3436 7177 3464 8191
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 584 480 612 3470
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 480 1716 3402
rect 2884 480 2912 3538
rect 4080 480 4108 42094
rect 5448 42084 5500 42090
rect 5448 42026 5500 42032
rect 5460 4842 5488 42026
rect 5276 4814 5488 4842
rect 7656 4820 7708 4826
rect 5276 480 5304 4814
rect 7656 4762 7708 4768
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6472 480 6500 3606
rect 7668 480 7696 4762
rect 9600 3398 9628 42434
rect 13636 42424 13688 42430
rect 13636 42366 13688 42372
rect 12348 42288 12400 42294
rect 12348 42230 12400 42236
rect 10968 42220 11020 42226
rect 10968 42162 11020 42168
rect 10980 3398 11008 42162
rect 12360 3398 12388 42230
rect 12440 4888 12492 4894
rect 12440 4830 12492 4836
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 8864 480 8892 3334
rect 10060 480 10088 3334
rect 11256 480 11284 3334
rect 12452 480 12480 4830
rect 13648 480 13676 42366
rect 16488 42356 16540 42362
rect 16488 42298 16540 42304
rect 16500 4146 16528 42298
rect 17224 4956 17276 4962
rect 17224 4898 17276 4904
rect 16028 4140 16080 4146
rect 16028 4082 16080 4088
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 14832 3868 14884 3874
rect 14832 3810 14884 3816
rect 14844 480 14872 3810
rect 16040 480 16068 4082
rect 17236 480 17264 4898
rect 19260 4146 19288 42570
rect 20628 42560 20680 42566
rect 20628 42502 20680 42508
rect 20640 4146 20668 42502
rect 21928 4146 21956 42706
rect 23388 42696 23440 42702
rect 23388 42638 23440 42644
rect 22008 5024 22060 5030
rect 22008 4966 22060 4972
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 21916 4140 21968 4146
rect 21916 4082 21968 4088
rect 18340 480 18368 4082
rect 19536 480 19564 4082
rect 20732 480 20760 4082
rect 22020 2530 22048 4966
rect 23400 2854 23428 42638
rect 25516 35902 25544 644506
rect 25608 539578 25636 645662
rect 40684 645584 40736 645590
rect 40684 645526 40736 645532
rect 25596 539572 25648 539578
rect 25596 539514 25648 539520
rect 40696 367062 40724 645526
rect 53944 643892 53972 646847
rect 104440 646740 104492 646746
rect 104440 646682 104492 646688
rect 66534 646504 66590 646513
rect 66534 646439 66590 646448
rect 62394 646232 62450 646241
rect 62394 646167 62450 646176
rect 62408 643892 62436 646167
rect 66548 643892 66576 646439
rect 83372 644972 83424 644978
rect 83372 644914 83424 644920
rect 70768 644836 70820 644842
rect 70768 644778 70820 644784
rect 70780 643892 70808 644778
rect 83384 643892 83412 644914
rect 104452 643892 104480 646682
rect 112902 646368 112958 646377
rect 112902 646303 112958 646312
rect 108672 645108 108724 645114
rect 108672 645050 108724 645056
rect 108684 643892 108712 645050
rect 112916 643892 112944 646303
rect 125520 643892 125548 647090
rect 167644 647080 167696 647086
rect 167644 647022 167696 647028
rect 150808 646944 150860 646950
rect 150808 646886 150860 646892
rect 140044 646740 140096 646746
rect 140044 646682 140096 646688
rect 142344 646740 142396 646746
rect 142344 646682 142396 646688
rect 138112 646672 138164 646678
rect 138112 646614 138164 646620
rect 129740 646604 129792 646610
rect 129740 646546 129792 646552
rect 129752 643892 129780 646546
rect 133972 645448 134024 645454
rect 133972 645390 134024 645396
rect 133984 643892 134012 645390
rect 138124 643892 138152 646614
rect 140056 643958 140084 646682
rect 140044 643952 140096 643958
rect 140044 643894 140096 643900
rect 142356 643892 142384 646682
rect 146602 643890 146984 643906
rect 150820 643892 150848 646886
rect 154948 646808 155000 646814
rect 154948 646750 155000 646756
rect 154960 643892 154988 646750
rect 163410 646504 163466 646513
rect 163410 646439 163466 646448
rect 159180 645652 159232 645658
rect 159180 645594 159232 645600
rect 159192 643892 159220 645594
rect 163424 643892 163452 646439
rect 167656 643892 167684 647022
rect 168208 645250 168236 647090
rect 168196 645244 168248 645250
rect 168196 645186 168248 645192
rect 176016 644156 176068 644162
rect 176016 644098 176068 644104
rect 176028 643892 176056 644098
rect 180260 643892 180288 647158
rect 191840 647148 191892 647154
rect 191840 647090 191892 647096
rect 188618 646640 188674 646649
rect 188618 646575 188674 646584
rect 184480 644292 184532 644298
rect 184480 644234 184532 644240
rect 184492 643892 184520 644234
rect 188632 643892 188660 646575
rect 191852 644366 191880 647090
rect 201314 646776 201370 646785
rect 201314 646711 201370 646720
rect 191840 644360 191892 644366
rect 191840 644302 191892 644308
rect 197084 644360 197136 644366
rect 197084 644302 197136 644308
rect 192852 644224 192904 644230
rect 192852 644166 192904 644172
rect 192864 643892 192892 644166
rect 197096 643892 197124 644302
rect 201328 643892 201356 646711
rect 209688 644428 209740 644434
rect 209688 644370 209740 644376
rect 209700 643892 209728 644370
rect 146602 643884 146996 643890
rect 146602 643878 146944 643884
rect 146944 643826 146996 643832
rect 125782 643784 125838 643793
rect 215220 643770 215248 650014
rect 223500 643770 223528 673474
rect 227640 644042 227668 696934
rect 231768 685908 231820 685914
rect 231768 685850 231820 685856
rect 226996 644014 227668 644042
rect 226996 643770 227024 644014
rect 231780 643770 231808 685850
rect 235920 648174 235948 699654
rect 235908 648168 235960 648174
rect 235908 648110 235960 648116
rect 234988 647896 235040 647902
rect 234988 647838 235040 647844
rect 235000 643892 235028 647838
rect 240060 643770 240088 700470
rect 244188 700392 244240 700398
rect 244188 700334 244240 700340
rect 244200 643770 244228 700334
rect 247592 647964 247644 647970
rect 247592 647906 247644 647912
rect 247604 643892 247632 647906
rect 252480 643770 252508 700810
rect 256608 700732 256660 700738
rect 256608 700674 256660 700680
rect 256620 643770 256648 700674
rect 264888 700120 264940 700126
rect 264888 700062 264940 700068
rect 260196 648032 260248 648038
rect 260196 647974 260248 647980
rect 260208 643892 260236 647974
rect 264900 643770 264928 700062
rect 267660 699786 267688 703520
rect 269028 700256 269080 700262
rect 269028 700198 269080 700204
rect 267648 699780 267700 699786
rect 267648 699722 267700 699728
rect 269040 643906 269068 700198
rect 281448 699916 281500 699922
rect 281448 699858 281500 699864
rect 277308 699848 277360 699854
rect 277308 699790 277360 699796
rect 272892 648100 272944 648106
rect 272892 648042 272944 648048
rect 268686 643878 269068 643906
rect 272904 643892 272932 648042
rect 277320 643906 277348 699790
rect 281460 643906 281488 699858
rect 283852 699718 283880 703520
rect 288440 699780 288492 699786
rect 288440 699722 288492 699728
rect 283840 699712 283892 699718
rect 283840 699654 283892 699660
rect 285496 648236 285548 648242
rect 285496 648178 285548 648184
rect 277058 643878 277348 643906
rect 281290 643878 281488 643906
rect 285508 643892 285536 648178
rect 288452 644042 288480 699722
rect 293960 699712 294012 699718
rect 293960 699654 294012 699660
rect 288452 644014 289308 644042
rect 171810 643754 172192 643770
rect 171810 643748 172204 643754
rect 171810 643742 172152 643748
rect 125782 643719 125784 643728
rect 125836 643719 125838 643728
rect 125784 643690 125836 643696
rect 213946 643742 215248 643770
rect 222410 643742 223528 643770
rect 226550 643742 227024 643770
rect 230782 643742 231808 643770
rect 239246 643742 240088 643770
rect 243386 643742 244228 643770
rect 251850 643742 252508 643770
rect 256082 643742 256648 643770
rect 264454 643742 264928 643770
rect 289280 643770 289308 644014
rect 293972 643892 294000 699654
rect 300136 688634 300164 703520
rect 318800 701004 318852 701010
rect 318800 700946 318852 700952
rect 314660 700936 314712 700942
rect 314660 700878 314712 700884
rect 310520 700188 310572 700194
rect 310520 700130 310572 700136
rect 302240 700052 302292 700058
rect 302240 699994 302292 700000
rect 299664 688628 299716 688634
rect 299664 688570 299716 688576
rect 300124 688628 300176 688634
rect 300124 688570 300176 688576
rect 299676 685930 299704 688570
rect 299584 685902 299704 685930
rect 299584 684486 299612 685902
rect 299572 684480 299624 684486
rect 299572 684422 299624 684428
rect 299756 666596 299808 666602
rect 299756 666538 299808 666544
rect 299768 659734 299796 666538
rect 299756 659728 299808 659734
rect 299756 659670 299808 659676
rect 299664 657008 299716 657014
rect 299584 656956 299664 656962
rect 299584 656950 299716 656956
rect 299584 656934 299704 656950
rect 299584 656878 299612 656934
rect 299572 656872 299624 656878
rect 299572 656814 299624 656820
rect 298100 648168 298152 648174
rect 298100 648110 298152 648116
rect 298112 643892 298140 648110
rect 302252 643906 302280 699994
rect 306380 699984 306432 699990
rect 306380 699926 306432 699932
rect 306392 643906 306420 699926
rect 310532 643906 310560 700130
rect 314672 643906 314700 700878
rect 318812 643906 318840 700946
rect 322940 700800 322992 700806
rect 322940 700742 322992 700748
rect 302252 643878 302358 643906
rect 306392 643878 306590 643906
rect 310532 643878 310822 643906
rect 314672 643878 314962 643906
rect 318812 643878 319194 643906
rect 322952 643770 322980 700742
rect 331220 700664 331272 700670
rect 331220 700606 331272 700612
rect 327080 700596 327132 700602
rect 327080 700538 327132 700544
rect 327092 643770 327120 700538
rect 331232 643770 331260 700606
rect 332520 699854 332548 703520
rect 335360 700460 335412 700466
rect 335360 700402 335412 700408
rect 332508 699848 332560 699854
rect 332508 699790 332560 699796
rect 335372 643770 335400 700402
rect 339498 700360 339554 700369
rect 339498 700295 339554 700304
rect 343640 700324 343692 700330
rect 339512 643770 339540 700295
rect 343640 700266 343692 700272
rect 343652 643770 343680 700266
rect 348804 699922 348832 703520
rect 364996 703474 365024 703520
rect 364996 703446 365116 703474
rect 348792 699916 348844 699922
rect 348792 699858 348844 699864
rect 365088 686089 365116 703446
rect 397472 700126 397500 703520
rect 413664 700262 413692 703520
rect 413652 700256 413704 700262
rect 413652 700198 413704 700204
rect 397460 700120 397512 700126
rect 397460 700062 397512 700068
rect 429856 688634 429884 703520
rect 462332 700874 462360 703520
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 478524 700738 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 700732 478564 700738
rect 478512 700674 478564 700680
rect 429384 688628 429436 688634
rect 429384 688570 429436 688576
rect 429844 688628 429896 688634
rect 429844 688570 429896 688576
rect 365074 686080 365130 686089
rect 365074 686015 365130 686024
rect 364522 685944 364578 685953
rect 429396 685930 429424 688570
rect 494900 686089 494928 703446
rect 527192 700534 527220 703520
rect 527180 700528 527232 700534
rect 527180 700470 527232 700476
rect 543476 700398 543504 703520
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 559668 688634 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 559104 688628 559156 688634
rect 559104 688570 559156 688576
rect 559656 688628 559708 688634
rect 559656 688570 559708 688576
rect 494886 686080 494942 686089
rect 494886 686015 494942 686024
rect 364522 685879 364578 685888
rect 429304 685902 429424 685930
rect 494242 685944 494298 685953
rect 347780 681760 347832 681766
rect 347780 681702 347832 681708
rect 347792 643770 347820 681702
rect 364536 678994 364564 685879
rect 429304 684486 429332 685902
rect 559116 685930 559144 688570
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 494242 685879 494298 685888
rect 559024 685902 559144 685930
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 429292 684480 429344 684486
rect 429292 684422 429344 684428
rect 494256 678994 494284 685879
rect 559024 684486 559052 685902
rect 580172 685850 580224 685856
rect 559012 684480 559064 684486
rect 559012 684422 559064 684428
rect 364352 678966 364564 678994
rect 494072 678966 494284 678994
rect 364352 676190 364380 678966
rect 494072 676190 494100 678966
rect 364340 676184 364392 676190
rect 364340 676126 364392 676132
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 356060 667956 356112 667962
rect 356060 667898 356112 667904
rect 351920 652792 351972 652798
rect 351920 652734 351972 652740
rect 351932 643770 351960 652734
rect 356072 643770 356100 667898
rect 364432 666596 364484 666602
rect 364432 666538 364484 666544
rect 429476 666596 429528 666602
rect 429476 666538 429528 666544
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 559196 666596 559248 666602
rect 559196 666538 559248 666544
rect 364444 659682 364472 666538
rect 429488 659682 429516 666538
rect 364444 659654 364564 659682
rect 364536 654158 364564 659654
rect 429304 659654 429516 659682
rect 494164 659682 494192 666538
rect 559208 659682 559236 666538
rect 494164 659654 494284 659682
rect 429304 656878 429332 659654
rect 429292 656872 429344 656878
rect 429292 656814 429344 656820
rect 494256 654158 494284 659654
rect 559024 659654 559236 659682
rect 559024 656878 559052 659654
rect 559012 656872 559064 656878
rect 559012 656814 559064 656820
rect 364340 654152 364392 654158
rect 364340 654094 364392 654100
rect 364524 654152 364576 654158
rect 364524 654094 364576 654100
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 364352 648106 364380 654094
rect 364340 648100 364392 648106
rect 364340 648042 364392 648048
rect 494072 647970 494100 654094
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 494060 647964 494112 647970
rect 494060 647906 494112 647912
rect 386604 647216 386656 647222
rect 386604 647158 386656 647164
rect 365536 647012 365588 647018
rect 365536 646954 365588 646960
rect 361304 644088 361356 644094
rect 361304 644030 361356 644036
rect 361316 643892 361344 644030
rect 365548 643892 365576 646954
rect 382372 646876 382424 646882
rect 382372 646818 382424 646824
rect 378140 645720 378192 645726
rect 378140 645662 378192 645668
rect 373540 644020 373592 644026
rect 373540 643962 373592 643968
rect 373552 643906 373580 643962
rect 373552 643878 373934 643906
rect 378152 643892 378180 645662
rect 382384 643892 382412 646818
rect 386616 645522 386644 647158
rect 407580 647148 407632 647154
rect 407580 647090 407632 647096
rect 386512 645516 386564 645522
rect 386512 645458 386564 645464
rect 386604 645516 386656 645522
rect 386604 645458 386656 645464
rect 386524 643892 386552 645458
rect 399208 645380 399260 645386
rect 399208 645322 399260 645328
rect 399220 643892 399248 645322
rect 407592 643892 407620 647090
rect 522672 647080 522724 647086
rect 522672 647022 522724 647028
rect 432880 646536 432932 646542
rect 432880 646478 432932 646484
rect 416044 645584 416096 645590
rect 416044 645526 416096 645532
rect 411812 645312 411864 645318
rect 411812 645254 411864 645260
rect 411824 643892 411852 645254
rect 416056 643892 416084 645526
rect 424416 645176 424468 645182
rect 424416 645118 424468 645124
rect 424428 643892 424456 645118
rect 432892 643892 432920 646478
rect 441252 646468 441304 646474
rect 441252 646410 441304 646416
rect 437020 645040 437072 645046
rect 437020 644982 437072 644988
rect 437032 643892 437060 644982
rect 441264 643892 441292 646410
rect 445484 646400 445536 646406
rect 445484 646342 445536 646348
rect 445496 643892 445524 646342
rect 458088 646332 458140 646338
rect 458088 646274 458140 646280
rect 449716 644904 449768 644910
rect 449716 644846 449768 644852
rect 449728 643892 449756 644846
rect 458100 643892 458128 646274
rect 466552 646264 466604 646270
rect 466552 646206 466604 646212
rect 462320 644768 462372 644774
rect 462320 644710 462372 644716
rect 462332 643892 462360 644710
rect 466564 643892 466592 646206
rect 470784 646196 470836 646202
rect 470784 646138 470836 646144
rect 470796 643892 470824 646138
rect 483388 646128 483440 646134
rect 483388 646070 483440 646076
rect 504454 646096 504510 646105
rect 479154 645960 479210 645969
rect 479154 645895 479210 645904
rect 474924 644700 474976 644706
rect 474924 644642 474976 644648
rect 474936 643892 474964 644642
rect 479168 643892 479196 645895
rect 483400 643892 483428 646070
rect 495992 646060 496044 646066
rect 504454 646031 504510 646040
rect 495992 646002 496044 646008
rect 491760 645992 491812 645998
rect 491760 645934 491812 645940
rect 487620 644632 487672 644638
rect 487620 644574 487672 644580
rect 487632 643892 487660 644574
rect 491772 643892 491800 645934
rect 496004 643892 496032 646002
rect 500224 644496 500276 644502
rect 500224 644438 500276 644444
rect 500236 643892 500264 644438
rect 504468 643892 504496 646031
rect 508596 645924 508648 645930
rect 508596 645866 508648 645872
rect 508608 643892 508636 645866
rect 522580 644972 522632 644978
rect 522580 644914 522632 644920
rect 522488 644836 522540 644842
rect 522488 644778 522540 644784
rect 512828 644564 512880 644570
rect 512828 644506 512880 644512
rect 512840 643892 512868 644506
rect 402980 643816 403032 643822
rect 289280 643742 289754 643770
rect 322952 643742 323426 643770
rect 327092 643742 327658 643770
rect 331232 643742 331798 643770
rect 335372 643742 336030 643770
rect 339512 643742 340262 643770
rect 343652 643742 344494 643770
rect 347792 643742 348634 643770
rect 351932 643742 352866 643770
rect 356072 643742 357098 643770
rect 403032 643764 403374 643770
rect 402980 643758 403374 643764
rect 402992 643742 403374 643758
rect 172152 643690 172204 643696
rect 117228 643680 117280 643686
rect 117070 643628 117228 643634
rect 121368 643680 121420 643686
rect 117070 643622 117280 643628
rect 121302 643628 121368 643634
rect 121302 643622 121420 643628
rect 117070 643606 117268 643622
rect 121302 643606 121408 643622
rect 419920 643618 420210 643634
rect 419908 643612 420210 643618
rect 419960 643606 420210 643612
rect 419908 643554 419960 643560
rect 96344 643544 96396 643550
rect 91862 643482 92152 643498
rect 96094 643492 96344 643498
rect 96094 643486 96396 643492
rect 91862 643476 92164 643482
rect 91862 643470 92112 643476
rect 96094 643470 96384 643486
rect 92112 643418 92164 643424
rect 79600 643408 79652 643414
rect 49974 643376 50030 643385
rect 45586 643346 45876 643362
rect 45586 643340 45888 643346
rect 45586 643334 45836 643340
rect 49726 643334 49974 643362
rect 75274 643376 75330 643385
rect 58190 643346 58480 643362
rect 58190 643340 58492 643346
rect 58190 643334 58440 643340
rect 49974 643311 50030 643320
rect 45836 643282 45888 643288
rect 75026 643334 75274 643362
rect 79258 643356 79600 643362
rect 87880 643408 87932 643414
rect 79258 643350 79652 643356
rect 87630 643356 87880 643362
rect 100482 643376 100538 643385
rect 87630 643350 87932 643356
rect 79258 643334 79640 643350
rect 87630 643334 87920 643350
rect 100234 643334 100482 643362
rect 75274 643311 75330 643320
rect 100482 643311 100538 643320
rect 205454 643376 205510 643385
rect 218426 643376 218482 643385
rect 205510 643334 205574 643362
rect 218178 643334 218426 643362
rect 205454 643311 205510 643320
rect 218426 643311 218482 643320
rect 369398 643376 369454 643385
rect 390558 643376 390614 643385
rect 369454 643334 369702 643362
rect 369398 643311 369454 643320
rect 394790 643376 394846 643385
rect 390614 643334 390770 643362
rect 390558 643311 390614 643320
rect 428462 643376 428518 643385
rect 394846 643334 395002 643362
rect 394790 643311 394846 643320
rect 453670 643376 453726 643385
rect 428518 643334 428674 643362
rect 428462 643311 428518 643320
rect 516690 643376 516746 643385
rect 453726 643334 453974 643362
rect 453670 643311 453726 643320
rect 520922 643376 520978 643385
rect 516746 643334 517086 643362
rect 516690 643311 516746 643320
rect 520978 643334 521318 643362
rect 522396 643340 522448 643346
rect 520922 643311 520978 643320
rect 58440 643282 58492 643288
rect 522396 643282 522448 643288
rect 522304 643204 522356 643210
rect 522304 643146 522356 643152
rect 522118 616856 522174 616865
rect 522118 616791 522174 616800
rect 522132 610201 522160 616791
rect 522118 610192 522174 610201
rect 522118 610127 522174 610136
rect 40684 367056 40736 367062
rect 40684 366998 40736 367004
rect 246132 44254 246698 44282
rect 42904 44118 44022 44146
rect 44284 44118 44942 44146
rect 45664 44118 45954 44146
rect 31668 42016 31720 42022
rect 31668 41958 31720 41964
rect 28908 41948 28960 41954
rect 28908 41890 28960 41896
rect 25504 35896 25556 35902
rect 25504 35838 25556 35844
rect 26700 5092 26752 5098
rect 26700 5034 26752 5040
rect 25504 4004 25556 4010
rect 25504 3946 25556 3952
rect 24308 3936 24360 3942
rect 24308 3878 24360 3884
rect 23112 2848 23164 2854
rect 23112 2790 23164 2796
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 21928 2502 22048 2530
rect 21928 480 21956 2502
rect 23124 480 23152 2790
rect 24320 480 24348 3878
rect 25516 480 25544 3946
rect 26712 480 26740 5034
rect 28920 3738 28948 41890
rect 31680 38622 31708 41958
rect 38476 41880 38528 41886
rect 38476 41822 38528 41828
rect 35808 41812 35860 41818
rect 35808 41754 35860 41760
rect 31668 38616 31720 38622
rect 31668 38558 31720 38564
rect 31668 29028 31720 29034
rect 31668 28970 31720 28976
rect 31680 19310 31708 28970
rect 31484 19304 31536 19310
rect 31484 19246 31536 19252
rect 31668 19304 31720 19310
rect 31668 19246 31720 19252
rect 31496 9761 31524 19246
rect 31482 9752 31538 9761
rect 31482 9687 31538 9696
rect 31666 9752 31722 9761
rect 31666 9687 31722 9696
rect 31680 9654 31708 9687
rect 31668 9648 31720 9654
rect 31668 9590 31720 9596
rect 33876 5228 33928 5234
rect 33876 5170 33928 5176
rect 30288 5160 30340 5166
rect 30288 5102 30340 5108
rect 29092 4072 29144 4078
rect 29092 4014 29144 4020
rect 27896 3732 27948 3738
rect 27896 3674 27948 3680
rect 28908 3732 28960 3738
rect 28908 3674 28960 3680
rect 27908 480 27936 3674
rect 29104 480 29132 4014
rect 30300 480 30328 5102
rect 32680 3732 32732 3738
rect 32680 3674 32732 3680
rect 31484 604 31536 610
rect 31484 546 31536 552
rect 31496 480 31524 546
rect 32692 480 32720 3674
rect 33888 480 33916 5170
rect 35820 3398 35848 41754
rect 37372 5296 37424 5302
rect 37372 5238 37424 5244
rect 36176 4140 36228 4146
rect 36176 4082 36228 4088
rect 34980 3392 35032 3398
rect 34980 3334 35032 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 34992 480 35020 3334
rect 36188 480 36216 4082
rect 37384 480 37412 5238
rect 38488 626 38516 41822
rect 42708 41744 42760 41750
rect 42708 41686 42760 41692
rect 41328 41608 41380 41614
rect 41328 41550 41380 41556
rect 39304 41472 39356 41478
rect 39304 41414 39356 41420
rect 39316 4078 39344 41414
rect 39304 4072 39356 4078
rect 39304 4014 39356 4020
rect 39764 3800 39816 3806
rect 39764 3742 39816 3748
rect 38488 598 38608 626
rect 38580 480 38608 598
rect 39776 480 39804 3742
rect 41340 610 41368 41550
rect 42720 3330 42748 41686
rect 42904 3466 42932 44118
rect 44086 42120 44142 42129
rect 44086 42055 44142 42064
rect 44100 3534 44128 42055
rect 43352 3528 43404 3534
rect 43352 3470 43404 3476
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 42892 3460 42944 3466
rect 42892 3402 42944 3408
rect 42156 3324 42208 3330
rect 42156 3266 42208 3272
rect 42708 3324 42760 3330
rect 42708 3266 42760 3272
rect 40960 604 41012 610
rect 40960 546 41012 552
rect 41328 604 41380 610
rect 41328 546 41380 552
rect 40972 480 41000 546
rect 42168 480 42196 3266
rect 43364 480 43392 3470
rect 44284 3262 44312 44118
rect 45468 41676 45520 41682
rect 45468 41618 45520 41624
rect 45480 3534 45508 41618
rect 45664 3670 45692 44118
rect 46860 42158 46888 44132
rect 46848 42152 46900 42158
rect 46848 42094 46900 42100
rect 46940 42152 46992 42158
rect 46940 42094 46992 42100
rect 46952 41970 46980 42094
rect 47872 42090 47900 44132
rect 47860 42084 47912 42090
rect 47860 42026 47912 42032
rect 46860 41942 46980 41970
rect 46204 41540 46256 41546
rect 46204 41482 46256 41488
rect 45652 3664 45704 3670
rect 45652 3606 45704 3612
rect 46216 3602 46244 41482
rect 46204 3596 46256 3602
rect 46204 3538 46256 3544
rect 46860 3534 46888 41942
rect 48884 41546 48912 44132
rect 49608 42084 49660 42090
rect 49608 42026 49660 42032
rect 48872 41540 48924 41546
rect 48872 41482 48924 41488
rect 46940 3596 46992 3602
rect 46940 3538 46992 3544
rect 44548 3528 44600 3534
rect 44548 3470 44600 3476
rect 45468 3528 45520 3534
rect 45468 3470 45520 3476
rect 45744 3528 45796 3534
rect 45744 3470 45796 3476
rect 46848 3528 46900 3534
rect 46848 3470 46900 3476
rect 44272 3256 44324 3262
rect 44272 3198 44324 3204
rect 44560 480 44588 3470
rect 45756 480 45784 3470
rect 46952 480 46980 3538
rect 48136 3392 48188 3398
rect 48136 3334 48188 3340
rect 48148 480 48176 3334
rect 49620 626 49648 42026
rect 49804 4826 49832 44132
rect 50816 42498 50844 44132
rect 50804 42492 50856 42498
rect 50804 42434 50856 42440
rect 50988 42492 51040 42498
rect 50988 42434 51040 42440
rect 50344 41540 50396 41546
rect 50344 41482 50396 41488
rect 49792 4820 49844 4826
rect 49792 4762 49844 4768
rect 50356 3874 50384 41482
rect 50344 3868 50396 3874
rect 50344 3810 50396 3816
rect 51000 3534 51028 42434
rect 51828 42226 51856 44132
rect 52748 42294 52776 44132
rect 53392 44118 53774 44146
rect 52736 42288 52788 42294
rect 52736 42230 52788 42236
rect 51816 42220 51868 42226
rect 51816 42162 51868 42168
rect 53392 38622 53420 44118
rect 54772 42430 54800 44132
rect 54760 42424 54812 42430
rect 54760 42366 54812 42372
rect 55128 42424 55180 42430
rect 55128 42366 55180 42372
rect 53748 42220 53800 42226
rect 53748 42162 53800 42168
rect 53380 38616 53432 38622
rect 53380 38558 53432 38564
rect 53288 29028 53340 29034
rect 53288 28970 53340 28976
rect 53300 22166 53328 28970
rect 52552 22160 52604 22166
rect 52552 22102 52604 22108
rect 53288 22160 53340 22166
rect 53288 22102 53340 22108
rect 52564 12458 52592 22102
rect 52564 12430 52684 12458
rect 52656 4894 52684 12430
rect 52644 4888 52696 4894
rect 52644 4830 52696 4836
rect 50528 3528 50580 3534
rect 50528 3470 50580 3476
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 51632 3528 51684 3534
rect 51632 3470 51684 3476
rect 49344 598 49648 626
rect 49344 480 49372 598
rect 50540 480 50568 3470
rect 51644 480 51672 3470
rect 53760 3466 53788 42162
rect 55140 4146 55168 42366
rect 55692 41546 55720 44132
rect 56704 42362 56732 44132
rect 57440 44118 57730 44146
rect 56692 42356 56744 42362
rect 56692 42298 56744 42304
rect 56508 42288 56560 42294
rect 56508 42230 56560 42236
rect 55680 41540 55732 41546
rect 55680 41482 55732 41488
rect 54024 4140 54076 4146
rect 54024 4082 54076 4088
rect 55128 4140 55180 4146
rect 55128 4082 55180 4088
rect 52828 3460 52880 3466
rect 52828 3402 52880 3408
rect 53748 3460 53800 3466
rect 53748 3402 53800 3408
rect 52840 480 52868 3402
rect 54036 480 54064 4082
rect 55220 3868 55272 3874
rect 55220 3810 55272 3816
rect 55232 480 55260 3810
rect 56520 3670 56548 42230
rect 57244 41540 57296 41546
rect 57244 41482 57296 41488
rect 56876 31816 56928 31822
rect 56876 31758 56928 31764
rect 56888 12458 56916 31758
rect 56704 12430 56916 12458
rect 56704 4962 56732 12430
rect 56692 4956 56744 4962
rect 56692 4898 56744 4904
rect 57256 4010 57284 41482
rect 57440 31822 57468 44118
rect 58636 42634 58664 44132
rect 58624 42628 58676 42634
rect 58624 42570 58676 42576
rect 59648 42566 59676 44132
rect 60568 42770 60596 44132
rect 60752 44118 61594 44146
rect 60556 42764 60608 42770
rect 60556 42706 60608 42712
rect 60648 42628 60700 42634
rect 60648 42570 60700 42576
rect 59636 42560 59688 42566
rect 59636 42502 59688 42508
rect 57888 42356 57940 42362
rect 57888 42298 57940 42304
rect 57428 31816 57480 31822
rect 57428 31758 57480 31764
rect 57244 4004 57296 4010
rect 57244 3946 57296 3952
rect 56508 3664 56560 3670
rect 56508 3606 56560 3612
rect 57900 2854 57928 42298
rect 59912 42084 59964 42090
rect 59912 42026 59964 42032
rect 59924 41954 59952 42026
rect 59912 41948 59964 41954
rect 59912 41890 59964 41896
rect 60004 41472 60056 41478
rect 60004 41414 60056 41420
rect 60016 4298 60044 41414
rect 59924 4270 60044 4298
rect 59924 3942 59952 4270
rect 60660 4146 60688 42570
rect 60752 5030 60780 44118
rect 62592 42702 62620 44132
rect 62580 42696 62632 42702
rect 62580 42638 62632 42644
rect 62028 42356 62080 42362
rect 62028 42298 62080 42304
rect 60740 5024 60792 5030
rect 60740 4966 60792 4972
rect 60004 4140 60056 4146
rect 60004 4082 60056 4088
rect 60648 4140 60700 4146
rect 60648 4082 60700 4088
rect 59912 3936 59964 3942
rect 59912 3878 59964 3884
rect 58808 3664 58860 3670
rect 58808 3606 58860 3612
rect 57888 2848 57940 2854
rect 57888 2790 57940 2796
rect 56416 604 56468 610
rect 56416 546 56468 552
rect 57612 604 57664 610
rect 57612 546 57664 552
rect 56428 480 56456 546
rect 57624 480 57652 546
rect 58820 480 58848 3606
rect 60016 480 60044 4082
rect 62040 3466 62068 42298
rect 63512 41478 63540 44132
rect 64524 41546 64552 44132
rect 64892 44118 65550 44146
rect 66272 44118 66470 44146
rect 64788 42696 64840 42702
rect 64788 42638 64840 42644
rect 64512 41540 64564 41546
rect 64512 41482 64564 41488
rect 63500 41472 63552 41478
rect 63500 41414 63552 41420
rect 62396 3936 62448 3942
rect 62396 3878 62448 3884
rect 61200 3460 61252 3466
rect 61200 3402 61252 3408
rect 62028 3460 62080 3466
rect 62028 3402 62080 3408
rect 61212 480 61240 3402
rect 62408 480 62436 3878
rect 64800 3466 64828 42638
rect 64892 5098 64920 44118
rect 66168 42560 66220 42566
rect 66272 42514 66300 44118
rect 67468 42770 67496 44132
rect 67652 44118 68494 44146
rect 69032 44118 69414 44146
rect 67456 42764 67508 42770
rect 67456 42706 67508 42712
rect 66220 42508 66300 42514
rect 66168 42502 66300 42508
rect 66180 42486 66300 42502
rect 66904 41812 66956 41818
rect 66904 41754 66956 41760
rect 64880 5092 64932 5098
rect 64880 5034 64932 5040
rect 65984 4004 66036 4010
rect 65984 3946 66036 3952
rect 63592 3460 63644 3466
rect 63592 3402 63644 3408
rect 64788 3460 64840 3466
rect 64788 3402 64840 3408
rect 63604 480 63632 3402
rect 64788 3120 64840 3126
rect 64788 3062 64840 3068
rect 64800 480 64828 3062
rect 65996 480 66024 3946
rect 66916 3126 66944 41754
rect 67548 41472 67600 41478
rect 67548 41414 67600 41420
rect 66904 3120 66956 3126
rect 66904 3062 66956 3068
rect 67560 626 67588 41414
rect 67652 5166 67680 44118
rect 69032 42838 69060 44118
rect 69020 42832 69072 42838
rect 69020 42774 69072 42780
rect 68928 42764 68980 42770
rect 68928 42706 68980 42712
rect 68284 41608 68336 41614
rect 68284 41550 68336 41556
rect 67640 5160 67692 5166
rect 67640 5102 67692 5108
rect 68296 4078 68324 41550
rect 68284 4072 68336 4078
rect 68284 4014 68336 4020
rect 68940 3466 68968 42706
rect 69480 4072 69532 4078
rect 69480 4014 69532 4020
rect 68284 3460 68336 3466
rect 68284 3402 68336 3408
rect 68928 3460 68980 3466
rect 68928 3402 68980 3408
rect 67192 598 67588 626
rect 67192 480 67220 598
rect 68296 480 68324 3402
rect 69492 480 69520 4014
rect 70412 3738 70440 44132
rect 70504 44118 71438 44146
rect 70504 5234 70532 44118
rect 72344 42634 72372 44132
rect 72332 42628 72384 42634
rect 72332 42570 72384 42576
rect 73356 41614 73384 44132
rect 73344 41608 73396 41614
rect 73344 41550 73396 41556
rect 73804 41608 73856 41614
rect 73804 41550 73856 41556
rect 71688 41472 71740 41478
rect 71688 41414 71740 41420
rect 70492 5228 70544 5234
rect 70492 5170 70544 5176
rect 70400 3732 70452 3738
rect 70400 3674 70452 3680
rect 71700 3262 71728 41414
rect 73434 38720 73490 38729
rect 73490 38678 73568 38706
rect 73434 38655 73490 38664
rect 73540 38622 73568 38678
rect 73528 38616 73580 38622
rect 73528 38558 73580 38564
rect 73620 29028 73672 29034
rect 73620 28970 73672 28976
rect 73632 22114 73660 28970
rect 73448 22086 73660 22114
rect 73448 12458 73476 22086
rect 73264 12430 73476 12458
rect 73264 5302 73292 12430
rect 73252 5296 73304 5302
rect 73252 5238 73304 5244
rect 73068 4820 73120 4826
rect 73068 4762 73120 4768
rect 71872 4140 71924 4146
rect 71872 4082 71924 4088
rect 70676 3256 70728 3262
rect 70676 3198 70728 3204
rect 71688 3256 71740 3262
rect 71688 3198 71740 3204
rect 70688 480 70716 3198
rect 71884 480 71912 4082
rect 73080 480 73108 4762
rect 73816 4146 73844 41550
rect 74368 38865 74396 44132
rect 75288 41886 75316 44132
rect 76116 44118 76314 44146
rect 75828 42016 75880 42022
rect 75828 41958 75880 41964
rect 75276 41880 75328 41886
rect 75276 41822 75328 41828
rect 74448 41812 74500 41818
rect 74448 41754 74500 41760
rect 74354 38856 74410 38865
rect 74354 38791 74410 38800
rect 73804 4140 73856 4146
rect 73804 4082 73856 4088
rect 74460 610 74488 41754
rect 75840 38622 75868 41958
rect 75736 38616 75788 38622
rect 75736 38558 75788 38564
rect 75828 38616 75880 38622
rect 75828 38558 75880 38564
rect 75748 37262 75776 38558
rect 75736 37256 75788 37262
rect 75736 37198 75788 37204
rect 75828 27668 75880 27674
rect 75828 27610 75880 27616
rect 75840 21010 75868 27610
rect 75828 21004 75880 21010
rect 75828 20946 75880 20952
rect 75460 9716 75512 9722
rect 75460 9658 75512 9664
rect 74264 604 74316 610
rect 74264 546 74316 552
rect 74448 604 74500 610
rect 74448 546 74500 552
rect 74276 480 74304 546
rect 75472 480 75500 9658
rect 76116 3806 76144 44118
rect 77220 41886 77248 44132
rect 77208 41880 77260 41886
rect 77208 41822 77260 41828
rect 78232 41750 78260 44132
rect 79244 42129 79272 44132
rect 79230 42120 79286 42129
rect 79230 42055 79286 42064
rect 78588 41880 78640 41886
rect 78588 41822 78640 41828
rect 78220 41744 78272 41750
rect 78220 41686 78272 41692
rect 76104 3800 76156 3806
rect 76104 3742 76156 3748
rect 76656 3732 76708 3738
rect 76656 3674 76708 3680
rect 76668 480 76696 3674
rect 78600 3194 78628 41822
rect 79968 41744 80020 41750
rect 79968 41686 80020 41692
rect 79980 3806 80008 41686
rect 80164 41682 80192 44132
rect 81176 42158 81204 44132
rect 81164 42152 81216 42158
rect 81164 42094 81216 42100
rect 80152 41676 80204 41682
rect 80152 41618 80204 41624
rect 82188 41546 82216 44132
rect 83016 44118 83122 44146
rect 83384 44118 84134 44146
rect 82728 42152 82780 42158
rect 82728 42094 82780 42100
rect 80704 41540 80756 41546
rect 80704 41482 80756 41488
rect 82176 41540 82228 41546
rect 82176 41482 82228 41488
rect 80716 4146 80744 41482
rect 80704 4140 80756 4146
rect 80704 4082 80756 4088
rect 82636 3868 82688 3874
rect 82636 3810 82688 3816
rect 79048 3800 79100 3806
rect 79048 3742 79100 3748
rect 79968 3800 80020 3806
rect 79968 3742 80020 3748
rect 80244 3800 80296 3806
rect 80244 3742 80296 3748
rect 77852 3188 77904 3194
rect 77852 3130 77904 3136
rect 78588 3188 78640 3194
rect 78588 3130 78640 3136
rect 77864 480 77892 3130
rect 79060 480 79088 3742
rect 80256 480 80284 3742
rect 81440 3460 81492 3466
rect 81440 3402 81492 3408
rect 81452 480 81480 3402
rect 82648 480 82676 3810
rect 82740 3466 82768 42094
rect 82728 3460 82780 3466
rect 82728 3402 82780 3408
rect 83016 3398 83044 44118
rect 83384 41682 83412 44118
rect 85132 42090 85160 44132
rect 85684 44118 86066 44146
rect 85120 42084 85172 42090
rect 85120 42026 85172 42032
rect 85488 42084 85540 42090
rect 85488 42026 85540 42032
rect 83372 41676 83424 41682
rect 83372 41618 83424 41624
rect 83464 41676 83516 41682
rect 83464 41618 83516 41624
rect 83476 3874 83504 41618
rect 85500 4146 85528 42026
rect 84936 4140 84988 4146
rect 84936 4082 84988 4088
rect 85488 4140 85540 4146
rect 85488 4082 85540 4088
rect 83464 3868 83516 3874
rect 83464 3810 83516 3816
rect 83004 3392 83056 3398
rect 83004 3334 83056 3340
rect 83832 3324 83884 3330
rect 83832 3266 83884 3272
rect 83844 480 83872 3266
rect 84948 480 84976 4082
rect 85684 3398 85712 44118
rect 87064 42226 87092 44132
rect 88076 42430 88104 44132
rect 88352 44118 89010 44146
rect 88064 42424 88116 42430
rect 88064 42366 88116 42372
rect 87052 42220 87104 42226
rect 87052 42162 87104 42168
rect 86868 41540 86920 41546
rect 86868 41482 86920 41488
rect 86880 4146 86908 41482
rect 86132 4140 86184 4146
rect 86132 4082 86184 4088
rect 86868 4140 86920 4146
rect 86868 4082 86920 4088
rect 85672 3392 85724 3398
rect 85672 3334 85724 3340
rect 86144 480 86172 4082
rect 88352 3602 88380 44118
rect 89628 42424 89680 42430
rect 89628 42366 89680 42372
rect 88340 3596 88392 3602
rect 88340 3538 88392 3544
rect 87328 3392 87380 3398
rect 87328 3334 87380 3340
rect 87340 480 87368 3334
rect 89640 3194 89668 42366
rect 90008 42294 90036 44132
rect 91020 42498 91048 44132
rect 91112 44118 91954 44146
rect 91008 42492 91060 42498
rect 91008 42434 91060 42440
rect 89996 42288 90048 42294
rect 89996 42230 90048 42236
rect 91008 42220 91060 42226
rect 91008 42162 91060 42168
rect 91020 3602 91048 42162
rect 91112 3670 91140 44118
rect 92952 42566 92980 44132
rect 92940 42560 92992 42566
rect 92940 42502 92992 42508
rect 92388 42492 92440 42498
rect 92388 42434 92440 42440
rect 91100 3664 91152 3670
rect 91100 3606 91152 3612
rect 89720 3596 89772 3602
rect 89720 3538 89772 3544
rect 91008 3596 91060 3602
rect 91008 3538 91060 3544
rect 88524 3188 88576 3194
rect 88524 3130 88576 3136
rect 89628 3188 89680 3194
rect 89628 3130 89680 3136
rect 88536 480 88564 3130
rect 89732 480 89760 3538
rect 90916 3528 90968 3534
rect 90916 3470 90968 3476
rect 90928 480 90956 3470
rect 92400 2854 92428 42434
rect 93872 42362 93900 44132
rect 93964 44118 94898 44146
rect 93860 42356 93912 42362
rect 93860 42298 93912 42304
rect 93768 42288 93820 42294
rect 93768 42230 93820 42236
rect 93780 4146 93808 42230
rect 93308 4140 93360 4146
rect 93308 4082 93360 4088
rect 93768 4140 93820 4146
rect 93768 4082 93820 4088
rect 92112 2848 92164 2854
rect 92112 2790 92164 2796
rect 92388 2848 92440 2854
rect 92388 2790 92440 2796
rect 92124 480 92152 2790
rect 93320 480 93348 4082
rect 93964 3942 93992 44118
rect 95896 42702 95924 44132
rect 95884 42696 95936 42702
rect 95884 42638 95936 42644
rect 96528 42560 96580 42566
rect 96528 42502 96580 42508
rect 93952 3936 94004 3942
rect 93952 3878 94004 3884
rect 94504 3664 94556 3670
rect 94504 3606 94556 3612
rect 94516 480 94544 3606
rect 96540 3262 96568 42502
rect 96816 41954 96844 44132
rect 97552 44118 97842 44146
rect 96804 41948 96856 41954
rect 96804 41890 96856 41896
rect 97552 29034 97580 44118
rect 98840 42770 98868 44132
rect 98828 42764 98880 42770
rect 98828 42706 98880 42712
rect 99288 42696 99340 42702
rect 99288 42638 99340 42644
rect 97908 42356 97960 42362
rect 97908 42298 97960 42304
rect 96620 29028 96672 29034
rect 96620 28970 96672 28976
rect 97540 29028 97592 29034
rect 97540 28970 97592 28976
rect 96632 19378 96660 28970
rect 96620 19372 96672 19378
rect 96620 19314 96672 19320
rect 96712 19372 96764 19378
rect 96712 19314 96764 19320
rect 96724 19258 96752 19314
rect 96724 19230 96844 19258
rect 96816 4010 96844 19230
rect 97920 4146 97948 42298
rect 96896 4140 96948 4146
rect 96896 4082 96948 4088
rect 97908 4140 97960 4146
rect 97908 4082 97960 4088
rect 96804 4004 96856 4010
rect 96804 3946 96856 3952
rect 95700 3256 95752 3262
rect 95700 3198 95752 3204
rect 96528 3256 96580 3262
rect 96528 3198 96580 3204
rect 95712 480 95740 3198
rect 96908 480 96936 4082
rect 98092 3936 98144 3942
rect 98092 3878 98144 3884
rect 98104 480 98132 3878
rect 99300 480 99328 42638
rect 99760 42634 99788 44132
rect 100786 44118 100892 44146
rect 99748 42628 99800 42634
rect 99748 42570 99800 42576
rect 100666 42120 100722 42129
rect 100666 42055 100722 42064
rect 100680 19582 100708 42055
rect 100668 19576 100720 19582
rect 100668 19518 100720 19524
rect 100668 19440 100720 19446
rect 100668 19382 100720 19388
rect 100680 9654 100708 19382
rect 100668 9648 100720 9654
rect 100668 9590 100720 9596
rect 100864 4078 100892 44118
rect 101784 41478 101812 44132
rect 102704 41614 102732 44132
rect 103624 44118 103730 44146
rect 102692 41608 102744 41614
rect 102692 41550 102744 41556
rect 103428 41608 103480 41614
rect 103428 41550 103480 41556
rect 101772 41472 101824 41478
rect 101772 41414 101824 41420
rect 103440 4146 103468 41550
rect 103624 4826 103652 44118
rect 104728 41818 104756 44132
rect 105648 42022 105676 44132
rect 106292 44118 106674 44146
rect 105636 42016 105688 42022
rect 105636 41958 105688 41964
rect 104808 41948 104860 41954
rect 104808 41890 104860 41896
rect 104716 41812 104768 41818
rect 104716 41754 104768 41760
rect 103612 4820 103664 4826
rect 103612 4762 103664 4768
rect 102784 4140 102836 4146
rect 102784 4082 102836 4088
rect 103428 4140 103480 4146
rect 103428 4082 103480 4088
rect 100852 4072 100904 4078
rect 100852 4014 100904 4020
rect 101588 3868 101640 3874
rect 101588 3810 101640 3816
rect 100484 604 100536 610
rect 100484 546 100536 552
rect 100496 480 100524 546
rect 101600 480 101628 3810
rect 102796 480 102824 4082
rect 104820 3194 104848 41890
rect 106188 41812 106240 41818
rect 106188 41754 106240 41760
rect 106200 3466 106228 41754
rect 106292 3738 106320 44118
rect 107568 42764 107620 42770
rect 107568 42706 107620 42712
rect 107476 42628 107528 42634
rect 107476 42570 107528 42576
rect 107488 4146 107516 42570
rect 106372 4140 106424 4146
rect 106372 4082 106424 4088
rect 107476 4140 107528 4146
rect 107476 4082 107528 4088
rect 106280 3732 106332 3738
rect 106280 3674 106332 3680
rect 105176 3460 105228 3466
rect 105176 3402 105228 3408
rect 106188 3460 106240 3466
rect 106188 3402 106240 3408
rect 103980 3188 104032 3194
rect 103980 3130 104032 3136
rect 104808 3188 104860 3194
rect 104808 3130 104860 3136
rect 103992 480 104020 3130
rect 105188 480 105216 3402
rect 106384 480 106412 4082
rect 107580 480 107608 42706
rect 107672 41886 107700 44132
rect 107660 41880 107712 41886
rect 107660 41822 107712 41828
rect 108592 41750 108620 44132
rect 109052 44118 109618 44146
rect 108580 41744 108632 41750
rect 108580 41686 108632 41692
rect 108948 38684 109000 38690
rect 108948 38626 109000 38632
rect 108960 38554 108988 38626
rect 108948 38548 109000 38554
rect 108948 38490 109000 38496
rect 108948 29028 109000 29034
rect 108948 28970 109000 28976
rect 108960 19310 108988 28970
rect 108764 19304 108816 19310
rect 108764 19246 108816 19252
rect 108948 19304 109000 19310
rect 108948 19246 109000 19252
rect 108776 9761 108804 19246
rect 108762 9752 108818 9761
rect 108762 9687 108818 9696
rect 108946 9752 109002 9761
rect 108946 9687 109002 9696
rect 108960 9654 108988 9687
rect 108948 9648 109000 9654
rect 108948 9590 109000 9596
rect 109052 3806 109080 44118
rect 110524 42158 110552 44132
rect 110512 42152 110564 42158
rect 110512 42094 110564 42100
rect 110328 41880 110380 41886
rect 110328 41822 110380 41828
rect 109040 3800 109092 3806
rect 109040 3742 109092 3748
rect 110340 2854 110368 41822
rect 111536 41682 111564 44132
rect 111904 44118 112562 44146
rect 111524 41676 111576 41682
rect 111524 41618 111576 41624
rect 111708 41676 111760 41682
rect 111708 41618 111760 41624
rect 111720 4146 111748 41618
rect 111156 4140 111208 4146
rect 111156 4082 111208 4088
rect 111708 4140 111760 4146
rect 111708 4082 111760 4088
rect 109960 2848 110012 2854
rect 109960 2790 110012 2796
rect 110328 2848 110380 2854
rect 110328 2790 110380 2796
rect 108764 604 108816 610
rect 108764 546 108816 552
rect 108776 480 108804 546
rect 109972 480 110000 2790
rect 111168 480 111196 4082
rect 111904 3398 111932 44118
rect 113468 42090 113496 44132
rect 114112 44118 114494 44146
rect 114664 44118 115506 44146
rect 113456 42084 113508 42090
rect 113456 42026 113508 42032
rect 114112 41546 114140 44118
rect 114100 41540 114152 41546
rect 114100 41482 114152 41488
rect 114468 41540 114520 41546
rect 114468 41482 114520 41488
rect 113088 41472 113140 41478
rect 113088 41414 113140 41420
rect 113100 4146 113128 41414
rect 114480 4146 114508 41482
rect 112352 4140 112404 4146
rect 112352 4082 112404 4088
rect 113088 4140 113140 4146
rect 113088 4082 113140 4088
rect 113548 4140 113600 4146
rect 113548 4082 113600 4088
rect 114468 4140 114520 4146
rect 114468 4082 114520 4088
rect 111892 3392 111944 3398
rect 111892 3334 111944 3340
rect 112364 480 112392 4082
rect 113560 480 113588 4082
rect 114664 3534 114692 44118
rect 116412 42430 116440 44132
rect 116400 42424 116452 42430
rect 116400 42366 116452 42372
rect 117424 42226 117452 44132
rect 118160 44118 118450 44146
rect 117412 42220 117464 42226
rect 117412 42162 117464 42168
rect 117136 42152 117188 42158
rect 117136 42094 117188 42100
rect 115848 41744 115900 41750
rect 115848 41686 115900 41692
rect 115860 3534 115888 41686
rect 115940 4140 115992 4146
rect 115940 4082 115992 4088
rect 114652 3528 114704 3534
rect 114652 3470 114704 3476
rect 114744 3528 114796 3534
rect 114744 3470 114796 3476
rect 115848 3528 115900 3534
rect 115848 3470 115900 3476
rect 114756 480 114784 3470
rect 115952 480 115980 4082
rect 117148 480 117176 42094
rect 117228 42084 117280 42090
rect 117228 42026 117280 42032
rect 117240 4146 117268 42026
rect 118160 29209 118188 44118
rect 119356 42498 119384 44132
rect 119344 42492 119396 42498
rect 119344 42434 119396 42440
rect 119988 42424 120040 42430
rect 119988 42366 120040 42372
rect 118608 42152 118660 42158
rect 118608 42094 118660 42100
rect 118146 29200 118202 29209
rect 118146 29135 118202 29144
rect 117410 29064 117466 29073
rect 117410 28999 117466 29008
rect 117424 27606 117452 28999
rect 117412 27600 117464 27606
rect 117412 27542 117464 27548
rect 117688 9716 117740 9722
rect 117688 9658 117740 9664
rect 117228 4140 117280 4146
rect 117228 4082 117280 4088
rect 117700 3602 117728 9658
rect 117688 3596 117740 3602
rect 117688 3538 117740 3544
rect 118620 2854 118648 42094
rect 120000 4146 120028 42366
rect 120368 42294 120396 44132
rect 121104 44118 121394 44146
rect 120356 42288 120408 42294
rect 120356 42230 120408 42236
rect 121104 27849 121132 44118
rect 122300 42566 122328 44132
rect 122288 42560 122340 42566
rect 122288 42502 122340 42508
rect 121368 42492 121420 42498
rect 121368 42434 121420 42440
rect 121090 27840 121146 27849
rect 121090 27775 121146 27784
rect 120170 27704 120226 27713
rect 120170 27639 120226 27648
rect 120184 27606 120212 27639
rect 120172 27600 120224 27606
rect 120172 27542 120224 27548
rect 120448 12436 120500 12442
rect 120448 12378 120500 12384
rect 120460 4418 120488 12378
rect 120448 4412 120500 4418
rect 120448 4354 120500 4360
rect 119436 4140 119488 4146
rect 119436 4082 119488 4088
rect 119988 4140 120040 4146
rect 119988 4082 120040 4088
rect 118240 2848 118292 2854
rect 118240 2790 118292 2796
rect 118608 2848 118660 2854
rect 118608 2790 118660 2796
rect 118252 480 118280 2790
rect 119448 480 119476 4082
rect 121380 3398 121408 42434
rect 123312 42362 123340 44132
rect 123300 42356 123352 42362
rect 123300 42298 123352 42304
rect 122748 42288 122800 42294
rect 122748 42230 122800 42236
rect 122760 3738 122788 42230
rect 124128 41812 124180 41818
rect 124128 41754 124180 41760
rect 121828 3732 121880 3738
rect 121828 3674 121880 3680
rect 122748 3732 122800 3738
rect 122748 3674 122800 3680
rect 120632 3392 120684 3398
rect 120632 3334 120684 3340
rect 121368 3392 121420 3398
rect 121368 3334 121420 3340
rect 120644 480 120672 3334
rect 121840 480 121868 3674
rect 124140 3670 124168 41754
rect 124324 3942 124352 44132
rect 125244 42702 125272 44132
rect 125232 42696 125284 42702
rect 125232 42638 125284 42644
rect 125416 42356 125468 42362
rect 125416 42298 125468 42304
rect 125324 12436 125376 12442
rect 125324 12378 125376 12384
rect 124312 3936 124364 3942
rect 124312 3878 124364 3884
rect 123024 3664 123076 3670
rect 123024 3606 123076 3612
rect 124128 3664 124180 3670
rect 124128 3606 124180 3612
rect 123036 480 123064 3606
rect 124220 3188 124272 3194
rect 124220 3130 124272 3136
rect 124232 480 124260 3130
rect 125336 3074 125364 12378
rect 125428 3194 125456 42298
rect 125692 42220 125744 42226
rect 125692 42162 125744 42168
rect 125704 42106 125732 42162
rect 126256 42129 126284 44132
rect 127084 44118 127190 44146
rect 127544 44118 128202 44146
rect 125520 42078 125732 42106
rect 126242 42120 126298 42129
rect 125520 12442 125548 42078
rect 126242 42055 126298 42064
rect 125508 12436 125560 12442
rect 125508 12378 125560 12384
rect 127084 3874 127112 44118
rect 127544 41886 127572 44118
rect 129200 41954 129228 44132
rect 129648 42696 129700 42702
rect 129648 42638 129700 42644
rect 129188 41948 129240 41954
rect 129188 41890 129240 41896
rect 127532 41880 127584 41886
rect 127532 41822 127584 41828
rect 128268 41608 128320 41614
rect 128268 41550 128320 41556
rect 128280 4146 128308 41550
rect 127808 4140 127860 4146
rect 127808 4082 127860 4088
rect 128268 4140 128320 4146
rect 128268 4082 128320 4088
rect 127072 3868 127124 3874
rect 127072 3810 127124 3816
rect 126612 3460 126664 3466
rect 126612 3402 126664 3408
rect 125416 3188 125468 3194
rect 125416 3130 125468 3136
rect 125336 3046 125456 3074
rect 125428 480 125456 3046
rect 126624 480 126652 3402
rect 127820 480 127848 4082
rect 129660 3058 129688 42638
rect 130120 41682 130148 44132
rect 131132 42634 131160 44132
rect 131224 44118 132158 44146
rect 131224 42770 131252 44118
rect 131212 42764 131264 42770
rect 131212 42706 131264 42712
rect 131120 42628 131172 42634
rect 131120 42570 131172 42576
rect 133064 42022 133092 44132
rect 133788 42764 133840 42770
rect 133788 42706 133840 42712
rect 133052 42016 133104 42022
rect 133052 41958 133104 41964
rect 133696 42016 133748 42022
rect 133696 41958 133748 41964
rect 131028 41948 131080 41954
rect 131028 41890 131080 41896
rect 130108 41676 130160 41682
rect 130108 41618 130160 41624
rect 131040 3534 131068 41890
rect 132408 41676 132460 41682
rect 132408 41618 132460 41624
rect 132420 3534 132448 41618
rect 133708 3534 133736 41958
rect 130200 3528 130252 3534
rect 130200 3470 130252 3476
rect 131028 3528 131080 3534
rect 131028 3470 131080 3476
rect 131396 3528 131448 3534
rect 131396 3470 131448 3476
rect 132408 3528 132460 3534
rect 132408 3470 132460 3476
rect 132592 3528 132644 3534
rect 132592 3470 132644 3476
rect 133696 3528 133748 3534
rect 133696 3470 133748 3476
rect 129004 3052 129056 3058
rect 129004 2994 129056 3000
rect 129648 3052 129700 3058
rect 129648 2994 129700 3000
rect 129016 480 129044 2994
rect 130212 480 130240 3470
rect 131408 480 131436 3470
rect 132604 480 132632 3470
rect 133800 480 133828 42706
rect 134076 42702 134104 44132
rect 134064 42696 134116 42702
rect 134064 42638 134116 42644
rect 135088 41886 135116 44132
rect 135076 41880 135128 41886
rect 135076 41822 135128 41828
rect 135168 41880 135220 41886
rect 135168 41822 135220 41828
rect 135180 3482 135208 41822
rect 136008 41478 136036 44132
rect 137020 41546 137048 44132
rect 137928 41880 137980 41886
rect 137928 41822 137980 41828
rect 137008 41540 137060 41546
rect 137008 41482 137060 41488
rect 135996 41472 136048 41478
rect 135996 41414 136048 41420
rect 136548 41472 136600 41478
rect 136548 41414 136600 41420
rect 134904 3454 135208 3482
rect 134904 480 134932 3454
rect 136560 2922 136588 41414
rect 137940 3534 137968 41822
rect 138032 41750 138060 44132
rect 138952 42498 138980 44132
rect 138940 42492 138992 42498
rect 138940 42434 138992 42440
rect 139308 42492 139360 42498
rect 139308 42434 139360 42440
rect 138020 41744 138072 41750
rect 138020 41686 138072 41692
rect 139320 3534 139348 42434
rect 139964 42090 139992 44132
rect 140976 42158 141004 44132
rect 141896 42430 141924 44132
rect 142908 42566 142936 44132
rect 142896 42560 142948 42566
rect 142896 42502 142948 42508
rect 141884 42424 141936 42430
rect 141884 42366 141936 42372
rect 141976 42424 142028 42430
rect 141976 42366 142028 42372
rect 140964 42152 141016 42158
rect 140964 42094 141016 42100
rect 139952 42084 140004 42090
rect 139952 42026 140004 42032
rect 140688 41744 140740 41750
rect 140688 41686 140740 41692
rect 140700 3534 140728 41686
rect 141988 3534 142016 42366
rect 143828 42294 143856 44132
rect 144644 42560 144696 42566
rect 144644 42502 144696 42508
rect 143816 42288 143868 42294
rect 143816 42230 143868 42236
rect 143448 42152 143500 42158
rect 143448 42094 143500 42100
rect 142068 42084 142120 42090
rect 142068 42026 142120 42032
rect 137284 3528 137336 3534
rect 137284 3470 137336 3476
rect 137928 3528 137980 3534
rect 137928 3470 137980 3476
rect 138480 3528 138532 3534
rect 138480 3470 138532 3476
rect 139308 3528 139360 3534
rect 139308 3470 139360 3476
rect 139676 3528 139728 3534
rect 139676 3470 139728 3476
rect 140688 3528 140740 3534
rect 140688 3470 140740 3476
rect 140872 3528 140924 3534
rect 140872 3470 140924 3476
rect 141976 3528 142028 3534
rect 141976 3470 142028 3476
rect 136088 2916 136140 2922
rect 136088 2858 136140 2864
rect 136548 2916 136600 2922
rect 136548 2858 136600 2864
rect 136100 480 136128 2858
rect 137296 480 137324 3470
rect 138492 480 138520 3470
rect 139688 480 139716 3470
rect 140884 480 140912 3470
rect 142080 480 142108 42026
rect 143460 3346 143488 42094
rect 144656 39250 144684 42502
rect 144840 41818 144868 44132
rect 145852 42362 145880 44132
rect 145840 42356 145892 42362
rect 145840 42298 145892 42304
rect 146208 42288 146260 42294
rect 146208 42230 146260 42236
rect 144828 41812 144880 41818
rect 144828 41754 144880 41760
rect 144656 39222 144868 39250
rect 144840 3346 144868 39222
rect 146220 3534 146248 42230
rect 146772 42226 146800 44132
rect 146760 42220 146812 42226
rect 146760 42162 146812 42168
rect 147588 42220 147640 42226
rect 147588 42162 147640 42168
rect 147600 3534 147628 42162
rect 145656 3528 145708 3534
rect 145656 3470 145708 3476
rect 146208 3528 146260 3534
rect 146208 3470 146260 3476
rect 146852 3528 146904 3534
rect 146852 3470 146904 3476
rect 147588 3528 147640 3534
rect 147588 3470 147640 3476
rect 143276 3318 143488 3346
rect 144472 3318 144868 3346
rect 143276 480 143304 3318
rect 144472 480 144500 3318
rect 145668 480 145696 3470
rect 146864 480 146892 3470
rect 147784 3466 147812 44132
rect 148796 41614 148824 44132
rect 149716 42702 149744 44132
rect 149704 42696 149756 42702
rect 149704 42638 149756 42644
rect 150728 41954 150756 44132
rect 151464 44118 151754 44146
rect 150716 41948 150768 41954
rect 150716 41890 150768 41896
rect 148968 41812 149020 41818
rect 148968 41754 149020 41760
rect 148784 41608 148836 41614
rect 148784 41550 148836 41556
rect 148980 3534 149008 41754
rect 151464 41682 151492 44118
rect 151636 42696 151688 42702
rect 151636 42638 151688 42644
rect 151452 41676 151504 41682
rect 151452 41618 151504 41624
rect 150348 41608 150400 41614
rect 150348 41550 150400 41556
rect 150360 3534 150388 41550
rect 151648 3602 151676 42638
rect 151728 42356 151780 42362
rect 151728 42298 151780 42304
rect 150440 3596 150492 3602
rect 150440 3538 150492 3544
rect 151636 3596 151688 3602
rect 151636 3538 151688 3544
rect 148048 3528 148100 3534
rect 148048 3470 148100 3476
rect 148968 3528 149020 3534
rect 148968 3470 149020 3476
rect 149244 3528 149296 3534
rect 149244 3470 149296 3476
rect 150348 3528 150400 3534
rect 150348 3470 150400 3476
rect 147772 3460 147824 3466
rect 147772 3402 147824 3408
rect 148060 480 148088 3470
rect 149256 480 149284 3470
rect 150452 480 150480 3538
rect 151740 3482 151768 42298
rect 152660 42022 152688 44132
rect 153672 42770 153700 44132
rect 153660 42764 153712 42770
rect 153660 42706 153712 42712
rect 154488 42764 154540 42770
rect 154488 42706 154540 42712
rect 152648 42016 152700 42022
rect 152648 41958 152700 41964
rect 153108 42016 153160 42022
rect 153108 41958 153160 41964
rect 153120 3482 153148 41958
rect 154500 3534 154528 42706
rect 154684 42634 154712 44132
rect 154672 42628 154724 42634
rect 154672 42570 154724 42576
rect 155604 41478 155632 44132
rect 155868 42628 155920 42634
rect 155868 42570 155920 42576
rect 155592 41472 155644 41478
rect 155592 41414 155644 41420
rect 155880 3534 155908 42570
rect 156616 41886 156644 44132
rect 157628 42498 157656 44132
rect 157616 42492 157668 42498
rect 157616 42434 157668 42440
rect 156604 41880 156656 41886
rect 156604 41822 156656 41828
rect 157248 41880 157300 41886
rect 157248 41822 157300 41828
rect 157260 3534 157288 41822
rect 158548 41750 158576 44132
rect 158628 42492 158680 42498
rect 158628 42434 158680 42440
rect 158536 41744 158588 41750
rect 158536 41686 158588 41692
rect 151556 3454 151768 3482
rect 152752 3454 153148 3482
rect 153936 3528 153988 3534
rect 153936 3470 153988 3476
rect 154488 3528 154540 3534
rect 154488 3470 154540 3476
rect 155132 3528 155184 3534
rect 155132 3470 155184 3476
rect 155868 3528 155920 3534
rect 155868 3470 155920 3476
rect 156328 3528 156380 3534
rect 156328 3470 156380 3476
rect 157248 3528 157300 3534
rect 157248 3470 157300 3476
rect 151556 480 151584 3454
rect 152752 480 152780 3454
rect 153948 480 153976 3470
rect 155144 480 155172 3470
rect 156340 480 156368 3470
rect 158640 3330 158668 42434
rect 159560 42430 159588 44132
rect 159548 42424 159600 42430
rect 159548 42366 159600 42372
rect 159916 42424 159968 42430
rect 159916 42366 159968 42372
rect 159928 3602 159956 42366
rect 160480 42090 160508 44132
rect 161492 42158 161520 44132
rect 162504 42566 162532 44132
rect 162492 42560 162544 42566
rect 162492 42502 162544 42508
rect 163424 42294 163452 44132
rect 163412 42288 163464 42294
rect 163412 42230 163464 42236
rect 164436 42226 164464 44132
rect 164424 42220 164476 42226
rect 164424 42162 164476 42168
rect 161480 42152 161532 42158
rect 161480 42094 161532 42100
rect 164148 42152 164200 42158
rect 164148 42094 164200 42100
rect 160468 42084 160520 42090
rect 160468 42026 160520 42032
rect 162768 42084 162820 42090
rect 162768 42026 162820 42032
rect 160008 41948 160060 41954
rect 160008 41890 160060 41896
rect 158720 3596 158772 3602
rect 158720 3538 158772 3544
rect 159916 3596 159968 3602
rect 159916 3538 159968 3544
rect 157524 3324 157576 3330
rect 157524 3266 157576 3272
rect 158628 3324 158680 3330
rect 158628 3266 158680 3272
rect 157536 480 157564 3266
rect 158732 480 158760 3538
rect 160020 3482 160048 41890
rect 161388 41744 161440 41750
rect 161388 41686 161440 41692
rect 161400 3482 161428 41686
rect 162780 3534 162808 42026
rect 164160 3534 164188 42094
rect 165448 41818 165476 44132
rect 165528 42288 165580 42294
rect 165528 42230 165580 42236
rect 165436 41812 165488 41818
rect 165436 41754 165488 41760
rect 159928 3454 160048 3482
rect 161124 3454 161428 3482
rect 162308 3528 162360 3534
rect 162308 3470 162360 3476
rect 162768 3528 162820 3534
rect 162768 3470 162820 3476
rect 163504 3528 163556 3534
rect 163504 3470 163556 3476
rect 164148 3528 164200 3534
rect 164148 3470 164200 3476
rect 159928 480 159956 3454
rect 161124 480 161152 3454
rect 162320 480 162348 3470
rect 163516 480 163544 3470
rect 165540 3466 165568 42230
rect 166368 41614 166396 44132
rect 167380 42702 167408 44132
rect 167368 42696 167420 42702
rect 167368 42638 167420 42644
rect 168288 42560 168340 42566
rect 168288 42502 168340 42508
rect 168196 42220 168248 42226
rect 168196 42162 168248 42168
rect 166908 41812 166960 41818
rect 166908 41754 166960 41760
rect 166356 41608 166408 41614
rect 166356 41550 166408 41556
rect 166920 3534 166948 41754
rect 165896 3528 165948 3534
rect 165896 3470 165948 3476
rect 166908 3528 166960 3534
rect 166908 3470 166960 3476
rect 164700 3460 164752 3466
rect 164700 3402 164752 3408
rect 165528 3460 165580 3466
rect 165528 3402 165580 3408
rect 164712 480 164740 3402
rect 165908 480 165936 3470
rect 167092 3120 167144 3126
rect 167092 3062 167144 3068
rect 167104 480 167132 3062
rect 168208 480 168236 42162
rect 168300 3126 168328 42502
rect 168392 42362 168420 44132
rect 168380 42356 168432 42362
rect 168380 42298 168432 42304
rect 169312 42022 169340 44132
rect 170324 42770 170352 44132
rect 170312 42764 170364 42770
rect 170312 42706 170364 42712
rect 169668 42696 169720 42702
rect 169668 42638 169720 42644
rect 169300 42016 169352 42022
rect 169300 41958 169352 41964
rect 168288 3120 168340 3126
rect 168288 3062 168340 3068
rect 169680 2854 169708 42638
rect 171336 42634 171364 44132
rect 171324 42628 171376 42634
rect 171324 42570 171376 42576
rect 171048 42356 171100 42362
rect 171048 42298 171100 42304
rect 171060 4146 171088 42298
rect 172256 41886 172284 44132
rect 172428 42628 172480 42634
rect 172428 42570 172480 42576
rect 172244 41880 172296 41886
rect 172244 41822 172296 41828
rect 172440 4146 172468 42570
rect 173268 42498 173296 44132
rect 173808 42764 173860 42770
rect 173808 42706 173860 42712
rect 173256 42492 173308 42498
rect 173256 42434 173308 42440
rect 170588 4140 170640 4146
rect 170588 4082 170640 4088
rect 171048 4140 171100 4146
rect 171048 4082 171100 4088
rect 171784 4140 171836 4146
rect 171784 4082 171836 4088
rect 172428 4140 172480 4146
rect 172428 4082 172480 4088
rect 169392 2848 169444 2854
rect 169392 2790 169444 2796
rect 169668 2848 169720 2854
rect 169668 2790 169720 2796
rect 169404 480 169432 2790
rect 170600 480 170628 4082
rect 171796 480 171824 4082
rect 173820 3534 173848 42706
rect 174280 42430 174308 44132
rect 174832 44118 175214 44146
rect 174268 42424 174320 42430
rect 174268 42366 174320 42372
rect 174832 41954 174860 44118
rect 175188 42492 175240 42498
rect 175188 42434 175240 42440
rect 174820 41948 174872 41954
rect 174820 41890 174872 41896
rect 175200 35902 175228 42434
rect 176212 41750 176240 44132
rect 176476 42424 176528 42430
rect 176476 42366 176528 42372
rect 176200 41744 176252 41750
rect 176200 41686 176252 41692
rect 175188 35896 175240 35902
rect 175188 35838 175240 35844
rect 175004 29028 175056 29034
rect 175004 28970 175056 28976
rect 175016 22166 175044 28970
rect 175004 22160 175056 22166
rect 175004 22102 175056 22108
rect 174820 22092 174872 22098
rect 174820 22034 174872 22040
rect 172980 3528 173032 3534
rect 172980 3470 173032 3476
rect 173808 3528 173860 3534
rect 173808 3470 173860 3476
rect 172992 480 173020 3470
rect 174832 3058 174860 22034
rect 176488 3330 176516 42366
rect 177132 42090 177160 44132
rect 178144 42158 178172 44132
rect 179156 42294 179184 44132
rect 179144 42288 179196 42294
rect 179144 42230 179196 42236
rect 178132 42152 178184 42158
rect 178132 42094 178184 42100
rect 179328 42152 179380 42158
rect 179328 42094 179380 42100
rect 177120 42084 177172 42090
rect 177120 42026 177172 42032
rect 177948 42084 178000 42090
rect 177948 42026 178000 42032
rect 176568 42016 176620 42022
rect 176568 41958 176620 41964
rect 175372 3324 175424 3330
rect 175372 3266 175424 3272
rect 176476 3324 176528 3330
rect 176476 3266 176528 3272
rect 174176 3052 174228 3058
rect 174176 2994 174228 3000
rect 174820 3052 174872 3058
rect 174820 2994 174872 3000
rect 174188 480 174216 2994
rect 175384 480 175412 3266
rect 176580 480 176608 41958
rect 177960 3482 177988 42026
rect 179340 3482 179368 42094
rect 180076 41818 180104 44132
rect 181088 42566 181116 44132
rect 181076 42560 181128 42566
rect 181076 42502 181128 42508
rect 180708 42288 180760 42294
rect 180708 42230 180760 42236
rect 180064 41812 180116 41818
rect 180064 41754 180116 41760
rect 180720 3534 180748 42230
rect 182100 42226 182128 44132
rect 183020 42702 183048 44132
rect 183008 42696 183060 42702
rect 183008 42638 183060 42644
rect 183468 42696 183520 42702
rect 183468 42638 183520 42644
rect 182180 42560 182232 42566
rect 182180 42502 182232 42508
rect 182088 42220 182140 42226
rect 182088 42162 182140 42168
rect 182192 42106 182220 42502
rect 182100 42078 182220 42106
rect 177776 3454 177988 3482
rect 178972 3454 179368 3482
rect 180156 3528 180208 3534
rect 180156 3470 180208 3476
rect 180708 3528 180760 3534
rect 180708 3470 180760 3476
rect 177776 480 177804 3454
rect 178972 480 179000 3454
rect 180168 480 180196 3470
rect 182100 3126 182128 42078
rect 183480 3534 183508 42638
rect 184032 42362 184060 44132
rect 185044 42634 185072 44132
rect 185964 42770 185992 44132
rect 185952 42764 186004 42770
rect 185952 42706 186004 42712
rect 185032 42628 185084 42634
rect 185032 42570 185084 42576
rect 186228 42628 186280 42634
rect 186228 42570 186280 42576
rect 184020 42356 184072 42362
rect 184020 42298 184072 42304
rect 184756 42220 184808 42226
rect 184756 42162 184808 42168
rect 183744 3596 183796 3602
rect 183744 3538 183796 3544
rect 182548 3528 182600 3534
rect 182548 3470 182600 3476
rect 183468 3528 183520 3534
rect 183468 3470 183520 3476
rect 181352 3120 181404 3126
rect 181352 3062 181404 3068
rect 182088 3120 182140 3126
rect 182088 3062 182140 3068
rect 181364 480 181392 3062
rect 182560 480 182588 3470
rect 183756 480 183784 3538
rect 184768 3482 184796 42162
rect 184848 41948 184900 41954
rect 184848 41890 184900 41896
rect 184860 3602 184888 41890
rect 184848 3596 184900 3602
rect 184848 3538 184900 3544
rect 186240 3482 186268 42570
rect 186976 42498 187004 44132
rect 186964 42492 187016 42498
rect 186964 42434 187016 42440
rect 187608 42492 187660 42498
rect 187608 42434 187660 42440
rect 187620 3482 187648 42434
rect 187988 42430 188016 44132
rect 187976 42424 188028 42430
rect 187976 42366 188028 42372
rect 188908 42022 188936 44132
rect 188988 42356 189040 42362
rect 188988 42298 189040 42304
rect 188896 42016 188948 42022
rect 188896 41958 188948 41964
rect 189000 3534 189028 42298
rect 189920 42090 189948 44132
rect 190368 42764 190420 42770
rect 190368 42706 190420 42712
rect 189908 42084 189960 42090
rect 189908 42026 189960 42032
rect 190380 3534 190408 42706
rect 190932 42158 190960 44132
rect 191748 42424 191800 42430
rect 191748 42366 191800 42372
rect 190920 42152 190972 42158
rect 190920 42094 190972 42100
rect 184768 3454 184888 3482
rect 184860 480 184888 3454
rect 186056 3454 186268 3482
rect 187252 3454 187648 3482
rect 188436 3528 188488 3534
rect 188436 3470 188488 3476
rect 188988 3528 189040 3534
rect 188988 3470 189040 3476
rect 189632 3528 189684 3534
rect 189632 3470 189684 3476
rect 190368 3528 190420 3534
rect 190368 3470 190420 3476
rect 186056 480 186084 3454
rect 187252 480 187280 3454
rect 188448 480 188476 3470
rect 189644 480 189672 3470
rect 191760 3058 191788 42366
rect 191852 42294 191880 44132
rect 192864 42566 192892 44132
rect 193784 42702 193812 44132
rect 193772 42696 193824 42702
rect 193772 42638 193824 42644
rect 192852 42560 192904 42566
rect 192852 42502 192904 42508
rect 191840 42288 191892 42294
rect 191840 42230 191892 42236
rect 193128 42152 193180 42158
rect 193128 42094 193180 42100
rect 193140 3534 193168 42094
rect 194416 42084 194468 42090
rect 194416 42026 194468 42032
rect 192024 3528 192076 3534
rect 192024 3470 192076 3476
rect 193128 3528 193180 3534
rect 193128 3470 193180 3476
rect 193220 3528 193272 3534
rect 193220 3470 193272 3476
rect 190828 3052 190880 3058
rect 190828 2994 190880 3000
rect 191748 3052 191800 3058
rect 191748 2994 191800 3000
rect 190840 480 190868 2994
rect 192036 480 192064 3470
rect 193232 480 193260 3470
rect 194428 480 194456 42026
rect 194796 41954 194824 44132
rect 195808 42226 195836 44132
rect 196728 42634 196756 44132
rect 196716 42628 196768 42634
rect 196716 42570 196768 42576
rect 197268 42628 197320 42634
rect 197268 42570 197320 42576
rect 195796 42220 195848 42226
rect 195796 42162 195848 42168
rect 195888 42220 195940 42226
rect 195888 42162 195940 42168
rect 194784 41948 194836 41954
rect 194784 41890 194836 41896
rect 194508 41472 194560 41478
rect 194508 41414 194560 41420
rect 194520 3534 194548 41414
rect 194508 3528 194560 3534
rect 195900 3482 195928 42162
rect 197280 3534 197308 42570
rect 197740 42498 197768 44132
rect 197728 42492 197780 42498
rect 197728 42434 197780 42440
rect 198648 42492 198700 42498
rect 198648 42434 198700 42440
rect 198660 3534 198688 42434
rect 198752 42362 198780 44132
rect 199672 42770 199700 44132
rect 199660 42764 199712 42770
rect 199660 42706 199712 42712
rect 200684 42430 200712 44132
rect 200672 42424 200724 42430
rect 200672 42366 200724 42372
rect 198740 42356 198792 42362
rect 198740 42298 198792 42304
rect 200028 42356 200080 42362
rect 200028 42298 200080 42304
rect 200040 3534 200068 42298
rect 201696 42158 201724 44132
rect 201684 42152 201736 42158
rect 201684 42094 201736 42100
rect 201408 41676 201460 41682
rect 201408 41618 201460 41624
rect 201420 3534 201448 41618
rect 202616 41478 202644 44132
rect 202788 42152 202840 42158
rect 202788 42094 202840 42100
rect 202696 41608 202748 41614
rect 202696 41550 202748 41556
rect 202604 41472 202656 41478
rect 202604 41414 202656 41420
rect 202708 3602 202736 41550
rect 201500 3596 201552 3602
rect 201500 3538 201552 3544
rect 202696 3596 202748 3602
rect 202696 3538 202748 3544
rect 194508 3470 194560 3476
rect 195624 3454 195928 3482
rect 196808 3528 196860 3534
rect 196808 3470 196860 3476
rect 197268 3528 197320 3534
rect 197268 3470 197320 3476
rect 198004 3528 198056 3534
rect 198004 3470 198056 3476
rect 198648 3528 198700 3534
rect 198648 3470 198700 3476
rect 199200 3528 199252 3534
rect 199200 3470 199252 3476
rect 200028 3528 200080 3534
rect 200028 3470 200080 3476
rect 200396 3528 200448 3534
rect 200396 3470 200448 3476
rect 201408 3528 201460 3534
rect 201408 3470 201460 3476
rect 195624 480 195652 3454
rect 196820 480 196848 3470
rect 198016 480 198044 3470
rect 199212 480 199240 3470
rect 200408 480 200436 3470
rect 201512 480 201540 3538
rect 202800 3482 202828 42094
rect 203628 42090 203656 44132
rect 204640 42226 204668 44132
rect 205560 42634 205588 44132
rect 205548 42628 205600 42634
rect 205548 42570 205600 42576
rect 206572 42498 206600 44132
rect 206560 42492 206612 42498
rect 206560 42434 206612 42440
rect 207584 42362 207612 44132
rect 207572 42356 207624 42362
rect 207572 42298 207624 42304
rect 208308 42356 208360 42362
rect 208308 42298 208360 42304
rect 204628 42220 204680 42226
rect 204628 42162 204680 42168
rect 206928 42220 206980 42226
rect 206928 42162 206980 42168
rect 203616 42084 203668 42090
rect 203616 42026 203668 42032
rect 204168 41540 204220 41546
rect 204168 41482 204220 41488
rect 204180 3482 204208 41482
rect 205548 41472 205600 41478
rect 205548 41414 205600 41420
rect 205560 3534 205588 41414
rect 202708 3454 202828 3482
rect 203904 3454 204208 3482
rect 205088 3528 205140 3534
rect 205088 3470 205140 3476
rect 205548 3528 205600 3534
rect 205548 3470 205600 3476
rect 202708 480 202736 3454
rect 203904 480 203932 3454
rect 205100 480 205128 3470
rect 206940 3058 206968 42162
rect 208320 3534 208348 42298
rect 208504 41682 208532 44132
rect 208492 41676 208544 41682
rect 208492 41618 208544 41624
rect 209516 41614 209544 44132
rect 209688 42288 209740 42294
rect 209688 42230 209740 42236
rect 209504 41608 209556 41614
rect 209504 41550 209556 41556
rect 209700 3534 209728 42230
rect 210436 42158 210464 44132
rect 210424 42152 210476 42158
rect 210424 42094 210476 42100
rect 211068 41744 211120 41750
rect 211068 41686 211120 41692
rect 210976 41608 211028 41614
rect 210976 41550 211028 41556
rect 210988 3534 211016 41550
rect 207480 3528 207532 3534
rect 207480 3470 207532 3476
rect 208308 3528 208360 3534
rect 208308 3470 208360 3476
rect 208676 3528 208728 3534
rect 208676 3470 208728 3476
rect 209688 3528 209740 3534
rect 209688 3470 209740 3476
rect 209872 3528 209924 3534
rect 209872 3470 209924 3476
rect 210976 3528 211028 3534
rect 210976 3470 211028 3476
rect 206284 3052 206336 3058
rect 206284 2994 206336 3000
rect 206928 3052 206980 3058
rect 206928 2994 206980 3000
rect 206296 480 206324 2994
rect 207492 480 207520 3470
rect 208688 480 208716 3470
rect 209884 480 209912 3470
rect 211080 480 211108 41686
rect 211448 41546 211476 44132
rect 211436 41540 211488 41546
rect 211436 41482 211488 41488
rect 212460 41478 212488 44132
rect 213380 42226 213408 44132
rect 214392 42362 214420 44132
rect 214380 42356 214432 42362
rect 214380 42298 214432 42304
rect 215404 42294 215432 44132
rect 215392 42288 215444 42294
rect 215392 42230 215444 42236
rect 213368 42220 213420 42226
rect 213368 42162 213420 42168
rect 213828 42220 213880 42226
rect 213828 42162 213880 42168
rect 212540 41676 212592 41682
rect 212540 41618 212592 41624
rect 212448 41472 212500 41478
rect 212448 41414 212500 41420
rect 212552 41290 212580 41618
rect 212460 41262 212580 41290
rect 212460 3482 212488 41262
rect 213840 3482 213868 42162
rect 216324 41614 216352 44132
rect 217336 41750 217364 44132
rect 217968 42152 218020 42158
rect 217968 42094 218020 42100
rect 217324 41744 217376 41750
rect 217324 41686 217376 41692
rect 216312 41608 216364 41614
rect 216312 41550 216364 41556
rect 215208 41540 215260 41546
rect 215208 41482 215260 41488
rect 215220 3534 215248 41482
rect 216588 41472 216640 41478
rect 216588 41414 216640 41420
rect 216600 3534 216628 41414
rect 217980 3534 218008 42094
rect 218348 41682 218376 44132
rect 219268 42226 219296 44132
rect 219348 42424 219400 42430
rect 219348 42366 219400 42372
rect 219256 42220 219308 42226
rect 219256 42162 219308 42168
rect 219256 42084 219308 42090
rect 219256 42026 219308 42032
rect 218336 41676 218388 41682
rect 218336 41618 218388 41624
rect 212276 3454 212488 3482
rect 213472 3454 213868 3482
rect 214656 3528 214708 3534
rect 214656 3470 214708 3476
rect 215208 3528 215260 3534
rect 215208 3470 215260 3476
rect 215852 3528 215904 3534
rect 215852 3470 215904 3476
rect 216588 3528 216640 3534
rect 216588 3470 216640 3476
rect 217048 3528 217100 3534
rect 217048 3470 217100 3476
rect 217968 3528 218020 3534
rect 217968 3470 218020 3476
rect 212276 480 212304 3454
rect 213472 480 213500 3454
rect 214668 480 214696 3470
rect 215864 480 215892 3470
rect 217060 480 217088 3470
rect 218152 3052 218204 3058
rect 218152 2994 218204 3000
rect 218164 480 218192 2994
rect 219268 1578 219296 42026
rect 219360 3058 219388 42366
rect 220280 41546 220308 44132
rect 220728 41676 220780 41682
rect 220728 41618 220780 41624
rect 220268 41540 220320 41546
rect 220268 41482 220320 41488
rect 220740 3482 220768 41618
rect 221292 41478 221320 44132
rect 222212 42158 222240 44132
rect 223224 42430 223252 44132
rect 223212 42424 223264 42430
rect 223212 42366 223264 42372
rect 222200 42152 222252 42158
rect 222200 42094 222252 42100
rect 224236 42090 224264 44132
rect 224224 42084 224276 42090
rect 224224 42026 224276 42032
rect 225156 41682 225184 44132
rect 225144 41676 225196 41682
rect 225144 41618 225196 41624
rect 224868 41608 224920 41614
rect 224868 41550 224920 41556
rect 222108 41540 222160 41546
rect 222108 41482 222160 41488
rect 221280 41472 221332 41478
rect 221280 41414 221332 41420
rect 222120 3482 222148 41482
rect 223488 41472 223540 41478
rect 223488 41414 223540 41420
rect 223500 3534 223528 41414
rect 224880 3534 224908 41550
rect 226168 41546 226196 44132
rect 226156 41540 226208 41546
rect 226156 41482 226208 41488
rect 226248 41540 226300 41546
rect 226248 41482 226300 41488
rect 226260 3534 226288 41482
rect 227088 41478 227116 44132
rect 228100 41614 228128 44132
rect 229008 42084 229060 42090
rect 229008 42026 229060 42032
rect 228088 41608 228140 41614
rect 228088 41550 228140 41556
rect 227076 41472 227128 41478
rect 227076 41414 227128 41420
rect 227628 41472 227680 41478
rect 227628 41414 227680 41420
rect 220556 3454 220768 3482
rect 221752 3454 222148 3482
rect 222936 3528 222988 3534
rect 222936 3470 222988 3476
rect 223488 3528 223540 3534
rect 223488 3470 223540 3476
rect 224132 3528 224184 3534
rect 224132 3470 224184 3476
rect 224868 3528 224920 3534
rect 224868 3470 224920 3476
rect 225328 3528 225380 3534
rect 225328 3470 225380 3476
rect 226248 3528 226300 3534
rect 226248 3470 226300 3476
rect 219348 3052 219400 3058
rect 219348 2994 219400 3000
rect 219268 1550 219388 1578
rect 219360 480 219388 1550
rect 220556 480 220584 3454
rect 221752 480 221780 3454
rect 222948 480 222976 3470
rect 224144 480 224172 3470
rect 225340 480 225368 3470
rect 227640 3330 227668 41414
rect 227720 3732 227772 3738
rect 227720 3674 227772 3680
rect 226524 3324 226576 3330
rect 226524 3266 226576 3272
rect 227628 3324 227680 3330
rect 227628 3266 227680 3272
rect 226536 480 226564 3266
rect 227732 480 227760 3674
rect 229020 3482 229048 42026
rect 229112 41546 229140 44132
rect 229100 41540 229152 41546
rect 229100 41482 229152 41488
rect 230032 41478 230060 44132
rect 230584 44118 231058 44146
rect 230388 41540 230440 41546
rect 230388 41482 230440 41488
rect 230020 41472 230072 41478
rect 230020 41414 230072 41420
rect 230400 3482 230428 41482
rect 230584 3738 230612 44118
rect 232056 42090 232084 44132
rect 232044 42084 232096 42090
rect 232044 42026 232096 42032
rect 232976 41546 233004 44132
rect 232964 41540 233016 41546
rect 232964 41482 233016 41488
rect 233148 41540 233200 41546
rect 233148 41482 233200 41488
rect 231768 41472 231820 41478
rect 231768 41414 231820 41420
rect 230572 3732 230624 3738
rect 230572 3674 230624 3680
rect 231780 3534 231808 41414
rect 233160 3534 233188 41482
rect 233988 41478 234016 44132
rect 235000 41546 235028 44132
rect 234988 41540 235040 41546
rect 234988 41482 235040 41488
rect 235920 41478 235948 44132
rect 236196 44118 236946 44146
rect 237392 44118 237958 44146
rect 233976 41472 234028 41478
rect 233976 41414 234028 41420
rect 234528 41472 234580 41478
rect 234528 41414 234580 41420
rect 235908 41472 235960 41478
rect 235908 41414 235960 41420
rect 234540 3534 234568 41414
rect 236000 3596 236052 3602
rect 236000 3538 236052 3544
rect 228928 3454 229048 3482
rect 230124 3454 230428 3482
rect 231308 3528 231360 3534
rect 231308 3470 231360 3476
rect 231768 3528 231820 3534
rect 231768 3470 231820 3476
rect 232504 3528 232556 3534
rect 232504 3470 232556 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 233700 3528 233752 3534
rect 233700 3470 233752 3476
rect 234528 3528 234580 3534
rect 234528 3470 234580 3476
rect 234804 3528 234856 3534
rect 234804 3470 234856 3476
rect 228928 480 228956 3454
rect 230124 480 230152 3454
rect 231320 480 231348 3470
rect 232516 480 232544 3470
rect 233712 480 233740 3470
rect 234816 480 234844 3470
rect 236012 480 236040 3538
rect 236196 3534 236224 44118
rect 237288 42764 237340 42770
rect 237288 42706 237340 42712
rect 236184 3528 236236 3534
rect 237300 3482 237328 42706
rect 237392 3602 237420 44118
rect 238864 42770 238892 44132
rect 239600 44118 239890 44146
rect 238852 42764 238904 42770
rect 238852 42706 238904 42712
rect 239600 40050 239628 44118
rect 240888 42770 240916 44132
rect 241624 44118 241822 44146
rect 242544 44118 242834 44146
rect 242912 44118 243754 44146
rect 244292 44118 244766 44146
rect 241624 42786 241652 44118
rect 240048 42764 240100 42770
rect 240048 42706 240100 42712
rect 240876 42764 240928 42770
rect 240876 42706 240928 42712
rect 241440 42758 241652 42786
rect 238852 40044 238904 40050
rect 238852 39986 238904 39992
rect 239588 40044 239640 40050
rect 239588 39986 239640 39992
rect 238864 4146 238892 39986
rect 238392 4140 238444 4146
rect 238392 4082 238444 4088
rect 238852 4140 238904 4146
rect 238852 4082 238904 4088
rect 237380 3596 237432 3602
rect 237380 3538 237432 3544
rect 236184 3470 236236 3476
rect 237208 3454 237328 3482
rect 237208 480 237236 3454
rect 238404 480 238432 4082
rect 240060 3534 240088 42706
rect 241440 4146 241468 42758
rect 242544 35970 242572 44118
rect 241612 35964 241664 35970
rect 241612 35906 241664 35912
rect 242532 35964 242584 35970
rect 242532 35906 242584 35912
rect 241624 4842 241652 35906
rect 242912 4842 242940 44118
rect 244292 38622 244320 44118
rect 245764 42786 245792 44132
rect 245580 42758 245792 42786
rect 244280 38616 244332 38622
rect 244280 38558 244332 38564
rect 244372 38616 244424 38622
rect 244372 38558 244424 38564
rect 244384 37262 244412 38558
rect 244372 37256 244424 37262
rect 244372 37198 244424 37204
rect 244280 27668 244332 27674
rect 244280 27610 244332 27616
rect 244292 22778 244320 27610
rect 244280 22772 244332 22778
rect 244280 22714 244332 22720
rect 244372 9716 244424 9722
rect 244372 9658 244424 9664
rect 241624 4814 242020 4842
rect 242912 4814 243216 4842
rect 240784 4140 240836 4146
rect 240784 4082 240836 4088
rect 241428 4140 241480 4146
rect 241428 4082 241480 4088
rect 239588 3528 239640 3534
rect 239588 3470 239640 3476
rect 240048 3528 240100 3534
rect 240048 3470 240100 3476
rect 239600 480 239628 3470
rect 240796 480 240824 4082
rect 241992 480 242020 4814
rect 243188 480 243216 4814
rect 244384 480 244412 9658
rect 245580 480 245608 42758
rect 246132 41426 246160 44254
rect 246040 41398 246160 41426
rect 247052 44118 247710 44146
rect 248524 44118 248722 44146
rect 249642 44118 249748 44146
rect 250654 44118 251128 44146
rect 246040 38622 246068 41398
rect 246028 38616 246080 38622
rect 246028 38558 246080 38564
rect 245936 29028 245988 29034
rect 245936 28970 245988 28976
rect 245948 22114 245976 28970
rect 245856 22098 245976 22114
rect 245844 22092 245976 22098
rect 245896 22086 245976 22092
rect 246028 22092 246080 22098
rect 245844 22034 245896 22040
rect 246028 22034 246080 22040
rect 246040 19310 246068 22034
rect 246028 19304 246080 19310
rect 246028 19246 246080 19252
rect 246028 9716 246080 9722
rect 246028 9658 246080 9664
rect 246040 4146 246068 9658
rect 247052 4146 247080 44118
rect 248524 4146 248552 44118
rect 249720 4146 249748 44118
rect 246028 4140 246080 4146
rect 246028 4082 246080 4088
rect 246764 4140 246816 4146
rect 246764 4082 246816 4088
rect 247040 4140 247092 4146
rect 247040 4082 247092 4088
rect 247960 4140 248012 4146
rect 247960 4082 248012 4088
rect 248512 4140 248564 4146
rect 248512 4082 248564 4088
rect 249156 4140 249208 4146
rect 249156 4082 249208 4088
rect 249708 4140 249760 4146
rect 249708 4082 249760 4088
rect 250352 4140 250404 4146
rect 250352 4082 250404 4088
rect 246776 480 246804 4082
rect 247972 480 248000 4082
rect 249168 480 249196 4082
rect 250364 480 250392 4082
rect 251100 4026 251128 44118
rect 251652 42770 251680 44132
rect 251640 42764 251692 42770
rect 251640 42706 251692 42712
rect 252468 42764 252520 42770
rect 252468 42706 252520 42712
rect 252480 12442 252508 42706
rect 252284 12436 252336 12442
rect 252284 12378 252336 12384
rect 252468 12436 252520 12442
rect 252468 12378 252520 12384
rect 252296 4078 252324 12378
rect 252572 4146 252600 44132
rect 253598 44118 253888 44146
rect 254610 44118 255268 44146
rect 253860 41426 253888 44118
rect 253860 41398 254072 41426
rect 252560 4140 252612 4146
rect 252560 4082 252612 4088
rect 253848 4140 253900 4146
rect 253848 4082 253900 4088
rect 252284 4072 252336 4078
rect 251100 3998 251496 4026
rect 252284 4014 252336 4020
rect 252652 4072 252704 4078
rect 252652 4014 252704 4020
rect 251468 480 251496 3998
rect 252664 480 252692 4014
rect 253860 480 253888 4082
rect 254044 610 254072 41398
rect 255240 3534 255268 44118
rect 255516 41478 255544 44132
rect 256542 44118 256648 44146
rect 255504 41472 255556 41478
rect 255504 41414 255556 41420
rect 255228 3528 255280 3534
rect 255228 3470 255280 3476
rect 256240 3528 256292 3534
rect 256240 3470 256292 3476
rect 254032 604 254084 610
rect 254032 546 254084 552
rect 255044 604 255096 610
rect 255044 546 255096 552
rect 255056 480 255084 546
rect 256252 480 256280 3470
rect 256620 3330 256648 44118
rect 257540 41546 257568 44132
rect 257528 41540 257580 41546
rect 257528 41482 257580 41488
rect 258460 41478 258488 44132
rect 258724 41540 258776 41546
rect 258724 41482 258776 41488
rect 256700 41472 256752 41478
rect 256700 41414 256752 41420
rect 258448 41472 258500 41478
rect 258448 41414 258500 41420
rect 256608 3324 256660 3330
rect 256608 3266 256660 3272
rect 256712 610 256740 41414
rect 258736 3534 258764 41482
rect 259472 41478 259500 44132
rect 260406 44118 260788 44146
rect 261418 44118 262168 44146
rect 259368 41472 259420 41478
rect 259368 41414 259420 41420
rect 259460 41472 259512 41478
rect 259460 41414 259512 41420
rect 258724 3528 258776 3534
rect 258724 3470 258776 3476
rect 259380 3466 259408 41414
rect 259828 3528 259880 3534
rect 259828 3470 259880 3476
rect 259368 3460 259420 3466
rect 259368 3402 259420 3408
rect 258632 3324 258684 3330
rect 258632 3266 258684 3272
rect 256700 604 256752 610
rect 256700 546 256752 552
rect 257436 604 257488 610
rect 257436 546 257488 552
rect 257448 480 257476 546
rect 258644 480 258672 3266
rect 259840 480 259868 3470
rect 260760 3398 260788 44118
rect 261484 41472 261536 41478
rect 261484 41414 261536 41420
rect 261496 3534 261524 41414
rect 261484 3528 261536 3534
rect 261484 3470 261536 3476
rect 261024 3460 261076 3466
rect 261024 3402 261076 3408
rect 260748 3392 260800 3398
rect 260748 3334 260800 3340
rect 261036 480 261064 3402
rect 262140 3126 262168 44118
rect 262416 41478 262444 44132
rect 263350 44118 263548 44146
rect 262404 41472 262456 41478
rect 262404 41414 262456 41420
rect 263416 41472 263468 41478
rect 263416 41414 263468 41420
rect 263428 3534 263456 41414
rect 263520 3602 263548 44118
rect 264348 41546 264376 44132
rect 264336 41540 264388 41546
rect 264336 41482 264388 41488
rect 265360 41478 265388 44132
rect 265348 41472 265400 41478
rect 265348 41414 265400 41420
rect 266176 41472 266228 41478
rect 266176 41414 266228 41420
rect 263508 3596 263560 3602
rect 263508 3538 263560 3544
rect 262220 3528 262272 3534
rect 262220 3470 262272 3476
rect 263416 3528 263468 3534
rect 263416 3470 263468 3476
rect 265808 3528 265860 3534
rect 265808 3470 265860 3476
rect 262128 3120 262180 3126
rect 262128 3062 262180 3068
rect 262232 480 262260 3470
rect 263416 3392 263468 3398
rect 263416 3334 263468 3340
rect 263428 480 263456 3334
rect 264612 3120 264664 3126
rect 264612 3062 264664 3068
rect 264624 480 264652 3062
rect 265820 480 265848 3470
rect 266188 3466 266216 41414
rect 266280 3534 266308 44132
rect 267306 44118 267688 44146
rect 267004 41540 267056 41546
rect 267004 41482 267056 41488
rect 267016 4146 267044 41482
rect 267004 4140 267056 4146
rect 267004 4082 267056 4088
rect 267660 3738 267688 44118
rect 268304 41478 268332 44132
rect 269224 41478 269252 44132
rect 270250 44118 270356 44146
rect 268292 41472 268344 41478
rect 268292 41414 268344 41420
rect 269028 41472 269080 41478
rect 269028 41414 269080 41420
rect 269212 41472 269264 41478
rect 269212 41414 269264 41420
rect 268108 4140 268160 4146
rect 268108 4082 268160 4088
rect 267648 3732 267700 3738
rect 267648 3674 267700 3680
rect 267004 3596 267056 3602
rect 267004 3538 267056 3544
rect 266268 3528 266320 3534
rect 266268 3470 266320 3476
rect 266176 3460 266228 3466
rect 266176 3402 266228 3408
rect 267016 480 267044 3538
rect 268120 480 268148 4082
rect 269040 3194 269068 41414
rect 270328 3466 270356 44118
rect 271248 41546 271276 44132
rect 271236 41540 271288 41546
rect 271236 41482 271288 41488
rect 272168 41478 272196 44132
rect 272524 41540 272576 41546
rect 272524 41482 272576 41488
rect 270408 41472 270460 41478
rect 270408 41414 270460 41420
rect 272156 41472 272208 41478
rect 272156 41414 272208 41420
rect 270420 3602 270448 41414
rect 271696 3732 271748 3738
rect 271696 3674 271748 3680
rect 270408 3596 270460 3602
rect 270408 3538 270460 3544
rect 270500 3528 270552 3534
rect 270500 3470 270552 3476
rect 269304 3460 269356 3466
rect 269304 3402 269356 3408
rect 270316 3460 270368 3466
rect 270316 3402 270368 3408
rect 269028 3188 269080 3194
rect 269028 3130 269080 3136
rect 269316 480 269344 3402
rect 270512 480 270540 3470
rect 271708 480 271736 3674
rect 272536 3330 272564 41482
rect 273076 41472 273128 41478
rect 273076 41414 273128 41420
rect 272524 3324 272576 3330
rect 272524 3266 272576 3272
rect 272892 3188 272944 3194
rect 272892 3130 272944 3136
rect 272904 480 272932 3130
rect 273088 3126 273116 41414
rect 273180 3874 273208 44132
rect 274206 44118 274588 44146
rect 273168 3868 273220 3874
rect 273168 3810 273220 3816
rect 274088 3596 274140 3602
rect 274088 3538 274140 3544
rect 273076 3120 273128 3126
rect 273076 3062 273128 3068
rect 274100 480 274128 3538
rect 274560 2990 274588 44118
rect 275112 41478 275140 44132
rect 276124 41478 276152 44132
rect 277058 44118 277256 44146
rect 278070 44118 278728 44146
rect 275100 41472 275152 41478
rect 275100 41414 275152 41420
rect 275928 41472 275980 41478
rect 275928 41414 275980 41420
rect 276112 41472 276164 41478
rect 276112 41414 276164 41420
rect 275940 3670 275968 41414
rect 275928 3664 275980 3670
rect 275928 3606 275980 3612
rect 277228 3466 277256 44118
rect 277308 41472 277360 41478
rect 277308 41414 277360 41420
rect 277320 3806 277348 41414
rect 277308 3800 277360 3806
rect 277308 3742 277360 3748
rect 275284 3460 275336 3466
rect 275284 3402 275336 3408
rect 277216 3460 277268 3466
rect 277216 3402 277268 3408
rect 274548 2984 274600 2990
rect 274548 2926 274600 2932
rect 275296 480 275324 3402
rect 278700 3330 278728 44118
rect 279068 41478 279096 44132
rect 279056 41472 279108 41478
rect 279056 41414 279108 41420
rect 278872 3868 278924 3874
rect 278872 3810 278924 3816
rect 276480 3324 276532 3330
rect 276480 3266 276532 3272
rect 278688 3324 278740 3330
rect 278688 3266 278740 3272
rect 276492 480 276520 3266
rect 277676 3120 277728 3126
rect 277676 3062 277728 3068
rect 277688 480 277716 3062
rect 278884 480 278912 3810
rect 279988 3602 280016 44132
rect 281014 44118 281488 44146
rect 280068 41472 280120 41478
rect 280068 41414 280120 41420
rect 279976 3596 280028 3602
rect 279976 3538 280028 3544
rect 280080 3534 280108 41414
rect 281264 3664 281316 3670
rect 281264 3606 281316 3612
rect 280068 3528 280120 3534
rect 280068 3470 280120 3476
rect 280068 2984 280120 2990
rect 280068 2926 280120 2932
rect 280080 480 280108 2926
rect 281276 480 281304 3606
rect 281460 3398 281488 44118
rect 282012 41478 282040 44132
rect 282932 41478 282960 44132
rect 283958 44118 284248 44146
rect 284970 44118 285628 44146
rect 282000 41472 282052 41478
rect 282000 41414 282052 41420
rect 282828 41472 282880 41478
rect 282828 41414 282880 41420
rect 282920 41472 282972 41478
rect 282920 41414 282972 41420
rect 284116 41472 284168 41478
rect 284116 41414 284168 41420
rect 282460 3800 282512 3806
rect 282460 3742 282512 3748
rect 281448 3392 281500 3398
rect 281448 3334 281500 3340
rect 282472 480 282500 3742
rect 282840 3058 282868 41414
rect 284128 3670 284156 41414
rect 284220 3806 284248 44118
rect 285600 3874 285628 44118
rect 285876 41478 285904 44132
rect 286902 44118 287008 44146
rect 287914 44118 288388 44146
rect 285864 41472 285916 41478
rect 285864 41414 285916 41420
rect 286876 41472 286928 41478
rect 286876 41414 286928 41420
rect 285588 3868 285640 3874
rect 285588 3810 285640 3816
rect 284208 3800 284260 3806
rect 284208 3742 284260 3748
rect 284116 3664 284168 3670
rect 284116 3606 284168 3612
rect 286888 3602 286916 41414
rect 286876 3596 286928 3602
rect 286876 3538 286928 3544
rect 285956 3528 286008 3534
rect 285956 3470 286008 3476
rect 283656 3460 283708 3466
rect 283656 3402 283708 3408
rect 282828 3052 282880 3058
rect 282828 2994 282880 3000
rect 283668 480 283696 3402
rect 284760 3324 284812 3330
rect 284760 3266 284812 3272
rect 284772 480 284800 3266
rect 285968 480 285996 3470
rect 286980 3466 287008 44118
rect 288360 3534 288388 44118
rect 288820 41478 288848 44132
rect 289832 41478 289860 44132
rect 290858 44118 291056 44146
rect 291778 44118 292528 44146
rect 288808 41472 288860 41478
rect 288808 41414 288860 41420
rect 289728 41472 289780 41478
rect 289728 41414 289780 41420
rect 289820 41472 289872 41478
rect 289820 41414 289872 41420
rect 289740 4078 289768 41414
rect 289728 4072 289780 4078
rect 289728 4014 289780 4020
rect 291028 3670 291056 44118
rect 291108 41472 291160 41478
rect 291108 41414 291160 41420
rect 290740 3664 290792 3670
rect 290740 3606 290792 3612
rect 291016 3664 291068 3670
rect 291016 3606 291068 3612
rect 287152 3528 287204 3534
rect 287152 3470 287204 3476
rect 288348 3528 288400 3534
rect 288348 3470 288400 3476
rect 286968 3460 287020 3466
rect 286968 3402 287020 3408
rect 287164 480 287192 3470
rect 288348 3392 288400 3398
rect 288348 3334 288400 3340
rect 288360 480 288388 3334
rect 289544 3052 289596 3058
rect 289544 2994 289596 3000
rect 289556 480 289584 2994
rect 290752 480 290780 3606
rect 291120 2990 291148 41414
rect 292500 3806 292528 44118
rect 292776 41478 292804 44132
rect 293710 44118 293908 44146
rect 294722 44118 295288 44146
rect 292764 41472 292816 41478
rect 292764 41414 292816 41420
rect 293776 41472 293828 41478
rect 293776 41414 293828 41420
rect 293788 3874 293816 41414
rect 293880 3942 293908 44118
rect 295260 4010 295288 44118
rect 295720 41478 295748 44132
rect 295708 41472 295760 41478
rect 295708 41414 295760 41420
rect 296536 41472 296588 41478
rect 296536 41414 296588 41420
rect 295248 4004 295300 4010
rect 295248 3946 295300 3952
rect 293868 3936 293920 3942
rect 293868 3878 293920 3884
rect 293132 3868 293184 3874
rect 293132 3810 293184 3816
rect 293776 3868 293828 3874
rect 293776 3810 293828 3816
rect 291936 3800 291988 3806
rect 291936 3742 291988 3748
rect 292488 3800 292540 3806
rect 292488 3742 292540 3748
rect 291108 2984 291160 2990
rect 291108 2926 291160 2932
rect 291948 480 291976 3742
rect 293144 480 293172 3810
rect 294328 3596 294380 3602
rect 294328 3538 294380 3544
rect 294340 480 294368 3538
rect 295524 3460 295576 3466
rect 295524 3402 295576 3408
rect 295536 480 295564 3402
rect 296548 3398 296576 41414
rect 296640 3466 296668 44132
rect 297666 44118 298048 44146
rect 297916 4072 297968 4078
rect 297916 4014 297968 4020
rect 296720 3528 296772 3534
rect 296720 3470 296772 3476
rect 296628 3460 296680 3466
rect 296628 3402 296680 3408
rect 296536 3392 296588 3398
rect 296536 3334 296588 3340
rect 296732 480 296760 3470
rect 297928 480 297956 4014
rect 298020 3602 298048 44118
rect 298664 41478 298692 44132
rect 299584 41478 299612 44132
rect 300610 44118 300716 44146
rect 301622 44118 302188 44146
rect 298652 41472 298704 41478
rect 298652 41414 298704 41420
rect 299388 41472 299440 41478
rect 299388 41414 299440 41420
rect 299572 41472 299624 41478
rect 299572 41414 299624 41420
rect 298008 3596 298060 3602
rect 298008 3538 298060 3544
rect 299400 3534 299428 41414
rect 300688 3738 300716 44118
rect 300768 41472 300820 41478
rect 300768 41414 300820 41420
rect 300676 3732 300728 3738
rect 300676 3674 300728 3680
rect 300780 3670 300808 41414
rect 302160 3806 302188 44118
rect 302528 41478 302556 44132
rect 303448 44118 303554 44146
rect 304566 44118 304948 44146
rect 302516 41472 302568 41478
rect 302516 41414 302568 41420
rect 303448 3874 303476 44118
rect 303528 41472 303580 41478
rect 303528 41414 303580 41420
rect 303540 4146 303568 41414
rect 303528 4140 303580 4146
rect 303528 4082 303580 4088
rect 303804 3936 303856 3942
rect 303804 3878 303856 3884
rect 302608 3868 302660 3874
rect 302608 3810 302660 3816
rect 303436 3868 303488 3874
rect 303436 3810 303488 3816
rect 301412 3800 301464 3806
rect 301412 3742 301464 3748
rect 302148 3800 302200 3806
rect 302148 3742 302200 3748
rect 300308 3664 300360 3670
rect 300308 3606 300360 3612
rect 300768 3664 300820 3670
rect 300768 3606 300820 3612
rect 299388 3528 299440 3534
rect 299388 3470 299440 3476
rect 299112 2984 299164 2990
rect 299112 2926 299164 2932
rect 299124 480 299152 2926
rect 300320 480 300348 3606
rect 301424 480 301452 3742
rect 302620 480 302648 3810
rect 303816 480 303844 3878
rect 304920 3330 304948 44118
rect 305472 41478 305500 44132
rect 306484 41478 306512 44132
rect 307510 44118 307708 44146
rect 308430 44118 309088 44146
rect 305460 41472 305512 41478
rect 305460 41414 305512 41420
rect 306288 41472 306340 41478
rect 306288 41414 306340 41420
rect 306472 41472 306524 41478
rect 306472 41414 306524 41420
rect 307576 41472 307628 41478
rect 307576 41414 307628 41420
rect 305000 4004 305052 4010
rect 305000 3946 305052 3952
rect 304908 3324 304960 3330
rect 304908 3266 304960 3272
rect 305012 480 305040 3946
rect 306300 3398 306328 41414
rect 307588 4010 307616 41414
rect 307576 4004 307628 4010
rect 307576 3946 307628 3952
rect 307680 3466 307708 44118
rect 309060 3602 309088 44118
rect 309428 41478 309456 44132
rect 310362 44118 310468 44146
rect 311374 44118 311848 44146
rect 309416 41472 309468 41478
rect 309416 41414 309468 41420
rect 310336 41472 310388 41478
rect 310336 41414 310388 41420
rect 310348 4078 310376 41414
rect 310336 4072 310388 4078
rect 310336 4014 310388 4020
rect 308588 3596 308640 3602
rect 308588 3538 308640 3544
rect 309048 3596 309100 3602
rect 309048 3538 309100 3544
rect 307392 3460 307444 3466
rect 307392 3402 307444 3408
rect 307668 3460 307720 3466
rect 307668 3402 307720 3408
rect 306196 3392 306248 3398
rect 306196 3334 306248 3340
rect 306288 3392 306340 3398
rect 306288 3334 306340 3340
rect 306208 480 306236 3334
rect 307404 480 307432 3402
rect 308600 480 308628 3538
rect 310440 3534 310468 44118
rect 311820 3670 311848 44118
rect 312372 41478 312400 44132
rect 313292 41478 313320 44132
rect 314318 44118 314516 44146
rect 315330 44118 315988 44146
rect 312360 41472 312412 41478
rect 312360 41414 312412 41420
rect 313188 41472 313240 41478
rect 313188 41414 313240 41420
rect 313280 41472 313332 41478
rect 313280 41414 313332 41420
rect 313200 3942 313228 41414
rect 314384 4140 314436 4146
rect 314384 4082 314436 4088
rect 313188 3936 313240 3942
rect 313188 3878 313240 3884
rect 313372 3800 313424 3806
rect 313372 3742 313424 3748
rect 312176 3732 312228 3738
rect 312176 3674 312228 3680
rect 310980 3664 311032 3670
rect 310980 3606 311032 3612
rect 311808 3664 311860 3670
rect 311808 3606 311860 3612
rect 309784 3528 309836 3534
rect 309784 3470 309836 3476
rect 310428 3528 310480 3534
rect 310428 3470 310480 3476
rect 309796 480 309824 3470
rect 310992 480 311020 3606
rect 312188 480 312216 3674
rect 313384 480 313412 3742
rect 314396 3618 314424 4082
rect 314488 3806 314516 44118
rect 314568 41472 314620 41478
rect 314568 41414 314620 41420
rect 314580 4146 314608 41414
rect 314568 4140 314620 4146
rect 314568 4082 314620 4088
rect 315960 3874 315988 44118
rect 316236 41478 316264 44132
rect 317262 44118 317368 44146
rect 318274 44118 318748 44146
rect 316224 41472 316276 41478
rect 316224 41414 316276 41420
rect 317236 41472 317288 41478
rect 317236 41414 317288 41420
rect 315764 3868 315816 3874
rect 315764 3810 315816 3816
rect 315948 3868 316000 3874
rect 315948 3810 316000 3816
rect 314476 3800 314528 3806
rect 314476 3742 314528 3748
rect 314396 3590 314608 3618
rect 314580 480 314608 3590
rect 315776 480 315804 3810
rect 317248 3738 317276 41414
rect 317236 3732 317288 3738
rect 317236 3674 317288 3680
rect 317340 3330 317368 44118
rect 318064 3392 318116 3398
rect 318064 3334 318116 3340
rect 316960 3324 317012 3330
rect 316960 3266 317012 3272
rect 317328 3324 317380 3330
rect 317328 3266 317380 3272
rect 316972 480 317000 3266
rect 318076 480 318104 3334
rect 318720 3194 318748 44118
rect 319180 41478 319208 44132
rect 320192 41478 320220 44132
rect 321218 44118 321416 44146
rect 322138 44118 322888 44146
rect 319168 41472 319220 41478
rect 319168 41414 319220 41420
rect 320088 41472 320140 41478
rect 320088 41414 320140 41420
rect 320180 41472 320232 41478
rect 320180 41414 320232 41420
rect 319260 4004 319312 4010
rect 319260 3946 319312 3952
rect 318708 3188 318760 3194
rect 318708 3130 318760 3136
rect 319272 480 319300 3946
rect 320100 3126 320128 41414
rect 321388 3466 321416 44118
rect 321468 41472 321520 41478
rect 321468 41414 321520 41420
rect 320456 3460 320508 3466
rect 320456 3402 320508 3408
rect 321376 3460 321428 3466
rect 321376 3402 321428 3408
rect 320088 3120 320140 3126
rect 320088 3062 320140 3068
rect 320468 480 320496 3402
rect 321480 2922 321508 41414
rect 322756 4072 322808 4078
rect 322756 4014 322808 4020
rect 321652 3596 321704 3602
rect 321652 3538 321704 3544
rect 321468 2916 321520 2922
rect 321468 2858 321520 2864
rect 321664 480 321692 3538
rect 322768 3482 322796 4014
rect 322860 3602 322888 44118
rect 323136 41478 323164 44132
rect 323124 41472 323176 41478
rect 323124 41414 323176 41420
rect 322848 3596 322900 3602
rect 322848 3538 322900 3544
rect 324148 3534 324176 44132
rect 325082 44118 325648 44146
rect 324228 41472 324280 41478
rect 324228 41414 324280 41420
rect 324044 3528 324096 3534
rect 322768 3454 322888 3482
rect 324044 3470 324096 3476
rect 324136 3528 324188 3534
rect 324136 3470 324188 3476
rect 322860 480 322888 3454
rect 324056 480 324084 3470
rect 324240 3262 324268 41414
rect 325620 4078 325648 44118
rect 326080 41478 326108 44132
rect 326068 41472 326120 41478
rect 326068 41414 326120 41420
rect 326896 41472 326948 41478
rect 326896 41414 326948 41420
rect 325608 4072 325660 4078
rect 325608 4014 325660 4020
rect 326436 3936 326488 3942
rect 326436 3878 326488 3884
rect 325240 3664 325292 3670
rect 325240 3606 325292 3612
rect 324228 3256 324280 3262
rect 324228 3198 324280 3204
rect 325252 480 325280 3606
rect 326448 480 326476 3878
rect 326908 3670 326936 41414
rect 327000 4010 327028 44132
rect 328026 44118 328408 44146
rect 328380 4146 328408 44118
rect 329024 41478 329052 44132
rect 329944 41478 329972 44132
rect 330970 44118 331168 44146
rect 331982 44118 332548 44146
rect 329012 41472 329064 41478
rect 329012 41414 329064 41420
rect 329748 41472 329800 41478
rect 329748 41414 329800 41420
rect 329932 41472 329984 41478
rect 329932 41414 329984 41420
rect 331036 41472 331088 41478
rect 331036 41414 331088 41420
rect 327632 4140 327684 4146
rect 327632 4082 327684 4088
rect 328368 4140 328420 4146
rect 328368 4082 328420 4088
rect 326988 4004 327040 4010
rect 326988 3946 327040 3952
rect 326896 3664 326948 3670
rect 326896 3606 326948 3612
rect 327644 480 327672 4082
rect 328828 3800 328880 3806
rect 328828 3742 328880 3748
rect 328840 480 328868 3742
rect 329760 3398 329788 41414
rect 331048 3942 331076 41414
rect 331036 3936 331088 3942
rect 331036 3878 331088 3884
rect 330024 3868 330076 3874
rect 330024 3810 330076 3816
rect 329748 3392 329800 3398
rect 329748 3334 329800 3340
rect 330036 480 330064 3810
rect 331140 2990 331168 44118
rect 331220 3732 331272 3738
rect 331220 3674 331272 3680
rect 331128 2984 331180 2990
rect 331128 2926 331180 2932
rect 331232 480 331260 3674
rect 332416 3324 332468 3330
rect 332416 3266 332468 3272
rect 332428 480 332456 3266
rect 332520 3058 332548 44118
rect 332888 41478 332916 44132
rect 332876 41472 332928 41478
rect 332876 41414 332928 41420
rect 333796 41472 333848 41478
rect 333796 41414 333848 41420
rect 333808 3330 333836 41414
rect 333900 3738 333928 44132
rect 334926 44118 335308 44146
rect 335280 3806 335308 44118
rect 335832 41478 335860 44132
rect 336844 41478 336872 44132
rect 337870 44118 337976 44146
rect 338790 44118 339448 44146
rect 335820 41472 335872 41478
rect 335820 41414 335872 41420
rect 336648 41472 336700 41478
rect 336648 41414 336700 41420
rect 336832 41472 336884 41478
rect 336832 41414 336884 41420
rect 336660 3874 336688 41414
rect 336648 3868 336700 3874
rect 336648 3810 336700 3816
rect 335268 3800 335320 3806
rect 335268 3742 335320 3748
rect 333888 3732 333940 3738
rect 333888 3674 333940 3680
rect 337948 3466 337976 44118
rect 338028 41472 338080 41478
rect 338028 41414 338080 41420
rect 337108 3460 337160 3466
rect 337108 3402 337160 3408
rect 337936 3460 337988 3466
rect 337936 3402 337988 3408
rect 333796 3324 333848 3330
rect 333796 3266 333848 3272
rect 333612 3188 333664 3194
rect 333612 3130 333664 3136
rect 332508 3052 332560 3058
rect 332508 2994 332560 3000
rect 333624 480 333652 3130
rect 334716 3120 334768 3126
rect 334716 3062 334768 3068
rect 334728 480 334756 3062
rect 335912 2916 335964 2922
rect 335912 2858 335964 2864
rect 335924 480 335952 2858
rect 337120 480 337148 3402
rect 338040 3194 338068 41414
rect 339420 3602 339448 44118
rect 339788 41478 339816 44132
rect 340708 44118 340814 44146
rect 341734 44118 342208 44146
rect 339776 41472 339828 41478
rect 339776 41414 339828 41420
rect 340512 5364 340564 5370
rect 340512 5306 340564 5312
rect 338304 3596 338356 3602
rect 338304 3538 338356 3544
rect 339408 3596 339460 3602
rect 339408 3538 339460 3544
rect 338028 3188 338080 3194
rect 338028 3130 338080 3136
rect 338316 480 338344 3538
rect 339500 3256 339552 3262
rect 339500 3198 339552 3204
rect 339512 480 339540 3198
rect 340524 3126 340552 5306
rect 340708 5250 340736 44118
rect 340788 41472 340840 41478
rect 340788 41414 340840 41420
rect 340800 5370 340828 41414
rect 340788 5364 340840 5370
rect 340788 5306 340840 5312
rect 340708 5222 340828 5250
rect 340800 3534 340828 5222
rect 341892 4072 341944 4078
rect 341892 4014 341944 4020
rect 340696 3528 340748 3534
rect 340696 3470 340748 3476
rect 340788 3528 340840 3534
rect 340788 3470 340840 3476
rect 340512 3120 340564 3126
rect 340512 3062 340564 3068
rect 340708 480 340736 3470
rect 341904 480 341932 4014
rect 342180 3262 342208 44118
rect 342732 41478 342760 44132
rect 343652 41478 343680 44132
rect 344664 42158 344692 44132
rect 345690 44118 346348 44146
rect 344652 42152 344704 42158
rect 344652 42094 344704 42100
rect 342720 41472 342772 41478
rect 342720 41414 342772 41420
rect 343548 41472 343600 41478
rect 343548 41414 343600 41420
rect 343640 41472 343692 41478
rect 343640 41414 343692 41420
rect 344928 41472 344980 41478
rect 344928 41414 344980 41420
rect 343560 3670 343588 41414
rect 344940 4078 344968 41414
rect 346320 4146 346348 44118
rect 346596 41478 346624 44132
rect 347608 42566 347636 44132
rect 348634 44118 349108 44146
rect 347596 42560 347648 42566
rect 347596 42502 347648 42508
rect 346584 41472 346636 41478
rect 346584 41414 346636 41420
rect 347688 41472 347740 41478
rect 347688 41414 347740 41420
rect 345480 4140 345532 4146
rect 345480 4082 345532 4088
rect 346308 4140 346360 4146
rect 346308 4082 346360 4088
rect 344928 4072 344980 4078
rect 344928 4014 344980 4020
rect 344284 4004 344336 4010
rect 344284 3946 344336 3952
rect 343088 3664 343140 3670
rect 343088 3606 343140 3612
rect 343548 3664 343600 3670
rect 343548 3606 343600 3612
rect 342168 3256 342220 3262
rect 342168 3198 342220 3204
rect 343100 480 343128 3606
rect 344296 480 344324 3946
rect 345492 480 345520 4082
rect 347700 3398 347728 41414
rect 349080 3942 349108 44118
rect 349540 41478 349568 44132
rect 350552 42090 350580 44132
rect 351578 44118 351868 44146
rect 352498 44118 353248 44146
rect 350540 42084 350592 42090
rect 350540 42026 350592 42032
rect 349528 41472 349580 41478
rect 349528 41414 349580 41420
rect 350448 41472 350500 41478
rect 350448 41414 350500 41420
rect 350460 4010 350488 41414
rect 350448 4004 350500 4010
rect 350448 3946 350500 3952
rect 347872 3936 347924 3942
rect 347872 3878 347924 3884
rect 349068 3936 349120 3942
rect 349068 3878 349120 3884
rect 346676 3392 346728 3398
rect 346676 3334 346728 3340
rect 347688 3392 347740 3398
rect 347688 3334 347740 3340
rect 346688 480 346716 3334
rect 347884 480 347912 3878
rect 351840 3330 351868 44118
rect 352564 3732 352616 3738
rect 352564 3674 352616 3680
rect 351368 3324 351420 3330
rect 351368 3266 351420 3272
rect 351828 3324 351880 3330
rect 351828 3266 351880 3272
rect 350264 3052 350316 3058
rect 350264 2994 350316 3000
rect 349068 2984 349120 2990
rect 349068 2926 349120 2932
rect 349080 480 349108 2926
rect 350276 480 350304 2994
rect 351380 480 351408 3266
rect 352576 480 352604 3674
rect 353220 3058 353248 44118
rect 353496 42430 353524 44132
rect 354522 44118 354628 44146
rect 355442 44118 356008 44146
rect 353484 42424 353536 42430
rect 353484 42366 353536 42372
rect 354600 3806 354628 44118
rect 355980 3874 356008 44118
rect 356440 42362 356468 44132
rect 356428 42356 356480 42362
rect 356428 42298 356480 42304
rect 357452 41478 357480 44132
rect 358386 44118 358676 44146
rect 357440 41472 357492 41478
rect 357440 41414 357492 41420
rect 354956 3868 355008 3874
rect 354956 3810 355008 3816
rect 355968 3868 356020 3874
rect 355968 3810 356020 3816
rect 353760 3800 353812 3806
rect 353760 3742 353812 3748
rect 354588 3800 354640 3806
rect 354588 3742 354640 3748
rect 353208 3052 353260 3058
rect 353208 2994 353260 3000
rect 353772 480 353800 3742
rect 354968 480 354996 3810
rect 358544 3596 358596 3602
rect 358544 3538 358596 3544
rect 357348 3460 357400 3466
rect 357348 3402 357400 3408
rect 356152 3188 356204 3194
rect 356152 3130 356204 3136
rect 356164 480 356192 3130
rect 357360 480 357388 3402
rect 358556 480 358584 3538
rect 358648 3466 358676 44118
rect 359384 42498 359412 44132
rect 359372 42492 359424 42498
rect 359372 42434 359424 42440
rect 360304 41478 360332 44132
rect 361330 44118 361436 44146
rect 358728 41472 358780 41478
rect 358728 41414 358780 41420
rect 360292 41472 360344 41478
rect 360292 41414 360344 41420
rect 358740 3738 358768 41414
rect 358728 3732 358780 3738
rect 358728 3674 358780 3680
rect 361408 3602 361436 44118
rect 362328 42294 362356 44132
rect 362316 42288 362368 42294
rect 362316 42230 362368 42236
rect 363248 41478 363276 44132
rect 364168 44118 364274 44146
rect 361488 41472 361540 41478
rect 361488 41414 361540 41420
rect 363236 41472 363288 41478
rect 363236 41414 363288 41420
rect 361396 3596 361448 3602
rect 361396 3538 361448 3544
rect 360936 3528 360988 3534
rect 360936 3470 360988 3476
rect 358636 3460 358688 3466
rect 358636 3402 358688 3408
rect 359740 3120 359792 3126
rect 359740 3062 359792 3068
rect 359752 480 359780 3062
rect 360948 480 360976 3470
rect 361500 3126 361528 41414
rect 363328 3664 363380 3670
rect 363328 3606 363380 3612
rect 362132 3256 362184 3262
rect 362132 3198 362184 3204
rect 361488 3120 361540 3126
rect 361488 3062 361540 3068
rect 362144 480 362172 3198
rect 363340 480 363368 3606
rect 364168 3534 364196 44118
rect 365272 42634 365300 44132
rect 365260 42628 365312 42634
rect 365260 42570 365312 42576
rect 365812 42152 365864 42158
rect 365812 42094 365864 42100
rect 364248 41472 364300 41478
rect 364248 41414 364300 41420
rect 364260 3670 364288 41414
rect 364524 4072 364576 4078
rect 364524 4014 364576 4020
rect 364248 3664 364300 3670
rect 364248 3606 364300 3612
rect 364156 3528 364208 3534
rect 364156 3470 364208 3476
rect 364536 480 364564 4014
rect 365824 3482 365852 42094
rect 366192 41478 366220 44132
rect 367204 41478 367232 44132
rect 368216 42226 368244 44132
rect 369150 44118 369808 44146
rect 368572 42560 368624 42566
rect 368572 42502 368624 42508
rect 368204 42220 368256 42226
rect 368204 42162 368256 42168
rect 366180 41472 366232 41478
rect 366180 41414 366232 41420
rect 367008 41472 367060 41478
rect 367008 41414 367060 41420
rect 367192 41472 367244 41478
rect 367192 41414 367244 41420
rect 368388 41472 368440 41478
rect 368388 41414 368440 41420
rect 366916 4140 366968 4146
rect 366916 4082 366968 4088
rect 365732 3454 365852 3482
rect 365732 480 365760 3454
rect 366928 480 366956 4082
rect 367020 3194 367048 41414
rect 368400 4146 368428 41414
rect 368388 4140 368440 4146
rect 368388 4082 368440 4088
rect 368020 3392 368072 3398
rect 368020 3334 368072 3340
rect 367008 3188 367060 3194
rect 367008 3130 367060 3136
rect 368032 480 368060 3334
rect 368584 610 368612 42502
rect 369780 3398 369808 44118
rect 370148 41478 370176 44132
rect 371160 42158 371188 44132
rect 372094 44118 372568 44146
rect 371148 42152 371200 42158
rect 371148 42094 371200 42100
rect 370136 41472 370188 41478
rect 370136 41414 370188 41420
rect 371148 41472 371200 41478
rect 371148 41414 371200 41420
rect 371160 4078 371188 41414
rect 371148 4072 371200 4078
rect 371148 4014 371200 4020
rect 371608 4004 371660 4010
rect 371608 3946 371660 3952
rect 370412 3936 370464 3942
rect 370412 3878 370464 3884
rect 369768 3392 369820 3398
rect 369768 3334 369820 3340
rect 368572 604 368624 610
rect 368572 546 368624 552
rect 369216 604 369268 610
rect 369216 546 369268 552
rect 369228 480 369256 546
rect 370424 480 370452 3878
rect 371620 480 371648 3946
rect 372540 3942 372568 44118
rect 372712 42084 372764 42090
rect 372712 42026 372764 42032
rect 372528 3936 372580 3942
rect 372528 3878 372580 3884
rect 372724 3482 372752 42026
rect 373092 41478 373120 44132
rect 374104 42566 374132 44132
rect 375038 44118 375328 44146
rect 376050 44118 376708 44146
rect 374092 42560 374144 42566
rect 374092 42502 374144 42508
rect 373080 41472 373132 41478
rect 373080 41414 373132 41420
rect 373908 41472 373960 41478
rect 373908 41414 373960 41420
rect 373920 4010 373948 41414
rect 373908 4004 373960 4010
rect 373908 3946 373960 3952
rect 372724 3454 372844 3482
rect 372816 480 372844 3454
rect 375300 3330 375328 44118
rect 375472 42424 375524 42430
rect 375472 42366 375524 42372
rect 374000 3324 374052 3330
rect 374000 3266 374052 3272
rect 375288 3324 375340 3330
rect 375288 3266 375340 3272
rect 374012 480 374040 3266
rect 375196 3052 375248 3058
rect 375196 2994 375248 3000
rect 375208 480 375236 2994
rect 375484 610 375512 42366
rect 376680 3262 376708 44118
rect 376956 42090 376984 44132
rect 377982 44118 378088 44146
rect 378994 44118 379468 44146
rect 376944 42084 376996 42090
rect 376944 42026 376996 42032
rect 378060 3806 378088 44118
rect 379440 3874 379468 44118
rect 379900 42430 379928 44132
rect 379888 42424 379940 42430
rect 379888 42366 379940 42372
rect 379520 42356 379572 42362
rect 379520 42298 379572 42304
rect 378784 3868 378836 3874
rect 378784 3810 378836 3816
rect 379428 3868 379480 3874
rect 379428 3810 379480 3816
rect 377588 3800 377640 3806
rect 377588 3742 377640 3748
rect 378048 3800 378100 3806
rect 378048 3742 378100 3748
rect 376668 3256 376720 3262
rect 376668 3198 376720 3204
rect 375472 604 375524 610
rect 375472 546 375524 552
rect 376392 604 376444 610
rect 376392 546 376444 552
rect 376404 480 376432 546
rect 377600 480 377628 3742
rect 378796 480 378824 3810
rect 379532 610 379560 42298
rect 380912 41478 380940 44132
rect 381938 44118 382136 44146
rect 380900 41472 380952 41478
rect 380900 41414 380952 41420
rect 382108 3738 382136 44118
rect 382844 42770 382872 44132
rect 382832 42764 382884 42770
rect 382832 42706 382884 42712
rect 382464 42492 382516 42498
rect 382464 42434 382516 42440
rect 382188 41472 382240 41478
rect 382188 41414 382240 41420
rect 381176 3732 381228 3738
rect 381176 3674 381228 3680
rect 382096 3732 382148 3738
rect 382096 3674 382148 3680
rect 379520 604 379572 610
rect 379520 546 379572 552
rect 379980 604 380032 610
rect 379980 546 380032 552
rect 379992 480 380020 546
rect 381188 480 381216 3674
rect 382200 2922 382228 41414
rect 382372 3460 382424 3466
rect 382372 3402 382424 3408
rect 382188 2916 382240 2922
rect 382188 2858 382240 2864
rect 382384 480 382412 3402
rect 382476 610 382504 42434
rect 383856 41478 383884 44132
rect 383844 41472 383896 41478
rect 383844 41414 383896 41420
rect 384868 3466 384896 44132
rect 385788 42362 385816 44132
rect 385776 42356 385828 42362
rect 385776 42298 385828 42304
rect 386512 42288 386564 42294
rect 386512 42230 386564 42236
rect 384948 41472 385000 41478
rect 384948 41414 385000 41420
rect 384856 3460 384908 3466
rect 384856 3402 384908 3408
rect 384672 3120 384724 3126
rect 384672 3062 384724 3068
rect 382464 604 382516 610
rect 382464 546 382516 552
rect 383568 604 383620 610
rect 383568 546 383620 552
rect 383580 480 383608 546
rect 384684 480 384712 3062
rect 384960 2990 384988 41414
rect 385868 3596 385920 3602
rect 385868 3538 385920 3544
rect 384948 2984 385000 2990
rect 384948 2926 385000 2932
rect 385880 480 385908 3538
rect 386524 610 386552 42230
rect 386800 41478 386828 44132
rect 387812 41478 387840 44132
rect 388732 42294 388760 44132
rect 388720 42288 388772 42294
rect 388720 42230 388772 42236
rect 389744 41478 389772 44132
rect 390652 42628 390704 42634
rect 390652 42570 390704 42576
rect 386788 41472 386840 41478
rect 386788 41414 386840 41420
rect 387708 41472 387760 41478
rect 387708 41414 387760 41420
rect 387800 41472 387852 41478
rect 387800 41414 387852 41420
rect 389088 41472 389140 41478
rect 389088 41414 389140 41420
rect 389732 41472 389784 41478
rect 389732 41414 389784 41420
rect 390468 41472 390520 41478
rect 390468 41414 390520 41420
rect 387720 3602 387748 41414
rect 388260 3664 388312 3670
rect 388260 3606 388312 3612
rect 387708 3596 387760 3602
rect 387708 3538 387760 3544
rect 386512 604 386564 610
rect 386512 546 386564 552
rect 387064 604 387116 610
rect 387064 546 387116 552
rect 387076 480 387104 546
rect 388272 480 388300 3606
rect 389100 3058 389128 41414
rect 390480 3670 390508 41414
rect 390468 3664 390520 3670
rect 390468 3606 390520 3612
rect 389456 3528 389508 3534
rect 389456 3470 389508 3476
rect 389088 3052 389140 3058
rect 389088 2994 389140 3000
rect 389468 480 389496 3470
rect 390664 480 390692 42570
rect 390756 41478 390784 44132
rect 391690 44118 391796 44146
rect 392702 44118 393268 44146
rect 390744 41472 390796 41478
rect 390744 41414 390796 41420
rect 391768 4826 391796 44118
rect 391848 41472 391900 41478
rect 391848 41414 391900 41420
rect 391756 4820 391808 4826
rect 391756 4762 391808 4768
rect 391860 4706 391888 41414
rect 391768 4678 391888 4706
rect 391768 3126 391796 4678
rect 393044 4140 393096 4146
rect 393044 4082 393096 4088
rect 391848 3188 391900 3194
rect 391848 3130 391900 3136
rect 391756 3120 391808 3126
rect 391756 3062 391808 3068
rect 391860 480 391888 3130
rect 393056 480 393084 4082
rect 393240 3534 393268 44118
rect 393504 42220 393556 42226
rect 393504 42162 393556 42168
rect 393228 3528 393280 3534
rect 393228 3470 393280 3476
rect 393516 610 393544 42162
rect 393608 41478 393636 44132
rect 394620 42022 394648 44132
rect 395646 44118 396028 44146
rect 394608 42016 394660 42022
rect 394608 41958 394660 41964
rect 393596 41472 393648 41478
rect 393596 41414 393648 41420
rect 394608 41472 394660 41478
rect 394608 41414 394660 41420
rect 394620 4146 394648 41414
rect 394608 4140 394660 4146
rect 394608 4082 394660 4088
rect 396000 4010 396028 44118
rect 396552 41546 396580 44132
rect 396540 41540 396592 41546
rect 396540 41482 396592 41488
rect 397564 41478 397592 44132
rect 398590 44118 398788 44146
rect 397644 42152 397696 42158
rect 397644 42094 397696 42100
rect 397552 41472 397604 41478
rect 397552 41414 397604 41420
rect 396632 4072 396684 4078
rect 396632 4014 396684 4020
rect 395988 4004 396040 4010
rect 395988 3946 396040 3952
rect 395436 3392 395488 3398
rect 395436 3334 395488 3340
rect 393504 604 393556 610
rect 393504 546 393556 552
rect 394240 604 394292 610
rect 394240 546 394292 552
rect 394252 480 394280 546
rect 395448 480 395476 3334
rect 396644 480 396672 4014
rect 397656 610 397684 42094
rect 398656 41472 398708 41478
rect 398656 41414 398708 41420
rect 398668 5234 398696 41414
rect 398656 5228 398708 5234
rect 398656 5170 398708 5176
rect 398760 4078 398788 44118
rect 399496 42702 399524 44132
rect 399484 42696 399536 42702
rect 399484 42638 399536 42644
rect 400404 42560 400456 42566
rect 400404 42502 400456 42508
rect 399484 41336 399536 41342
rect 399484 41278 399536 41284
rect 399496 31770 399524 41278
rect 399496 31742 399616 31770
rect 399588 26874 399616 31742
rect 399496 26846 399616 26874
rect 399496 12458 399524 26846
rect 399496 12430 399616 12458
rect 398748 4072 398800 4078
rect 398748 4014 398800 4020
rect 399024 3936 399076 3942
rect 399024 3878 399076 3884
rect 397644 604 397696 610
rect 397644 546 397696 552
rect 397828 604 397880 610
rect 397828 546 397880 552
rect 397840 480 397868 546
rect 399036 480 399064 3878
rect 399588 3126 399616 12430
rect 400220 3392 400272 3398
rect 400220 3334 400272 3340
rect 399576 3120 399628 3126
rect 399576 3062 399628 3068
rect 400232 480 400260 3334
rect 400416 610 400444 42502
rect 400508 42158 400536 44132
rect 400496 42152 400548 42158
rect 400496 42094 400548 42100
rect 401520 4010 401548 44132
rect 402244 42696 402296 42702
rect 402244 42638 402296 42644
rect 401508 4004 401560 4010
rect 401508 3946 401560 3952
rect 402256 3942 402284 42638
rect 402440 42498 402468 44132
rect 403452 42702 403480 44132
rect 404464 42702 404492 44132
rect 403440 42696 403492 42702
rect 403440 42638 403492 42644
rect 404268 42696 404320 42702
rect 404268 42638 404320 42644
rect 404452 42696 404504 42702
rect 404452 42638 404504 42644
rect 402428 42492 402480 42498
rect 402428 42434 402480 42440
rect 404280 5166 404308 42638
rect 405384 42634 405412 44132
rect 406410 44118 407068 44146
rect 405648 42696 405700 42702
rect 405648 42638 405700 42644
rect 405372 42628 405424 42634
rect 405372 42570 405424 42576
rect 404544 42084 404596 42090
rect 404544 42026 404596 42032
rect 404556 31770 404584 42026
rect 404556 31742 404676 31770
rect 404648 24426 404676 31742
rect 404648 24398 404768 24426
rect 404740 19310 404768 24398
rect 404728 19304 404780 19310
rect 404728 19246 404780 19252
rect 404452 9716 404504 9722
rect 404452 9658 404504 9664
rect 404268 5160 404320 5166
rect 404268 5102 404320 5108
rect 402244 3936 402296 3942
rect 402244 3878 402296 3884
rect 402796 3936 402848 3942
rect 402796 3878 402848 3884
rect 402808 3330 402836 3878
rect 402520 3324 402572 3330
rect 402520 3266 402572 3272
rect 402796 3324 402848 3330
rect 402796 3266 402848 3272
rect 400404 604 400456 610
rect 400404 546 400456 552
rect 401324 604 401376 610
rect 401324 546 401376 552
rect 401336 480 401364 546
rect 402532 480 402560 3266
rect 403716 3256 403768 3262
rect 403716 3198 403768 3204
rect 403728 480 403756 3198
rect 404464 678 404492 9658
rect 405660 3262 405688 42638
rect 407040 5098 407068 44118
rect 407408 42226 407436 44132
rect 407396 42220 407448 42226
rect 407396 42162 407448 42168
rect 408328 42090 408356 44132
rect 409354 44118 409828 44146
rect 408592 42424 408644 42430
rect 408592 42366 408644 42372
rect 408408 42220 408460 42226
rect 408408 42162 408460 42168
rect 408316 42084 408368 42090
rect 408316 42026 408368 42032
rect 407028 5092 407080 5098
rect 407028 5034 407080 5040
rect 407304 3868 407356 3874
rect 407304 3810 407356 3816
rect 406108 3800 406160 3806
rect 406108 3742 406160 3748
rect 405648 3256 405700 3262
rect 405648 3198 405700 3204
rect 404452 672 404504 678
rect 404452 614 404504 620
rect 404912 604 404964 610
rect 404912 546 404964 552
rect 404924 480 404952 546
rect 406120 480 406148 3742
rect 407316 480 407344 3810
rect 408420 3806 408448 42162
rect 408408 3800 408460 3806
rect 408408 3742 408460 3748
rect 408604 626 408632 42366
rect 409800 5030 409828 44118
rect 410260 41478 410288 44132
rect 411272 42566 411300 44132
rect 412298 44118 412588 44146
rect 413218 44118 413968 44146
rect 411444 42764 411496 42770
rect 411444 42706 411496 42712
rect 411260 42560 411312 42566
rect 411260 42502 411312 42508
rect 410248 41472 410300 41478
rect 410248 41414 410300 41420
rect 411168 41472 411220 41478
rect 411168 41414 411220 41420
rect 409788 5024 409840 5030
rect 409788 4966 409840 4972
rect 411180 3874 411208 41414
rect 411168 3868 411220 3874
rect 411168 3810 411220 3816
rect 410892 3732 410944 3738
rect 410892 3674 410944 3680
rect 409696 2916 409748 2922
rect 409696 2858 409748 2864
rect 408512 598 408632 626
rect 408512 480 408540 598
rect 409708 480 409736 2858
rect 410904 480 410932 3674
rect 411456 610 411484 42706
rect 412560 4894 412588 44118
rect 412548 4888 412600 4894
rect 412548 4830 412600 4836
rect 413940 3738 413968 44118
rect 414216 42770 414244 44132
rect 415242 44118 415348 44146
rect 416162 44118 416728 44146
rect 414204 42764 414256 42770
rect 414204 42706 414256 42712
rect 415320 4962 415348 44118
rect 415492 42356 415544 42362
rect 415492 42298 415544 42304
rect 415308 4956 415360 4962
rect 415308 4898 415360 4904
rect 413928 3732 413980 3738
rect 413928 3674 413980 3680
rect 414480 3460 414532 3466
rect 414480 3402 414532 3408
rect 413284 2984 413336 2990
rect 413284 2926 413336 2932
rect 411444 604 411496 610
rect 411444 546 411496 552
rect 412088 604 412140 610
rect 412088 546 412140 552
rect 412100 480 412128 546
rect 413296 480 413324 2926
rect 414492 480 414520 3402
rect 415504 610 415532 42298
rect 416700 3806 416728 44118
rect 417160 42498 417188 44132
rect 417424 42696 417476 42702
rect 417424 42638 417476 42644
rect 417148 42492 417200 42498
rect 417148 42434 417200 42440
rect 416688 3800 416740 3806
rect 416688 3742 416740 3748
rect 416872 3596 416924 3602
rect 416872 3538 416924 3544
rect 415492 604 415544 610
rect 415492 546 415544 552
rect 415676 604 415728 610
rect 415676 546 415728 552
rect 415688 480 415716 546
rect 416884 480 416912 3538
rect 417436 2854 417464 42638
rect 418172 42430 418200 44132
rect 419106 44118 419488 44146
rect 418160 42424 418212 42430
rect 418160 42366 418212 42372
rect 418252 42288 418304 42294
rect 418252 42230 418304 42236
rect 417976 3052 418028 3058
rect 417976 2994 418028 3000
rect 417424 2848 417476 2854
rect 417424 2790 417476 2796
rect 417988 480 418016 2994
rect 418264 610 418292 42230
rect 419460 3602 419488 44118
rect 420104 41478 420132 44132
rect 421116 41478 421144 44132
rect 422050 44118 422248 44146
rect 420092 41472 420144 41478
rect 420092 41414 420144 41420
rect 420828 41472 420880 41478
rect 420828 41414 420880 41420
rect 421104 41472 421156 41478
rect 421104 41414 421156 41420
rect 422116 41472 422168 41478
rect 422116 41414 422168 41420
rect 420840 3670 420868 41414
rect 422128 5370 422156 41414
rect 422116 5364 422168 5370
rect 422116 5306 422168 5312
rect 420368 3664 420420 3670
rect 420368 3606 420420 3612
rect 420828 3664 420880 3670
rect 420828 3606 420880 3612
rect 419448 3596 419500 3602
rect 419448 3538 419500 3544
rect 418252 604 418304 610
rect 418252 546 418304 552
rect 419172 604 419224 610
rect 419172 546 419224 552
rect 419184 480 419212 546
rect 420380 480 420408 3606
rect 422220 3466 422248 44118
rect 422944 42764 422996 42770
rect 422944 42706 422996 42712
rect 422760 4820 422812 4826
rect 422760 4762 422812 4768
rect 422208 3460 422260 3466
rect 422208 3402 422260 3408
rect 421564 3188 421616 3194
rect 421564 3130 421616 3136
rect 421576 480 421604 3130
rect 422772 480 422800 4762
rect 422956 2990 422984 42706
rect 423048 42294 423076 44132
rect 423036 42288 423088 42294
rect 423036 42230 423088 42236
rect 424060 41478 424088 44132
rect 424048 41472 424100 41478
rect 424048 41414 424100 41420
rect 424876 41472 424928 41478
rect 424876 41414 424928 41420
rect 424888 4826 424916 41414
rect 424876 4820 424928 4826
rect 424876 4762 424928 4768
rect 424980 3534 425008 44132
rect 425992 42226 426020 44132
rect 425980 42220 426032 42226
rect 425980 42162 426032 42168
rect 425244 42016 425296 42022
rect 425244 41958 425296 41964
rect 425152 4140 425204 4146
rect 425152 4082 425204 4088
rect 423956 3528 424008 3534
rect 423956 3470 424008 3476
rect 424968 3528 425020 3534
rect 424968 3470 425020 3476
rect 422944 2984 422996 2990
rect 422944 2926 422996 2932
rect 423968 480 423996 3470
rect 425164 480 425192 4082
rect 425256 610 425284 41958
rect 426912 41478 426940 44132
rect 427924 41478 427952 44132
rect 428936 42362 428964 44132
rect 429870 44118 430528 44146
rect 428924 42356 428976 42362
rect 428924 42298 428976 42304
rect 426900 41472 426952 41478
rect 426900 41414 426952 41420
rect 427728 41472 427780 41478
rect 427728 41414 427780 41420
rect 427912 41472 427964 41478
rect 427912 41414 427964 41420
rect 429108 41472 429160 41478
rect 429108 41414 429160 41420
rect 427740 4146 427768 41414
rect 427728 4140 427780 4146
rect 427728 4082 427780 4088
rect 429120 4010 429148 41414
rect 429936 5228 429988 5234
rect 429936 5170 429988 5176
rect 429108 4004 429160 4010
rect 429108 3946 429160 3952
rect 427544 3392 427596 3398
rect 427544 3334 427596 3340
rect 425244 604 425296 610
rect 425244 546 425296 552
rect 426348 604 426400 610
rect 426348 546 426400 552
rect 426360 480 426388 546
rect 427556 480 427584 3334
rect 428740 3120 428792 3126
rect 428740 3062 428792 3068
rect 428752 480 428780 3062
rect 429948 480 429976 5170
rect 430500 3058 430528 44118
rect 430868 41478 430896 44132
rect 431788 44118 431894 44146
rect 432814 44118 433288 44146
rect 430856 41472 430908 41478
rect 430856 41414 430908 41420
rect 431132 4072 431184 4078
rect 431132 4014 431184 4020
rect 430488 3052 430540 3058
rect 430488 2994 430540 3000
rect 431144 480 431172 4014
rect 431788 3126 431816 44118
rect 431868 41472 431920 41478
rect 431868 41414 431920 41420
rect 431776 3120 431828 3126
rect 431776 3062 431828 3068
rect 431880 2990 431908 41414
rect 433260 4010 433288 44118
rect 433432 42152 433484 42158
rect 433432 42094 433484 42100
rect 433444 37262 433472 42094
rect 433812 41478 433840 44132
rect 433984 42628 434036 42634
rect 433984 42570 434036 42576
rect 433800 41472 433852 41478
rect 433800 41414 433852 41420
rect 433432 37256 433484 37262
rect 433432 37198 433484 37204
rect 433432 27668 433484 27674
rect 433432 27610 433484 27616
rect 433444 17950 433472 27610
rect 433432 17944 433484 17950
rect 433432 17886 433484 17892
rect 433432 8424 433484 8430
rect 433432 8366 433484 8372
rect 433444 8294 433472 8366
rect 433432 8288 433484 8294
rect 433432 8230 433484 8236
rect 433996 4146 434024 42570
rect 434824 41750 434852 44132
rect 435758 44118 436048 44146
rect 434812 41744 434864 41750
rect 434812 41686 434864 41692
rect 434628 41472 434680 41478
rect 434628 41414 434680 41420
rect 434640 7834 434668 41414
rect 434548 7806 434668 7834
rect 433984 4140 434036 4146
rect 433984 4082 434036 4088
rect 433248 4004 433300 4010
rect 433248 3946 433300 3952
rect 432328 3324 432380 3330
rect 432328 3266 432380 3272
rect 431868 2984 431920 2990
rect 431868 2926 431920 2932
rect 432340 480 432368 3266
rect 434548 3194 434576 7806
rect 436020 4146 436048 44118
rect 436756 41546 436784 44132
rect 436744 41540 436796 41546
rect 436744 41482 436796 41488
rect 437768 41478 437796 44132
rect 437756 41472 437808 41478
rect 437756 41414 437808 41420
rect 437020 5160 437072 5166
rect 437020 5102 437072 5108
rect 435824 4140 435876 4146
rect 435824 4082 435876 4088
rect 436008 4140 436060 4146
rect 436008 4082 436060 4088
rect 434628 3392 434680 3398
rect 434628 3334 434680 3340
rect 434536 3188 434588 3194
rect 434536 3130 434588 3136
rect 433524 604 433576 610
rect 433524 546 433576 552
rect 433536 480 433564 546
rect 434640 480 434668 3334
rect 435836 480 435864 4082
rect 437032 480 437060 5102
rect 438688 4010 438716 44132
rect 439714 44118 440188 44146
rect 438768 41472 438820 41478
rect 438768 41414 438820 41420
rect 438676 4004 438728 4010
rect 438676 3946 438728 3952
rect 438780 3330 438808 41414
rect 440160 4078 440188 44118
rect 440712 41682 440740 44132
rect 440700 41676 440752 41682
rect 440700 41618 440752 41624
rect 441632 41478 441660 44132
rect 442658 44118 442948 44146
rect 441620 41472 441672 41478
rect 441620 41414 441672 41420
rect 442816 41472 442868 41478
rect 442816 41414 442868 41420
rect 442828 5166 442856 41414
rect 442816 5160 442868 5166
rect 442816 5102 442868 5108
rect 440608 5092 440660 5098
rect 440608 5034 440660 5040
rect 440148 4072 440200 4078
rect 440148 4014 440200 4020
rect 438768 3324 438820 3330
rect 438768 3266 438820 3272
rect 438216 3256 438268 3262
rect 438216 3198 438268 3204
rect 438228 480 438256 3198
rect 439412 2304 439464 2310
rect 439412 2246 439464 2252
rect 439424 480 439452 2246
rect 440620 480 440648 5034
rect 441804 3936 441856 3942
rect 441804 3878 441856 3884
rect 441434 3088 441490 3097
rect 441434 3023 441436 3032
rect 441488 3023 441490 3032
rect 441436 2994 441488 3000
rect 441816 480 441844 3878
rect 442920 3369 442948 44118
rect 443564 42158 443592 44132
rect 443552 42152 443604 42158
rect 443552 42094 443604 42100
rect 443000 42084 443052 42090
rect 443000 42026 443052 42032
rect 442906 3360 442962 3369
rect 442264 3324 442316 3330
rect 442906 3295 442962 3304
rect 442264 3266 442316 3272
rect 442276 3194 442304 3266
rect 442264 3188 442316 3194
rect 442264 3130 442316 3136
rect 443012 480 443040 42026
rect 443644 41540 443696 41546
rect 443644 41482 443696 41488
rect 443656 3942 443684 41482
rect 444576 41478 444604 44132
rect 445588 42090 445616 44132
rect 445760 42560 445812 42566
rect 445760 42502 445812 42508
rect 445576 42084 445628 42090
rect 445576 42026 445628 42032
rect 444564 41472 444616 41478
rect 444564 41414 444616 41420
rect 445668 41472 445720 41478
rect 445668 41414 445720 41420
rect 445680 5234 445708 41414
rect 445668 5228 445720 5234
rect 445668 5170 445720 5176
rect 444196 5024 444248 5030
rect 444196 4966 444248 4972
rect 443644 3936 443696 3942
rect 443644 3878 443696 3884
rect 444208 480 444236 4966
rect 445392 3868 445444 3874
rect 445392 3810 445444 3816
rect 445404 480 445432 3810
rect 445772 610 445800 42502
rect 446508 41886 446536 44132
rect 446496 41880 446548 41886
rect 446496 41822 446548 41828
rect 447520 41478 447548 44132
rect 448532 41478 448560 44132
rect 449466 44118 449848 44146
rect 447508 41472 447560 41478
rect 447508 41414 447560 41420
rect 448428 41472 448480 41478
rect 448428 41414 448480 41420
rect 448520 41472 448572 41478
rect 448520 41414 448572 41420
rect 449716 41472 449768 41478
rect 449716 41414 449768 41420
rect 448440 5098 448468 41414
rect 448428 5092 448480 5098
rect 448428 5034 448480 5040
rect 447784 4888 447836 4894
rect 447784 4830 447836 4836
rect 447046 3088 447102 3097
rect 447046 3023 447102 3032
rect 447060 2990 447088 3023
rect 447048 2984 447100 2990
rect 447048 2926 447100 2932
rect 445760 604 445812 610
rect 445760 546 445812 552
rect 446588 604 446640 610
rect 446588 546 446640 552
rect 446600 480 446628 546
rect 447796 480 447824 4830
rect 449728 3806 449756 41414
rect 449820 3942 449848 44118
rect 450464 41478 450492 44132
rect 451476 41478 451504 44132
rect 452396 42634 452424 44132
rect 453422 44118 453988 44146
rect 452384 42628 452436 42634
rect 452384 42570 452436 42576
rect 451924 42492 451976 42498
rect 451924 42434 451976 42440
rect 450452 41472 450504 41478
rect 450452 41414 450504 41420
rect 451188 41472 451240 41478
rect 451188 41414 451240 41420
rect 451464 41472 451516 41478
rect 451464 41414 451516 41420
rect 451200 4894 451228 41414
rect 451280 4956 451332 4962
rect 451280 4898 451332 4904
rect 451188 4888 451240 4894
rect 451188 4830 451240 4836
rect 449808 3936 449860 3942
rect 449808 3878 449860 3884
rect 449716 3800 449768 3806
rect 449716 3742 449768 3748
rect 448980 3732 449032 3738
rect 448980 3674 449032 3680
rect 448992 480 449020 3674
rect 450176 2848 450228 2854
rect 450176 2790 450228 2796
rect 450188 480 450216 2790
rect 451292 480 451320 4898
rect 451936 3942 451964 42434
rect 452568 41472 452620 41478
rect 452568 41414 452620 41420
rect 451924 3936 451976 3942
rect 451924 3878 451976 3884
rect 452476 3868 452528 3874
rect 452476 3810 452528 3816
rect 452488 480 452516 3810
rect 452580 3466 452608 41414
rect 453960 5030 453988 44118
rect 454132 42424 454184 42430
rect 454132 42366 454184 42372
rect 453948 5024 454000 5030
rect 453948 4966 454000 4972
rect 453672 3936 453724 3942
rect 453672 3878 453724 3884
rect 452568 3460 452620 3466
rect 452568 3402 452620 3408
rect 453684 480 453712 3878
rect 454144 610 454172 42366
rect 454420 41478 454448 44132
rect 455340 42770 455368 44132
rect 456366 44118 456748 44146
rect 457378 44118 458128 44146
rect 455328 42764 455380 42770
rect 455328 42706 455380 42712
rect 454408 41472 454460 41478
rect 454408 41414 454460 41420
rect 455328 41472 455380 41478
rect 455328 41414 455380 41420
rect 455340 3806 455368 41414
rect 456720 5302 456748 44118
rect 456708 5296 456760 5302
rect 456708 5238 456760 5244
rect 457260 3936 457312 3942
rect 457260 3878 457312 3884
rect 455328 3800 455380 3806
rect 455328 3742 455380 3748
rect 456064 3596 456116 3602
rect 456064 3538 456116 3544
rect 454132 604 454184 610
rect 454132 546 454184 552
rect 454868 604 454920 610
rect 454868 546 454920 552
rect 454880 480 454908 546
rect 456076 480 456104 3538
rect 457272 480 457300 3878
rect 458100 3602 458128 44118
rect 458284 41954 458312 44132
rect 459310 44118 459508 44146
rect 460230 44118 460888 44146
rect 458272 41948 458324 41954
rect 458272 41890 458324 41896
rect 458456 4956 458508 4962
rect 458456 4898 458508 4904
rect 458088 3596 458140 3602
rect 458088 3538 458140 3544
rect 458468 480 458496 4898
rect 459480 4758 459508 44118
rect 459652 42288 459704 42294
rect 459652 42230 459704 42236
rect 459468 4752 459520 4758
rect 459468 4694 459520 4700
rect 459560 3664 459612 3670
rect 459560 3606 459612 3612
rect 459572 3346 459600 3606
rect 459664 3466 459692 42230
rect 460860 3602 460888 44118
rect 461228 42702 461256 44132
rect 461216 42696 461268 42702
rect 461216 42638 461268 42644
rect 462240 4826 462268 44132
rect 462964 42220 463016 42226
rect 462964 42162 463016 42168
rect 462044 4820 462096 4826
rect 462044 4762 462096 4768
rect 462228 4820 462280 4826
rect 462228 4762 462280 4768
rect 460848 3596 460900 3602
rect 460848 3538 460900 3544
rect 459652 3460 459704 3466
rect 459652 3402 459704 3408
rect 460848 3460 460900 3466
rect 460848 3402 460900 3408
rect 459572 3318 459692 3346
rect 459664 480 459692 3318
rect 460860 480 460888 3402
rect 462056 480 462084 4762
rect 462976 3534 463004 42162
rect 463160 41818 463188 44132
rect 464172 42022 464200 44132
rect 464344 42356 464396 42362
rect 464344 42298 464396 42304
rect 464160 42016 464212 42022
rect 464160 41958 464212 41964
rect 463148 41812 463200 41818
rect 463148 41754 463200 41760
rect 462964 3528 463016 3534
rect 462964 3470 463016 3476
rect 464356 3466 464384 42298
rect 465184 41478 465212 44132
rect 466118 44118 466408 44146
rect 465172 41472 465224 41478
rect 465172 41414 465224 41420
rect 466276 41472 466328 41478
rect 466276 41414 466328 41420
rect 466288 5506 466316 41414
rect 466276 5500 466328 5506
rect 466276 5442 466328 5448
rect 466380 3534 466408 44118
rect 467116 42498 467144 44132
rect 467104 42492 467156 42498
rect 467104 42434 467156 42440
rect 467104 41744 467156 41750
rect 467104 41686 467156 41692
rect 464436 3528 464488 3534
rect 464436 3470 464488 3476
rect 466368 3528 466420 3534
rect 466368 3470 466420 3476
rect 463240 3460 463292 3466
rect 463240 3402 463292 3408
rect 464344 3460 464396 3466
rect 464344 3402 464396 3408
rect 463252 480 463280 3402
rect 464448 480 464476 3470
rect 467116 3126 467144 41686
rect 468128 41478 468156 44132
rect 469048 42294 469076 44132
rect 470074 44118 470548 44146
rect 469036 42288 469088 42294
rect 469036 42230 469088 42236
rect 468484 41676 468536 41682
rect 468484 41618 468536 41624
rect 468116 41472 468168 41478
rect 468116 41414 468168 41420
rect 468496 3466 468524 41618
rect 469128 41472 469180 41478
rect 469128 41414 469180 41420
rect 469140 6186 469168 41414
rect 469128 6180 469180 6186
rect 469128 6122 469180 6128
rect 470520 3466 470548 44118
rect 471072 41478 471100 44132
rect 471992 42566 472020 44132
rect 471980 42560 472032 42566
rect 471980 42502 472032 42508
rect 473004 42362 473032 44132
rect 474030 44118 474688 44146
rect 472992 42356 473044 42362
rect 472992 42298 473044 42304
rect 471060 41472 471112 41478
rect 471060 41414 471112 41420
rect 471888 41472 471940 41478
rect 471888 41414 471940 41420
rect 471900 6594 471928 41414
rect 471888 6588 471940 6594
rect 471888 6530 471940 6536
rect 474660 6526 474688 44118
rect 474936 41478 474964 44132
rect 475948 41750 475976 44132
rect 476882 44118 477448 44146
rect 475936 41744 475988 41750
rect 475936 41686 475988 41692
rect 474924 41472 474976 41478
rect 474924 41414 474976 41420
rect 476028 41472 476080 41478
rect 476028 41414 476080 41420
rect 474648 6520 474700 6526
rect 474648 6462 474700 6468
rect 467932 3460 467984 3466
rect 467932 3402 467984 3408
rect 468484 3460 468536 3466
rect 468484 3402 468536 3408
rect 470508 3460 470560 3466
rect 470508 3402 470560 3408
rect 466828 3120 466880 3126
rect 466828 3062 466880 3068
rect 467104 3120 467156 3126
rect 467104 3062 467156 3068
rect 465632 2916 465684 2922
rect 465632 2858 465684 2864
rect 465644 480 465672 2858
rect 466840 480 466868 3062
rect 467944 480 467972 3402
rect 471520 3392 471572 3398
rect 471520 3334 471572 3340
rect 470324 3052 470376 3058
rect 470324 2994 470376 3000
rect 469128 2984 469180 2990
rect 469128 2926 469180 2932
rect 469140 480 469168 2926
rect 470336 480 470364 2994
rect 471532 480 471560 3334
rect 476040 3330 476068 41414
rect 477420 6458 477448 44118
rect 477880 42226 477908 44132
rect 478892 42294 478920 44132
rect 479826 44118 480208 44146
rect 478144 42288 478196 42294
rect 478144 42230 478196 42236
rect 478880 42288 478932 42294
rect 478880 42230 478932 42236
rect 477868 42220 477920 42226
rect 477868 42162 477920 42168
rect 477408 6452 477460 6458
rect 477408 6394 477460 6400
rect 476304 4140 476356 4146
rect 476304 4082 476356 4088
rect 473912 3324 473964 3330
rect 473912 3266 473964 3272
rect 476028 3324 476080 3330
rect 476028 3266 476080 3272
rect 472716 3188 472768 3194
rect 472716 3130 472768 3136
rect 472728 480 472756 3130
rect 473924 480 473952 3266
rect 475108 3120 475160 3126
rect 475108 3062 475160 3068
rect 475120 480 475148 3062
rect 476316 480 476344 4082
rect 478156 3058 478184 42230
rect 480180 5438 480208 44118
rect 480824 41478 480852 44132
rect 481836 41478 481864 44132
rect 482770 44118 482876 44146
rect 480812 41472 480864 41478
rect 480812 41414 480864 41420
rect 481548 41472 481600 41478
rect 481548 41414 481600 41420
rect 481824 41472 481876 41478
rect 481824 41414 481876 41420
rect 480168 5432 480220 5438
rect 480168 5374 480220 5380
rect 481088 4072 481140 4078
rect 481088 4014 481140 4020
rect 479892 4004 479944 4010
rect 479892 3946 479944 3952
rect 478696 3256 478748 3262
rect 478696 3198 478748 3204
rect 478144 3052 478196 3058
rect 478144 2994 478196 3000
rect 477500 2848 477552 2854
rect 477500 2790 477552 2796
rect 477512 480 477540 2790
rect 478708 480 478736 3198
rect 479904 480 479932 3946
rect 481100 480 481128 4014
rect 481560 3126 481588 41414
rect 482848 5302 482876 44118
rect 483664 42560 483716 42566
rect 483664 42502 483716 42508
rect 482928 41472 482980 41478
rect 482928 41414 482980 41420
rect 482836 5296 482888 5302
rect 482836 5238 482888 5244
rect 482940 3194 482968 41414
rect 483480 5160 483532 5166
rect 483480 5102 483532 5108
rect 482928 3188 482980 3194
rect 482928 3130 482980 3136
rect 481548 3120 481600 3126
rect 481548 3062 481600 3068
rect 482284 2984 482336 2990
rect 482284 2926 482336 2932
rect 482296 480 482324 2926
rect 483492 480 483520 5102
rect 483676 2990 483704 42502
rect 483768 42430 483796 44132
rect 483756 42424 483808 42430
rect 483756 42366 483808 42372
rect 484780 42090 484808 44132
rect 483756 42084 483808 42090
rect 483756 42026 483808 42032
rect 484768 42084 484820 42090
rect 484768 42026 484820 42032
rect 483768 3262 483796 42026
rect 485700 5166 485728 44132
rect 486712 42566 486740 44132
rect 487738 44118 488488 44146
rect 486700 42560 486752 42566
rect 486700 42502 486752 42508
rect 485780 42152 485832 42158
rect 485780 42094 485832 42100
rect 485688 5160 485740 5166
rect 485688 5102 485740 5108
rect 484582 3360 484638 3369
rect 484582 3295 484638 3304
rect 483756 3256 483808 3262
rect 483756 3198 483808 3204
rect 483664 2984 483716 2990
rect 483664 2926 483716 2932
rect 484596 480 484624 3295
rect 485792 480 485820 42094
rect 486424 41880 486476 41886
rect 486424 41822 486476 41828
rect 486436 3398 486464 41822
rect 486976 5228 487028 5234
rect 486976 5170 487028 5176
rect 486424 3392 486476 3398
rect 486424 3334 486476 3340
rect 486988 480 487016 5170
rect 488460 3262 488488 44118
rect 488644 41478 488672 44132
rect 489670 44118 489868 44146
rect 488632 41472 488684 41478
rect 488632 41414 488684 41420
rect 489736 41472 489788 41478
rect 489736 41414 489788 41420
rect 489748 5370 489776 41414
rect 489736 5364 489788 5370
rect 489736 5306 489788 5312
rect 489840 3398 489868 44118
rect 490668 42158 490696 44132
rect 490656 42152 490708 42158
rect 490656 42094 490708 42100
rect 491588 41478 491616 44132
rect 491576 41472 491628 41478
rect 491576 41414 491628 41420
rect 492496 41472 492548 41478
rect 492496 41414 492548 41420
rect 492508 5098 492536 41414
rect 490564 5092 490616 5098
rect 490564 5034 490616 5040
rect 492496 5092 492548 5098
rect 492496 5034 492548 5040
rect 489368 3392 489420 3398
rect 489368 3334 489420 3340
rect 489828 3392 489880 3398
rect 489828 3334 489880 3340
rect 488172 3256 488224 3262
rect 488172 3198 488224 3204
rect 488448 3256 488500 3262
rect 488448 3198 488500 3204
rect 488184 480 488212 3198
rect 489380 480 489408 3334
rect 490576 480 490604 5034
rect 492600 4078 492628 44132
rect 493534 44118 494008 44146
rect 492588 4072 492640 4078
rect 492588 4014 492640 4020
rect 493980 4010 494008 44118
rect 494532 41478 494560 44132
rect 494704 42628 494756 42634
rect 494704 42570 494756 42576
rect 494520 41472 494572 41478
rect 494520 41414 494572 41420
rect 494152 4888 494204 4894
rect 494152 4830 494204 4836
rect 493968 4004 494020 4010
rect 493968 3946 494020 3952
rect 491760 3868 491812 3874
rect 491760 3810 491812 3816
rect 491772 480 491800 3810
rect 492956 3732 493008 3738
rect 492956 3674 493008 3680
rect 492968 480 492996 3674
rect 494164 480 494192 4830
rect 494716 3738 494744 42570
rect 495544 41886 495572 44132
rect 496464 42634 496492 44132
rect 497490 44118 498148 44146
rect 496452 42628 496504 42634
rect 496452 42570 496504 42576
rect 495532 41880 495584 41886
rect 495532 41822 495584 41828
rect 496084 41744 496136 41750
rect 496084 41686 496136 41692
rect 495348 41472 495400 41478
rect 495348 41414 495400 41420
rect 495360 5234 495388 41414
rect 495348 5228 495400 5234
rect 495348 5170 495400 5176
rect 495348 3936 495400 3942
rect 495348 3878 495400 3884
rect 494704 3732 494756 3738
rect 494704 3674 494756 3680
rect 495360 480 495388 3878
rect 496096 2922 496124 41686
rect 498120 5030 498148 44118
rect 498488 41478 498516 44132
rect 498476 41472 498528 41478
rect 498476 41414 498528 41420
rect 497740 5024 497792 5030
rect 497740 4966 497792 4972
rect 498108 5024 498160 5030
rect 498108 4966 498160 4972
rect 496544 3732 496596 3738
rect 496544 3674 496596 3680
rect 496084 2916 496136 2922
rect 496084 2858 496136 2864
rect 496556 480 496584 3674
rect 497752 480 497780 4966
rect 499408 3806 499436 44132
rect 500434 44118 500908 44146
rect 499672 42764 499724 42770
rect 499672 42706 499724 42712
rect 499488 41472 499540 41478
rect 499488 41414 499540 41420
rect 499500 4146 499528 41414
rect 499488 4140 499540 4146
rect 499488 4082 499540 4088
rect 498936 3800 498988 3806
rect 498936 3742 498988 3748
rect 499396 3800 499448 3806
rect 499396 3742 499448 3748
rect 498948 480 498976 3742
rect 499684 610 499712 42706
rect 500880 4894 500908 44118
rect 501432 41750 501460 44132
rect 502352 42770 502380 44132
rect 503378 44118 503668 44146
rect 504390 44118 505048 44146
rect 502340 42764 502392 42770
rect 502340 42706 502392 42712
rect 502432 41948 502484 41954
rect 502432 41890 502484 41896
rect 501604 41812 501656 41818
rect 501604 41754 501656 41760
rect 501420 41744 501472 41750
rect 501420 41686 501472 41692
rect 501236 4956 501288 4962
rect 501236 4898 501288 4904
rect 500868 4888 500920 4894
rect 500868 4830 500920 4836
rect 499672 604 499724 610
rect 499672 546 499724 552
rect 500132 604 500184 610
rect 500132 546 500184 552
rect 500144 480 500172 546
rect 501248 480 501276 4898
rect 501616 3874 501644 41754
rect 501604 3868 501656 3874
rect 501604 3810 501656 3816
rect 502444 3738 502472 41890
rect 503640 4962 503668 44118
rect 503628 4956 503680 4962
rect 503628 4898 503680 4904
rect 504824 4752 504876 4758
rect 504824 4694 504876 4700
rect 502432 3732 502484 3738
rect 502432 3674 502484 3680
rect 503628 3732 503680 3738
rect 503628 3674 503680 3680
rect 502340 3664 502392 3670
rect 502340 3606 502392 3612
rect 502352 3482 502380 3606
rect 502352 3454 502472 3482
rect 502444 480 502472 3454
rect 503640 480 503668 3674
rect 504836 480 504864 4694
rect 505020 3738 505048 44118
rect 505296 41478 505324 44132
rect 505284 41472 505336 41478
rect 505284 41414 505336 41420
rect 506308 6254 506336 44132
rect 506480 42696 506532 42702
rect 506480 42638 506532 42644
rect 506388 41472 506440 41478
rect 506388 41414 506440 41420
rect 506296 6248 506348 6254
rect 506296 6190 506348 6196
rect 506400 3874 506428 41414
rect 506388 3868 506440 3874
rect 506388 3810 506440 3816
rect 505008 3732 505060 3738
rect 505008 3674 505060 3680
rect 506020 3664 506072 3670
rect 506020 3606 506072 3612
rect 506032 480 506060 3606
rect 506492 610 506520 42638
rect 507320 41954 507348 44132
rect 508240 42702 508268 44132
rect 508228 42696 508280 42702
rect 508228 42638 508280 42644
rect 508504 42016 508556 42022
rect 508504 41958 508556 41964
rect 507308 41948 507360 41954
rect 507308 41890 507360 41896
rect 508412 4820 508464 4826
rect 508412 4762 508464 4768
rect 506480 604 506532 610
rect 506480 546 506532 552
rect 507216 604 507268 610
rect 507216 546 507268 552
rect 507228 480 507256 546
rect 508424 480 508452 4762
rect 508516 3942 508544 41958
rect 509252 41478 509280 44132
rect 510186 44118 510568 44146
rect 509240 41472 509292 41478
rect 509240 41414 509292 41420
rect 510436 41472 510488 41478
rect 510436 41414 510488 41420
rect 510448 4826 510476 41414
rect 510436 4820 510488 4826
rect 510436 4762 510488 4768
rect 508504 3936 508556 3942
rect 508504 3878 508556 3884
rect 509608 3732 509660 3738
rect 509608 3674 509660 3680
rect 509620 480 509648 3674
rect 510540 2854 510568 44118
rect 511184 41478 511212 44132
rect 512196 41478 512224 44132
rect 512644 42492 512696 42498
rect 512644 42434 512696 42440
rect 511172 41472 511224 41478
rect 511172 41414 511224 41420
rect 511908 41472 511960 41478
rect 511908 41414 511960 41420
rect 512184 41472 512236 41478
rect 512184 41414 512236 41420
rect 510804 3936 510856 3942
rect 510804 3878 510856 3884
rect 510528 2848 510580 2854
rect 510528 2790 510580 2796
rect 510816 480 510844 3878
rect 511920 3738 511948 41414
rect 512000 5500 512052 5506
rect 512000 5442 512052 5448
rect 511908 3732 511960 3738
rect 511908 3674 511960 3680
rect 512012 480 512040 5442
rect 512656 3534 512684 42434
rect 513116 41818 513144 44132
rect 514128 42498 514156 44132
rect 514116 42492 514168 42498
rect 514116 42434 514168 42440
rect 513104 41812 513156 41818
rect 513104 41754 513156 41760
rect 515140 41478 515168 44132
rect 513288 41472 513340 41478
rect 513288 41414 513340 41420
rect 515128 41472 515180 41478
rect 515128 41414 515180 41420
rect 515956 41472 516008 41478
rect 515956 41414 516008 41420
rect 513300 6390 513328 41414
rect 513288 6384 513340 6390
rect 513288 6326 513340 6332
rect 515968 6322 515996 41414
rect 515956 6316 516008 6322
rect 515956 6258 516008 6264
rect 515588 6180 515640 6186
rect 515588 6122 515640 6128
rect 512644 3528 512696 3534
rect 512644 3470 512696 3476
rect 514392 3528 514444 3534
rect 514392 3470 514444 3476
rect 513196 3460 513248 3466
rect 513196 3402 513248 3408
rect 513208 480 513236 3402
rect 514404 480 514432 3470
rect 515600 480 515628 6122
rect 516060 3670 516088 44132
rect 517086 44118 517468 44146
rect 518098 44118 518848 44146
rect 516048 3664 516100 3670
rect 516048 3606 516100 3612
rect 517440 3534 517468 44118
rect 518820 6186 518848 44118
rect 519004 41682 519032 44132
rect 520016 42022 520044 44132
rect 520464 42356 520516 42362
rect 520464 42298 520516 42304
rect 520004 42016 520056 42022
rect 520004 41958 520056 41964
rect 518992 41676 519044 41682
rect 518992 41618 519044 41624
rect 519084 6588 519136 6594
rect 519084 6530 519136 6536
rect 518808 6180 518860 6186
rect 518808 6122 518860 6128
rect 517888 3596 517940 3602
rect 517888 3538 517940 3544
rect 517428 3528 517480 3534
rect 517428 3470 517480 3476
rect 516784 3052 516836 3058
rect 516784 2994 516836 3000
rect 516796 480 516824 2994
rect 517900 480 517928 3538
rect 519096 480 519124 6530
rect 520476 3482 520504 42298
rect 521028 41614 521056 44132
rect 521016 41608 521068 41614
rect 521016 41550 521068 41556
rect 521948 41478 521976 44132
rect 521936 41472 521988 41478
rect 521936 41414 521988 41420
rect 522316 17950 522344 643146
rect 522408 66178 522436 643282
rect 522500 111790 522528 644778
rect 522592 158710 522620 644914
rect 522684 452606 522712 647022
rect 525524 646944 525576 646950
rect 525524 646886 525576 646892
rect 580262 646912 580318 646921
rect 525340 646740 525392 646746
rect 525340 646682 525392 646688
rect 525248 646604 525300 646610
rect 525248 646546 525300 646552
rect 524144 645448 524196 645454
rect 524144 645390 524196 645396
rect 523960 645108 524012 645114
rect 523960 645050 524012 645056
rect 523408 644428 523460 644434
rect 523408 644370 523460 644376
rect 523420 627910 523448 644370
rect 523500 644360 523552 644366
rect 523500 644302 523552 644308
rect 523408 627904 523460 627910
rect 523408 627846 523460 627852
rect 523420 627803 523448 627846
rect 523512 580990 523540 644302
rect 523592 644292 523644 644298
rect 523592 644234 523644 644240
rect 523500 580984 523552 580990
rect 523500 580926 523552 580932
rect 523604 534070 523632 644234
rect 523868 643544 523920 643550
rect 523868 643486 523920 643492
rect 523776 643408 523828 643414
rect 523776 643350 523828 643356
rect 523682 642696 523738 642705
rect 523682 642631 523738 642640
rect 523592 534064 523644 534070
rect 523592 534006 523644 534012
rect 522672 452600 522724 452606
rect 522672 452542 522724 452548
rect 522580 158704 522632 158710
rect 522580 158646 522632 158652
rect 523696 135250 523724 642631
rect 523788 182170 523816 643350
rect 523880 205630 523908 643486
rect 523972 252550 524000 645050
rect 524052 643680 524104 643686
rect 524052 643622 524104 643628
rect 524064 299470 524092 643622
rect 524156 346390 524184 645390
rect 524328 644156 524380 644162
rect 524328 644098 524380 644104
rect 524236 643884 524288 643890
rect 524236 643826 524288 643832
rect 524248 393310 524276 643826
rect 524340 510610 524368 644098
rect 525064 643476 525116 643482
rect 525064 643418 525116 643424
rect 524510 607064 524566 607073
rect 524510 606999 524566 607008
rect 524524 603265 524552 606999
rect 524510 603256 524566 603265
rect 524510 603191 524566 603200
rect 524328 510604 524380 510610
rect 524328 510546 524380 510552
rect 524236 393304 524288 393310
rect 524236 393246 524288 393252
rect 524144 346384 524196 346390
rect 524144 346326 524196 346332
rect 524052 299464 524104 299470
rect 524052 299406 524104 299412
rect 523960 252544 524012 252550
rect 523960 252486 524012 252492
rect 523868 205624 523920 205630
rect 523868 205566 523920 205572
rect 523776 182164 523828 182170
rect 523776 182106 523828 182112
rect 525076 171086 525104 643418
rect 525154 642832 525210 642841
rect 525154 642767 525210 642776
rect 525168 229090 525196 642767
rect 525260 311846 525288 646546
rect 525352 358766 525380 646682
rect 525432 646672 525484 646678
rect 525432 646614 525484 646620
rect 525444 369850 525472 646614
rect 525536 416770 525564 646886
rect 580262 646847 580318 646856
rect 537484 646808 537536 646814
rect 537484 646750 537536 646756
rect 525616 645652 525668 645658
rect 525616 645594 525668 645600
rect 525628 440230 525656 645594
rect 531964 644224 532016 644230
rect 531964 644166 532016 644172
rect 531976 546446 532004 644166
rect 531964 546440 532016 546446
rect 531964 546382 532016 546388
rect 526442 462632 526498 462641
rect 526442 462567 526498 462576
rect 533986 462632 534042 462641
rect 533986 462567 534042 462576
rect 526456 462097 526484 462567
rect 534000 462482 534028 462567
rect 534170 462496 534226 462505
rect 534000 462454 534170 462482
rect 534170 462431 534226 462440
rect 526442 462088 526498 462097
rect 526442 462023 526498 462032
rect 525616 440224 525668 440230
rect 525616 440166 525668 440172
rect 525524 416764 525576 416770
rect 525524 416706 525576 416712
rect 537496 405686 537524 646750
rect 567844 643748 567896 643754
rect 567844 643690 567896 643696
rect 544382 641880 544438 641889
rect 544382 641815 544438 641824
rect 544396 593366 544424 641815
rect 544384 593360 544436 593366
rect 544384 593302 544436 593308
rect 567856 487150 567884 643690
rect 571982 642016 572038 642025
rect 571982 641951 572038 641960
rect 571996 640286 572024 641951
rect 571984 640280 572036 640286
rect 571984 640222 572036 640228
rect 580172 640280 580224 640286
rect 580172 640222 580224 640228
rect 580184 639441 580212 640222
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 579804 627904 579856 627910
rect 579804 627846 579856 627852
rect 579816 627745 579844 627846
rect 579802 627736 579858 627745
rect 579802 627671 579858 627680
rect 579988 593360 580040 593366
rect 579988 593302 580040 593308
rect 580000 592521 580028 593302
rect 579986 592512 580042 592521
rect 579986 592447 580042 592456
rect 579804 580984 579856 580990
rect 579804 580926 579856 580932
rect 579816 580825 579844 580926
rect 579802 580816 579858 580825
rect 579802 580751 579858 580760
rect 579988 546440 580040 546446
rect 579988 546382 580040 546388
rect 580000 545601 580028 546382
rect 579986 545592 580042 545601
rect 579986 545527 580042 545536
rect 579804 534064 579856 534070
rect 579804 534006 579856 534012
rect 579816 533905 579844 534006
rect 579802 533896 579858 533905
rect 579802 533831 579858 533840
rect 580172 510604 580224 510610
rect 580172 510546 580224 510552
rect 580184 510377 580212 510546
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 567844 487144 567896 487150
rect 567844 487086 567896 487092
rect 579620 487144 579672 487150
rect 579620 487086 579672 487092
rect 579632 486849 579660 487086
rect 579618 486840 579674 486849
rect 579618 486775 579674 486784
rect 549166 462768 549222 462777
rect 549166 462703 549222 462712
rect 549180 462369 549208 462703
rect 560206 462632 560262 462641
rect 560206 462567 560262 462576
rect 560220 462534 560248 462567
rect 553308 462528 553360 462534
rect 553306 462496 553308 462505
rect 560208 462528 560260 462534
rect 553360 462496 553362 462505
rect 560208 462470 560260 462476
rect 553306 462431 553362 462440
rect 549166 462360 549222 462369
rect 549166 462295 549222 462304
rect 579988 452600 580040 452606
rect 579988 452542 580040 452548
rect 580000 451761 580028 452542
rect 579986 451752 580042 451761
rect 579986 451687 580042 451696
rect 579620 440224 579672 440230
rect 579620 440166 579672 440172
rect 579632 439929 579660 440166
rect 579618 439920 579674 439929
rect 579618 439855 579674 439864
rect 580172 416764 580224 416770
rect 580172 416706 580224 416712
rect 580184 416537 580212 416706
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 537484 405680 537536 405686
rect 537484 405622 537536 405628
rect 579988 405680 580040 405686
rect 579988 405622 580040 405628
rect 580000 404841 580028 405622
rect 579986 404832 580042 404841
rect 579986 404767 580042 404776
rect 579620 393304 579672 393310
rect 579620 393246 579672 393252
rect 579632 393009 579660 393246
rect 579618 393000 579674 393009
rect 579618 392935 579674 392944
rect 525432 369844 525484 369850
rect 525432 369786 525484 369792
rect 580172 369844 580224 369850
rect 580172 369786 580224 369792
rect 580184 369617 580212 369786
rect 580170 369608 580226 369617
rect 580170 369543 580226 369552
rect 525340 358760 525392 358766
rect 525340 358702 525392 358708
rect 579988 358760 580040 358766
rect 579988 358702 580040 358708
rect 580000 357921 580028 358702
rect 579986 357912 580042 357921
rect 579986 357847 580042 357856
rect 579620 346384 579672 346390
rect 579620 346326 579672 346332
rect 579632 346089 579660 346326
rect 579618 346080 579674 346089
rect 579618 346015 579674 346024
rect 525248 311840 525300 311846
rect 525248 311782 525300 311788
rect 580172 311840 580224 311846
rect 580172 311782 580224 311788
rect 580184 310865 580212 311782
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 299169 580212 299406
rect 580170 299160 580226 299169
rect 580170 299095 580226 299104
rect 549166 275088 549222 275097
rect 549166 275023 549222 275032
rect 526442 274952 526498 274961
rect 526442 274887 526498 274896
rect 533986 274952 534042 274961
rect 533986 274887 534042 274896
rect 526456 274417 526484 274887
rect 534000 274802 534028 274887
rect 534170 274816 534226 274825
rect 534000 274774 534170 274802
rect 534170 274751 534226 274760
rect 549180 274689 549208 275023
rect 560206 274952 560262 274961
rect 560206 274887 560262 274896
rect 560220 274854 560248 274887
rect 553308 274848 553360 274854
rect 553306 274816 553308 274825
rect 560208 274848 560260 274854
rect 553360 274816 553362 274825
rect 560208 274790 560260 274796
rect 553306 274751 553362 274760
rect 549166 274680 549222 274689
rect 549166 274615 549222 274624
rect 526442 274408 526498 274417
rect 526442 274343 526498 274352
rect 579712 252544 579764 252550
rect 579712 252486 579764 252492
rect 579724 252249 579752 252486
rect 579710 252240 579766 252249
rect 579710 252175 579766 252184
rect 525156 229084 525208 229090
rect 525156 229026 525208 229032
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 580172 205624 580224 205630
rect 580172 205566 580224 205572
rect 580184 205329 580212 205566
rect 580170 205320 580226 205329
rect 580170 205255 580226 205264
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 525064 171080 525116 171086
rect 525064 171022 525116 171028
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 580172 158704 580224 158710
rect 580172 158646 580224 158652
rect 580184 158409 580212 158646
rect 580170 158400 580226 158409
rect 580170 158335 580226 158344
rect 523684 135244 523736 135250
rect 523684 135186 523736 135192
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 522488 111784 522540 111790
rect 522488 111726 522540 111732
rect 579620 111784 579672 111790
rect 579620 111726 579672 111732
rect 579632 111489 579660 111726
rect 579618 111480 579674 111489
rect 579618 111415 579674 111424
rect 549166 87408 549222 87417
rect 549166 87343 549222 87352
rect 533986 87272 534042 87281
rect 533986 87207 534042 87216
rect 534000 87122 534028 87207
rect 534170 87136 534226 87145
rect 534000 87094 534170 87122
rect 534170 87071 534226 87080
rect 549180 87009 549208 87343
rect 560206 87272 560262 87281
rect 560206 87207 560262 87216
rect 560220 87174 560248 87207
rect 553308 87168 553360 87174
rect 553306 87136 553308 87145
rect 560208 87168 560260 87174
rect 553360 87136 553362 87145
rect 560208 87110 560260 87116
rect 553306 87071 553362 87080
rect 549166 87000 549222 87009
rect 549166 86935 549222 86944
rect 522408 66150 522528 66178
rect 522500 64870 522528 66150
rect 522488 64864 522540 64870
rect 522488 64806 522540 64812
rect 580172 64864 580224 64870
rect 580172 64806 580224 64812
rect 580184 64569 580212 64806
rect 580170 64560 580226 64569
rect 580170 64495 580226 64504
rect 524694 44704 524750 44713
rect 524694 44639 524750 44648
rect 522960 42362 522988 44132
rect 522948 42356 523000 42362
rect 522948 42298 523000 42304
rect 522948 41472 523000 41478
rect 522948 41414 523000 41420
rect 522304 17944 522356 17950
rect 522304 17886 522356 17892
rect 522672 6520 522724 6526
rect 522672 6462 522724 6468
rect 520476 3454 521516 3482
rect 520280 2984 520332 2990
rect 520280 2926 520332 2932
rect 520292 480 520320 2926
rect 521488 480 521516 3454
rect 522684 480 522712 6462
rect 522960 3466 522988 41414
rect 524708 40497 524736 44639
rect 543004 42764 543056 42770
rect 543004 42706 543056 42712
rect 541624 42628 541676 42634
rect 541624 42570 541676 42576
rect 531964 42560 532016 42566
rect 531964 42502 532016 42508
rect 530584 42424 530636 42430
rect 530584 42366 530636 42372
rect 528560 42288 528612 42294
rect 528560 42230 528612 42236
rect 527180 42220 527232 42226
rect 527180 42162 527232 42168
rect 524694 40488 524750 40497
rect 524694 40423 524750 40432
rect 526260 6452 526312 6458
rect 526260 6394 526312 6400
rect 522948 3460 523000 3466
rect 522948 3402 523000 3408
rect 523868 3324 523920 3330
rect 523868 3266 523920 3272
rect 523880 480 523908 3266
rect 525064 2916 525116 2922
rect 525064 2858 525116 2864
rect 525076 480 525104 2858
rect 526272 480 526300 6394
rect 527192 3482 527220 42162
rect 528572 3482 528600 42230
rect 529204 41608 529256 41614
rect 529204 41550 529256 41556
rect 527192 3454 527496 3482
rect 528572 3454 528692 3482
rect 527468 480 527496 3454
rect 528664 480 528692 3454
rect 529216 3058 529244 41550
rect 529848 5432 529900 5438
rect 529848 5374 529900 5380
rect 529204 3052 529256 3058
rect 529204 2994 529256 3000
rect 529860 480 529888 5374
rect 530596 3330 530624 42366
rect 530584 3324 530636 3330
rect 530584 3266 530636 3272
rect 531044 3120 531096 3126
rect 531044 3062 531096 3068
rect 531056 480 531084 3062
rect 531976 2990 532004 42502
rect 540244 42152 540296 42158
rect 540244 42094 540296 42100
rect 535460 42084 535512 42090
rect 535460 42026 535512 42032
rect 533344 41880 533396 41886
rect 533344 41822 533396 41828
rect 532240 3188 532292 3194
rect 532240 3130 532292 3136
rect 531964 2984 532016 2990
rect 531964 2926 532016 2932
rect 532252 480 532280 3130
rect 533356 2854 533384 41822
rect 534724 41744 534776 41750
rect 534724 41686 534776 41692
rect 533436 5296 533488 5302
rect 533436 5238 533488 5244
rect 533344 2848 533396 2854
rect 533344 2790 533396 2796
rect 533448 480 533476 5238
rect 534540 3324 534592 3330
rect 534540 3266 534592 3272
rect 534552 480 534580 3266
rect 534736 2922 534764 41686
rect 534724 2916 534776 2922
rect 534724 2858 534776 2864
rect 535472 626 535500 42026
rect 537484 41948 537536 41954
rect 537484 41890 537536 41896
rect 536932 5160 536984 5166
rect 536932 5102 536984 5108
rect 535472 598 535776 626
rect 535748 480 535776 598
rect 536944 480 536972 5102
rect 537496 3058 537524 41890
rect 537576 41812 537628 41818
rect 537576 41754 537628 41760
rect 537588 3126 537616 41754
rect 538864 41676 538916 41682
rect 538864 41618 538916 41624
rect 538876 3126 538904 41618
rect 540256 3398 540284 42094
rect 540886 40760 540942 40769
rect 540886 40695 540942 40704
rect 540900 40361 540928 40695
rect 540886 40352 540942 40361
rect 540886 40287 540942 40296
rect 540520 5364 540572 5370
rect 540520 5306 540572 5312
rect 540244 3392 540296 3398
rect 540244 3334 540296 3340
rect 539324 3256 539376 3262
rect 539324 3198 539376 3204
rect 537576 3120 537628 3126
rect 537576 3062 537628 3068
rect 538864 3120 538916 3126
rect 538864 3062 538916 3068
rect 537484 3052 537536 3058
rect 537484 2994 537536 3000
rect 538128 2984 538180 2990
rect 538128 2926 538180 2932
rect 538140 480 538168 2926
rect 539336 480 539364 3198
rect 540532 480 540560 5306
rect 541636 2990 541664 42570
rect 542912 3392 542964 3398
rect 542912 3334 542964 3340
rect 541716 3256 541768 3262
rect 541716 3198 541768 3204
rect 541624 2984 541676 2990
rect 541624 2926 541676 2932
rect 541728 480 541756 3198
rect 542924 480 542952 3334
rect 543016 2802 543044 42706
rect 544384 42696 544436 42702
rect 544384 42638 544436 42644
rect 544108 5092 544160 5098
rect 544108 5034 544160 5040
rect 543188 2916 543240 2922
rect 543188 2858 543240 2864
rect 543200 2802 543228 2858
rect 543016 2774 543228 2802
rect 544120 480 544148 5034
rect 544396 3398 544424 42638
rect 545764 42492 545816 42498
rect 545764 42434 545816 42440
rect 545776 4078 545804 42434
rect 547236 42356 547288 42362
rect 547236 42298 547288 42304
rect 547144 42016 547196 42022
rect 547144 41958 547196 41964
rect 545304 4072 545356 4078
rect 545304 4014 545356 4020
rect 545764 4072 545816 4078
rect 545764 4014 545816 4020
rect 544384 3392 544436 3398
rect 544384 3334 544436 3340
rect 545316 480 545344 4014
rect 547156 4010 547184 41958
rect 546500 4004 546552 4010
rect 546500 3946 546552 3952
rect 547144 4004 547196 4010
rect 547144 3946 547196 3952
rect 546512 480 546540 3946
rect 547248 3369 547276 42298
rect 565082 40488 565138 40497
rect 565082 40423 565138 40432
rect 560206 40216 560262 40225
rect 560206 40151 560262 40160
rect 560220 39817 560248 40151
rect 565096 40089 565124 40423
rect 572626 40216 572682 40225
rect 572626 40151 572682 40160
rect 565082 40080 565138 40089
rect 572640 40066 572668 40151
rect 572718 40080 572774 40089
rect 572640 40038 572718 40066
rect 565082 40015 565138 40024
rect 572718 40015 572774 40024
rect 560206 39808 560262 39817
rect 560206 39743 560262 39752
rect 580276 29345 580304 646847
rect 580816 645516 580868 645522
rect 580816 645458 580868 645464
rect 580724 645244 580776 645250
rect 580724 645186 580776 645192
rect 580540 643952 580592 643958
rect 580540 643894 580592 643900
rect 580448 643136 580500 643142
rect 580448 643078 580500 643084
rect 580356 641776 580408 641782
rect 580356 641718 580408 641724
rect 580368 76265 580396 641718
rect 580460 123185 580488 643078
rect 580552 217025 580580 643894
rect 580632 643272 580684 643278
rect 580632 643214 580684 643220
rect 580644 263945 580672 643214
rect 580736 322697 580764 645186
rect 580828 498681 580856 645458
rect 580814 498672 580870 498681
rect 580814 498607 580870 498616
rect 580722 322688 580778 322697
rect 580722 322623 580778 322632
rect 580630 263936 580686 263945
rect 580630 263871 580686 263880
rect 580538 217016 580594 217025
rect 580538 216951 580594 216960
rect 580446 123176 580502 123185
rect 580446 123111 580502 123120
rect 580354 76256 580410 76265
rect 580354 76191 580410 76200
rect 580262 29336 580318 29345
rect 580262 29271 580318 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 569040 6384 569092 6390
rect 569040 6326 569092 6332
rect 561956 6248 562008 6254
rect 561956 6190 562008 6196
rect 547696 5228 547748 5234
rect 547696 5170 547748 5176
rect 547234 3360 547290 3369
rect 547234 3295 547290 3304
rect 547708 480 547736 5170
rect 551192 5024 551244 5030
rect 551192 4966 551244 4972
rect 548892 2984 548944 2990
rect 548892 2926 548944 2932
rect 548904 480 548932 2926
rect 550088 2848 550140 2854
rect 550088 2790 550140 2796
rect 550100 480 550128 2790
rect 551204 480 551232 4966
rect 558368 4956 558420 4962
rect 558368 4898 558420 4904
rect 554780 4888 554832 4894
rect 554780 4830 554832 4836
rect 552388 4140 552440 4146
rect 552388 4082 552440 4088
rect 552400 480 552428 4082
rect 553584 3800 553636 3806
rect 553584 3742 553636 3748
rect 553596 480 553624 3742
rect 554792 480 554820 4830
rect 555976 3052 556028 3058
rect 555976 2994 556028 3000
rect 555988 480 556016 2994
rect 557172 2916 557224 2922
rect 557172 2858 557224 2864
rect 557184 480 557212 2858
rect 558380 480 558408 4898
rect 559564 3936 559616 3942
rect 559564 3878 559616 3884
rect 559576 480 559604 3878
rect 560760 3868 560812 3874
rect 560760 3810 560812 3816
rect 560772 480 560800 3810
rect 561968 480 561996 6190
rect 565544 4820 565596 4826
rect 565544 4762 565596 4768
rect 564348 3392 564400 3398
rect 564348 3334 564400 3340
rect 563152 3120 563204 3126
rect 563152 3062 563204 3068
rect 563164 480 563192 3062
rect 564360 480 564388 3334
rect 565556 480 565584 4762
rect 566740 3732 566792 3738
rect 566740 3674 566792 3680
rect 566752 480 566780 3674
rect 567844 3664 567896 3670
rect 567844 3606 567896 3612
rect 567856 480 567884 3606
rect 569052 480 569080 6326
rect 572628 6316 572680 6322
rect 572628 6258 572680 6264
rect 571432 4072 571484 4078
rect 571432 4014 571484 4020
rect 570236 3188 570288 3194
rect 570236 3130 570288 3136
rect 570248 480 570276 3130
rect 571444 480 571472 4014
rect 572640 480 572668 6258
rect 576216 6180 576268 6186
rect 576216 6122 576268 6128
rect 573824 3596 573876 3602
rect 573824 3538 573876 3544
rect 573836 480 573864 3538
rect 575020 3528 575072 3534
rect 575020 3470 575072 3476
rect 575032 480 575060 3470
rect 576228 480 576256 6122
rect 578608 4004 578660 4010
rect 578608 3946 578660 3952
rect 577412 3256 577464 3262
rect 577412 3198 577464 3204
rect 577424 480 577452 3198
rect 578620 480 578648 3946
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 579804 3324 579856 3330
rect 579804 3266 579856 3272
rect 579816 480 579844 3266
rect 581012 480 581040 3402
rect 582194 3360 582250 3369
rect 582194 3295 582250 3304
rect 582208 480 582236 3295
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 8114 700304 8170 700360
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3422 646040 3478 646096
rect 3330 624860 3332 624880
rect 3332 624860 3384 624880
rect 3384 624860 3386 624880
rect 3330 624824 3386 624860
rect 3330 610408 3386 610464
rect 3238 567296 3294 567352
rect 2778 553052 2780 553072
rect 2780 553052 2832 553072
rect 2832 553052 2834 553072
rect 2778 553016 2834 553052
rect 3054 538600 3110 538656
rect 3330 509940 3332 509960
rect 3332 509940 3384 509960
rect 3384 509940 3386 509960
rect 3330 509904 3386 509940
rect 3330 495524 3332 495544
rect 3332 495524 3384 495544
rect 3384 495524 3386 495544
rect 3330 495488 3386 495524
rect 3330 481108 3332 481128
rect 3332 481108 3384 481128
rect 3384 481108 3386 481128
rect 3330 481072 3386 481108
rect 3330 452376 3386 452432
rect 3330 423680 3386 423736
rect 3054 394984 3110 395040
rect 3146 366152 3202 366208
rect 3146 337456 3202 337512
rect 3330 308796 3332 308816
rect 3332 308796 3384 308816
rect 3384 308796 3386 308816
rect 3330 308760 3386 308796
rect 3238 280100 3240 280120
rect 3240 280100 3292 280120
rect 3292 280100 3294 280120
rect 3238 280064 3294 280100
rect 2778 265648 2834 265704
rect 3146 251268 3148 251288
rect 3148 251268 3200 251288
rect 3200 251268 3202 251288
rect 3146 251232 3202 251268
rect 3146 236952 3202 237008
rect 3330 208156 3332 208176
rect 3332 208156 3384 208176
rect 3384 208156 3386 208176
rect 3330 208120 3386 208156
rect 3054 193840 3110 193896
rect 2778 179460 2780 179480
rect 2780 179460 2832 179480
rect 2832 179460 2834 179480
rect 2778 179424 2834 179460
rect 3146 165008 3202 165064
rect 3330 150728 3386 150784
rect 2962 122032 3018 122088
rect 3238 107616 3294 107672
rect 2778 93236 2780 93256
rect 2780 93236 2832 93256
rect 2832 93236 2834 93256
rect 2778 93200 2834 93236
rect 3054 78920 3110 78976
rect 3330 64504 3386 64560
rect 3514 642368 3570 642424
rect 3698 642504 3754 642560
rect 3606 323040 3662 323096
rect 3606 294344 3662 294400
rect 53930 646856 53986 646912
rect 3974 595992 4030 596048
rect 3882 437960 3938 438016
rect 3790 380568 3846 380624
rect 3698 222536 3754 222592
rect 3514 136312 3570 136368
rect 8850 641688 8906 641744
rect 9310 642912 9366 642968
rect 9494 642232 9550 642288
rect 10414 642096 10470 642152
rect 3422 50088 3478 50144
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 3422 8200 3478 8256
rect 3422 7112 3478 7168
rect 66534 646448 66590 646504
rect 62394 646176 62450 646232
rect 112902 646312 112958 646368
rect 163410 646448 163466 646504
rect 188618 646584 188674 646640
rect 201314 646720 201370 646776
rect 125782 643748 125838 643784
rect 125782 643728 125784 643748
rect 125784 643728 125836 643748
rect 125836 643728 125838 643748
rect 339498 700304 339554 700360
rect 365074 686024 365130 686080
rect 364522 685888 364578 685944
rect 580170 697992 580226 698048
rect 494886 686024 494942 686080
rect 494242 685888 494298 685944
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 479154 645904 479210 645960
rect 504454 646040 504510 646096
rect 49974 643320 50030 643376
rect 75274 643320 75330 643376
rect 100482 643320 100538 643376
rect 205454 643320 205510 643376
rect 218426 643320 218482 643376
rect 369398 643320 369454 643376
rect 390558 643320 390614 643376
rect 394790 643320 394846 643376
rect 428462 643320 428518 643376
rect 453670 643320 453726 643376
rect 516690 643320 516746 643376
rect 520922 643320 520978 643376
rect 522118 616800 522174 616856
rect 522118 610136 522174 610192
rect 31482 9696 31538 9752
rect 31666 9696 31722 9752
rect 44086 42064 44142 42120
rect 73434 38664 73490 38720
rect 74354 38800 74410 38856
rect 79230 42064 79286 42120
rect 100666 42064 100722 42120
rect 108762 9696 108818 9752
rect 108946 9696 109002 9752
rect 118146 29144 118202 29200
rect 117410 29008 117466 29064
rect 121090 27784 121146 27840
rect 120170 27648 120226 27704
rect 126242 42064 126298 42120
rect 441434 3052 441490 3088
rect 441434 3032 441436 3052
rect 441436 3032 441488 3052
rect 441488 3032 441490 3052
rect 442906 3304 442962 3360
rect 447046 3032 447102 3088
rect 484582 3304 484638 3360
rect 523682 642640 523738 642696
rect 524510 607008 524566 607064
rect 524510 603200 524566 603256
rect 525154 642776 525210 642832
rect 580262 646856 580318 646912
rect 526442 462576 526498 462632
rect 533986 462576 534042 462632
rect 534170 462440 534226 462496
rect 526442 462032 526498 462088
rect 544382 641824 544438 641880
rect 571982 641960 572038 642016
rect 580170 639376 580226 639432
rect 579802 627680 579858 627736
rect 579986 592456 580042 592512
rect 579802 580760 579858 580816
rect 579986 545536 580042 545592
rect 579802 533840 579858 533896
rect 580170 510312 580226 510368
rect 579618 486784 579674 486840
rect 549166 462712 549222 462768
rect 560206 462576 560262 462632
rect 553306 462476 553308 462496
rect 553308 462476 553360 462496
rect 553360 462476 553362 462496
rect 553306 462440 553362 462476
rect 549166 462304 549222 462360
rect 579986 451696 580042 451752
rect 579618 439864 579674 439920
rect 580170 416472 580226 416528
rect 579986 404776 580042 404832
rect 579618 392944 579674 393000
rect 580170 369552 580226 369608
rect 579986 357856 580042 357912
rect 579618 346024 579674 346080
rect 580170 310800 580226 310856
rect 580170 299104 580226 299160
rect 549166 275032 549222 275088
rect 526442 274896 526498 274952
rect 533986 274896 534042 274952
rect 534170 274760 534226 274816
rect 560206 274896 560262 274952
rect 553306 274796 553308 274816
rect 553308 274796 553360 274816
rect 553360 274796 553362 274816
rect 553306 274760 553362 274796
rect 549166 274624 549222 274680
rect 526442 274352 526498 274408
rect 579710 252184 579766 252240
rect 580170 228792 580226 228848
rect 580170 205264 580226 205320
rect 580170 181872 580226 181928
rect 580170 170040 580226 170096
rect 580170 158344 580226 158400
rect 580170 134816 580226 134872
rect 579618 111424 579674 111480
rect 549166 87352 549222 87408
rect 533986 87216 534042 87272
rect 534170 87080 534226 87136
rect 560206 87216 560262 87272
rect 553306 87116 553308 87136
rect 553308 87116 553360 87136
rect 553360 87116 553362 87136
rect 553306 87080 553362 87116
rect 549166 86944 549222 87000
rect 580170 64504 580226 64560
rect 524694 44648 524750 44704
rect 524694 40432 524750 40488
rect 540886 40704 540942 40760
rect 540886 40296 540942 40352
rect 565082 40432 565138 40488
rect 560206 40160 560262 40216
rect 572626 40160 572682 40216
rect 565082 40024 565138 40080
rect 572718 40024 572774 40080
rect 560206 39752 560262 39808
rect 580814 498616 580870 498672
rect 580722 322632 580778 322688
rect 580630 263880 580686 263936
rect 580538 216960 580594 217016
rect 580446 123120 580502 123176
rect 580354 76200 580410 76256
rect 580262 29280 580318 29336
rect 579802 17584 579858 17640
rect 547234 3304 547290 3360
rect 582194 3304 582250 3360
<< metal3 >>
rect 8109 700362 8175 700365
rect 339493 700362 339559 700365
rect 8109 700360 339559 700362
rect 8109 700304 8114 700360
rect 8170 700304 339498 700360
rect 339554 700304 339559 700360
rect 8109 700302 339559 700304
rect 8109 700299 8175 700302
rect 339493 700299 339559 700302
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 365069 686082 365135 686085
rect 494881 686082 494947 686085
rect 364382 686080 365135 686082
rect 364382 686024 365074 686080
rect 365130 686024 365135 686080
rect 364382 686022 365135 686024
rect 364382 685946 364442 686022
rect 365069 686019 365135 686022
rect 494102 686080 494947 686082
rect 494102 686024 494886 686080
rect 494942 686024 494947 686080
rect 494102 686022 494947 686024
rect 364517 685946 364583 685949
rect 364382 685944 364583 685946
rect 364382 685888 364522 685944
rect 364578 685888 364583 685944
rect 364382 685886 364583 685888
rect 494102 685946 494162 686022
rect 494881 686019 494947 686022
rect 494237 685946 494303 685949
rect 494102 685944 494303 685946
rect 494102 685888 494242 685944
rect 494298 685888 494303 685944
rect 494102 685886 494303 685888
rect 364517 685883 364583 685886
rect 494237 685883 494303 685886
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 53925 646914 53991 646917
rect 580257 646914 580323 646917
rect 53925 646912 580323 646914
rect 53925 646856 53930 646912
rect 53986 646856 580262 646912
rect 580318 646856 580323 646912
rect 53925 646854 580323 646856
rect 53925 646851 53991 646854
rect 580257 646851 580323 646854
rect 201309 646778 201375 646781
rect 521510 646778 521516 646780
rect 201309 646776 521516 646778
rect 201309 646720 201314 646776
rect 201370 646720 521516 646776
rect 201309 646718 521516 646720
rect 201309 646715 201375 646718
rect 521510 646716 521516 646718
rect 521580 646716 521586 646780
rect 188613 646642 188679 646645
rect 520590 646642 520596 646644
rect 188613 646640 520596 646642
rect 188613 646584 188618 646640
rect 188674 646584 520596 646640
rect 188613 646582 520596 646584
rect 188613 646579 188679 646582
rect 520590 646580 520596 646582
rect 520660 646580 520666 646644
rect 66529 646506 66595 646509
rect 125726 646506 125732 646508
rect 66529 646504 125732 646506
rect 66529 646448 66534 646504
rect 66590 646448 125732 646504
rect 66529 646446 125732 646448
rect 66529 646443 66595 646446
rect 125726 646444 125732 646446
rect 125796 646444 125802 646508
rect 163405 646506 163471 646509
rect 521142 646506 521148 646508
rect 163405 646504 521148 646506
rect 163405 646448 163410 646504
rect 163466 646448 521148 646504
rect 163405 646446 521148 646448
rect 163405 646443 163471 646446
rect 521142 646444 521148 646446
rect 521212 646444 521218 646508
rect 112897 646370 112963 646373
rect 520958 646370 520964 646372
rect 112897 646368 520964 646370
rect 112897 646312 112902 646368
rect 112958 646312 520964 646368
rect 112897 646310 520964 646312
rect 112897 646307 112963 646310
rect 520958 646308 520964 646310
rect 521028 646308 521034 646372
rect 62389 646234 62455 646237
rect 520774 646234 520780 646236
rect 62389 646232 520780 646234
rect 62389 646176 62394 646232
rect 62450 646176 520780 646232
rect 62389 646174 520780 646176
rect 62389 646171 62455 646174
rect 520774 646172 520780 646174
rect 520844 646172 520850 646236
rect 3417 646098 3483 646101
rect 504449 646098 504515 646101
rect 3417 646096 504515 646098
rect 3417 646040 3422 646096
rect 3478 646040 504454 646096
rect 504510 646040 504515 646096
rect 3417 646038 504515 646040
rect 3417 646035 3483 646038
rect 504449 646035 504515 646038
rect 471278 645900 471284 645964
rect 471348 645962 471354 645964
rect 479149 645962 479215 645965
rect 471348 645960 479215 645962
rect 471348 645904 479154 645960
rect 479210 645904 479215 645960
rect 471348 645902 479215 645904
rect 471348 645900 471354 645902
rect 479149 645899 479215 645902
rect 125777 643788 125843 643789
rect 125726 643786 125732 643788
rect 125686 643726 125732 643786
rect 125796 643784 125843 643788
rect 125838 643728 125843 643784
rect 125726 643724 125732 643726
rect 125796 643724 125843 643728
rect 125777 643723 125843 643724
rect 49969 643378 50035 643381
rect 75269 643380 75335 643381
rect 100477 643380 100543 643381
rect 205449 643380 205515 643381
rect 50838 643378 50844 643380
rect 49969 643376 50844 643378
rect 49969 643320 49974 643376
rect 50030 643320 50844 643376
rect 49969 643318 50844 643320
rect 49969 643315 50035 643318
rect 50838 643316 50844 643318
rect 50908 643316 50914 643380
rect 75269 643376 75316 643380
rect 75380 643378 75386 643380
rect 75269 643320 75274 643376
rect 75269 643316 75316 643320
rect 75380 643318 75426 643378
rect 100477 643376 100524 643380
rect 100588 643378 100594 643380
rect 205398 643378 205404 643380
rect 100477 643320 100482 643376
rect 75380 643316 75386 643318
rect 100477 643316 100524 643320
rect 100588 643318 100634 643378
rect 205358 643318 205404 643378
rect 205468 643376 205515 643380
rect 205510 643320 205515 643376
rect 100588 643316 100594 643318
rect 205398 643316 205404 643318
rect 205468 643316 205515 643320
rect 75269 643315 75335 643316
rect 100477 643315 100543 643316
rect 205449 643315 205515 643316
rect 218421 643380 218487 643381
rect 369393 643380 369459 643381
rect 390553 643380 390619 643381
rect 394785 643380 394851 643381
rect 218421 643376 218468 643380
rect 218532 643378 218538 643380
rect 369342 643378 369348 643380
rect 218421 643320 218426 643376
rect 218421 643316 218468 643320
rect 218532 643318 218578 643378
rect 369302 643318 369348 643378
rect 369412 643376 369459 643380
rect 390502 643378 390508 643380
rect 369454 643320 369459 643376
rect 218532 643316 218538 643318
rect 369342 643316 369348 643318
rect 369412 643316 369459 643320
rect 390462 643318 390508 643378
rect 390572 643376 390619 643380
rect 394734 643378 394740 643380
rect 390614 643320 390619 643376
rect 390502 643316 390508 643318
rect 390572 643316 390619 643320
rect 394694 643318 394740 643378
rect 394804 643376 394851 643380
rect 428457 643378 428523 643381
rect 453665 643380 453731 643381
rect 453614 643378 453620 643380
rect 394846 643320 394851 643376
rect 394734 643316 394740 643318
rect 394804 643316 394851 643320
rect 218421 643315 218487 643316
rect 369393 643315 369459 643316
rect 390553 643315 390619 643316
rect 394785 643315 394851 643316
rect 428414 643376 428523 643378
rect 428414 643320 428462 643376
rect 428518 643320 428523 643376
rect 428414 643315 428523 643320
rect 453574 643318 453620 643378
rect 453684 643376 453731 643380
rect 453726 643320 453731 643376
rect 453614 643316 453620 643318
rect 453684 643316 453731 643320
rect 516358 643316 516364 643380
rect 516428 643378 516434 643380
rect 516685 643378 516751 643381
rect 516428 643376 516751 643378
rect 516428 643320 516690 643376
rect 516746 643320 516751 643376
rect 516428 643318 516751 643320
rect 516428 643316 516434 643318
rect 453665 643315 453731 643316
rect 516685 643315 516751 643318
rect 518014 643316 518020 643380
rect 518084 643378 518090 643380
rect 520917 643378 520983 643381
rect 518084 643376 520983 643378
rect 518084 643320 520922 643376
rect 520978 643320 520983 643376
rect 518084 643318 520983 643320
rect 518084 643316 518090 643318
rect 520917 643315 520983 643318
rect 240910 643044 240916 643108
rect 240980 643106 240986 643108
rect 253790 643106 253796 643108
rect 240980 643046 253796 643106
rect 240980 643044 240986 643046
rect 253790 643044 253796 643046
rect 253860 643044 253866 643108
rect 264462 643044 264468 643108
rect 264532 643106 264538 643108
rect 273110 643106 273116 643108
rect 264532 643046 273116 643106
rect 264532 643044 264538 643046
rect 273110 643044 273116 643046
rect 273180 643044 273186 643108
rect 282862 643044 282868 643108
rect 282932 643106 282938 643108
rect 311750 643106 311756 643108
rect 282932 643046 311756 643106
rect 282932 643044 282938 643046
rect 311750 643044 311756 643046
rect 311820 643044 311826 643108
rect 335302 643044 335308 643108
rect 335372 643106 335378 643108
rect 349654 643106 349660 643108
rect 335372 643046 349660 643106
rect 335372 643044 335378 643046
rect 349654 643044 349660 643046
rect 349724 643044 349730 643108
rect 350758 643044 350764 643108
rect 350828 643106 350834 643108
rect 369710 643106 369716 643108
rect 350828 643046 369716 643106
rect 350828 643044 350834 643046
rect 369710 643044 369716 643046
rect 369780 643044 369786 643108
rect 9305 642970 9371 642973
rect 428414 642970 428474 643315
rect 9305 642968 428474 642970
rect 9305 642912 9310 642968
rect 9366 642912 428474 642968
rect 9305 642910 428474 642912
rect 9305 642907 9371 642910
rect 100518 642772 100524 642836
rect 100588 642834 100594 642836
rect 525149 642834 525215 642837
rect 100588 642832 525215 642834
rect 100588 642776 525154 642832
rect 525210 642776 525215 642832
rect 100588 642774 525215 642776
rect 100588 642772 100594 642774
rect 525149 642771 525215 642774
rect 75310 642636 75316 642700
rect 75380 642698 75386 642700
rect 523677 642698 523743 642701
rect 75380 642696 523743 642698
rect 75380 642640 523682 642696
rect 523738 642640 523743 642696
rect 75380 642638 523743 642640
rect 75380 642636 75386 642638
rect 523677 642635 523743 642638
rect 3693 642562 3759 642565
rect 453614 642562 453620 642564
rect 3693 642560 453620 642562
rect 3693 642504 3698 642560
rect 3754 642504 453620 642560
rect 3693 642502 453620 642504
rect 3693 642499 3759 642502
rect 453614 642500 453620 642502
rect 453684 642500 453690 642564
rect 3509 642426 3575 642429
rect 471278 642426 471284 642428
rect 3509 642424 471284 642426
rect 3509 642368 3514 642424
rect 3570 642368 471284 642424
rect 3509 642366 471284 642368
rect 3509 642363 3575 642366
rect 471278 642364 471284 642366
rect 471348 642364 471354 642428
rect 9489 642290 9555 642293
rect 390502 642290 390508 642292
rect 9489 642288 390508 642290
rect 9489 642232 9494 642288
rect 9550 642232 390508 642288
rect 9489 642230 390508 642232
rect 9489 642227 9555 642230
rect 390502 642228 390508 642230
rect 390572 642228 390578 642292
rect 10409 642154 10475 642157
rect 369342 642154 369348 642156
rect 10409 642152 369348 642154
rect 10409 642096 10414 642152
rect 10470 642096 369348 642152
rect 10409 642094 369348 642096
rect 10409 642091 10475 642094
rect 369342 642092 369348 642094
rect 369412 642092 369418 642156
rect 379646 642092 379652 642156
rect 379716 642154 379722 642156
rect 391238 642154 391244 642156
rect 379716 642094 391244 642154
rect 379716 642092 379722 642094
rect 391238 642092 391244 642094
rect 391308 642092 391314 642156
rect 218462 641956 218468 642020
rect 218532 642018 218538 642020
rect 571977 642018 572043 642021
rect 218532 642016 572043 642018
rect 218532 641960 571982 642016
rect 572038 641960 572043 642016
rect 218532 641958 572043 641960
rect 218532 641956 218538 641958
rect 571977 641955 572043 641958
rect 75862 641820 75868 641884
rect 75932 641882 75938 641884
rect 85430 641882 85436 641884
rect 75932 641822 85436 641882
rect 75932 641820 75938 641822
rect 85430 641820 85436 641822
rect 85500 641820 85506 641884
rect 95182 641820 95188 641884
rect 95252 641882 95258 641884
rect 104750 641882 104756 641884
rect 95252 641822 104756 641882
rect 95252 641820 95258 641822
rect 104750 641820 104756 641822
rect 104820 641820 104826 641884
rect 153142 641820 153148 641884
rect 153212 641882 153218 641884
rect 162526 641882 162532 641884
rect 153212 641822 162532 641882
rect 153212 641820 153218 641822
rect 162526 641820 162532 641822
rect 162596 641820 162602 641884
rect 164182 641820 164188 641884
rect 164252 641882 164258 641884
rect 178718 641882 178724 641884
rect 164252 641822 178724 641882
rect 164252 641820 164258 641822
rect 178718 641820 178724 641822
rect 178788 641820 178794 641884
rect 186262 641820 186268 641884
rect 186332 641882 186338 641884
rect 195830 641882 195836 641884
rect 186332 641822 195836 641882
rect 186332 641820 186338 641822
rect 195830 641820 195836 641822
rect 195900 641820 195906 641884
rect 205398 641820 205404 641884
rect 205468 641882 205474 641884
rect 544377 641882 544443 641885
rect 205468 641880 544443 641882
rect 205468 641824 544382 641880
rect 544438 641824 544443 641880
rect 205468 641822 544443 641824
rect 205468 641820 205474 641822
rect 544377 641819 544443 641822
rect 8845 641746 8911 641749
rect 394734 641746 394740 641748
rect 8845 641744 394740 641746
rect 8845 641688 8850 641744
rect 8906 641688 394740 641744
rect 8845 641686 394740 641688
rect 8845 641683 8911 641686
rect 394734 641684 394740 641686
rect 394804 641684 394810 641748
rect 398782 641684 398788 641748
rect 398852 641746 398858 641748
rect 410558 641746 410564 641748
rect 398852 641686 410564 641746
rect 398852 641684 398858 641686
rect 410558 641684 410564 641686
rect 410628 641684 410634 641748
rect 418102 641684 418108 641748
rect 418172 641746 418178 641748
rect 427670 641746 427676 641748
rect 418172 641686 427676 641746
rect 418172 641684 418178 641686
rect 427670 641684 427676 641686
rect 427740 641684 427746 641748
rect 442942 641684 442948 641748
rect 443012 641746 443018 641748
rect 452510 641746 452516 641748
rect 443012 641686 452516 641746
rect 443012 641684 443018 641686
rect 452510 641684 452516 641686
rect 452580 641684 452586 641748
rect 462446 641684 462452 641748
rect 462516 641746 462522 641748
rect 471830 641746 471836 641748
rect 462516 641686 471836 641746
rect 462516 641684 462522 641686
rect 471830 641684 471836 641686
rect 471900 641684 471906 641748
rect 481582 641684 481588 641748
rect 481652 641746 481658 641748
rect 491150 641746 491156 641748
rect 481652 641686 491156 641746
rect 481652 641684 481658 641686
rect 491150 641684 491156 641686
rect 491220 641684 491226 641748
rect 500902 641684 500908 641748
rect 500972 641746 500978 641748
rect 519486 641746 519492 641748
rect 500972 641686 519492 641746
rect 500972 641684 500978 641686
rect 519486 641684 519492 641686
rect 519556 641684 519562 641748
rect 520590 641684 520596 641748
rect 520660 641746 520666 641748
rect 521326 641746 521332 641748
rect 520660 641686 521332 641746
rect 520660 641684 520666 641686
rect 521326 641684 521332 641686
rect 521396 641684 521402 641748
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 521510 636788 521516 636852
rect 521580 636788 521586 636852
rect 521518 636580 521578 636788
rect 521510 636516 521516 636580
rect 521580 636516 521586 636580
rect 521510 628764 521516 628828
rect 521580 628764 521586 628828
rect 521518 628012 521578 628764
rect 521510 627948 521516 628012
rect 521580 627948 521586 628012
rect 579797 627738 579863 627741
rect 583520 627738 584960 627828
rect 579797 627736 584960 627738
rect 579797 627680 579802 627736
rect 579858 627680 584960 627736
rect 579797 627678 584960 627680
rect 579797 627675 579863 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3325 624882 3391 624885
rect -960 624880 3391 624882
rect -960 624824 3330 624880
rect 3386 624824 3391 624880
rect -960 624822 3391 624824
rect -960 624732 480 624822
rect 3325 624819 3391 624822
rect 521510 616796 521516 616860
rect 521580 616858 521586 616860
rect 522113 616858 522179 616861
rect 521580 616856 522179 616858
rect 521580 616800 522118 616856
rect 522174 616800 522179 616856
rect 521580 616798 522179 616800
rect 521580 616796 521586 616798
rect 522113 616795 522179 616798
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3325 610466 3391 610469
rect -960 610464 3391 610466
rect -960 610408 3330 610464
rect 3386 610408 3391 610464
rect -960 610406 3391 610408
rect -960 610316 480 610406
rect 3325 610403 3391 610406
rect 521510 610132 521516 610196
rect 521580 610194 521586 610196
rect 522113 610194 522179 610197
rect 521580 610192 522179 610194
rect 521580 610136 522118 610192
rect 522174 610136 522179 610192
rect 521580 610134 522179 610136
rect 521580 610132 521586 610134
rect 522113 610131 522179 610134
rect 521510 607004 521516 607068
rect 521580 607066 521586 607068
rect 524505 607066 524571 607069
rect 521580 607064 524571 607066
rect 521580 607008 524510 607064
rect 524566 607008 524571 607064
rect 521580 607006 524571 607008
rect 521580 607004 521586 607006
rect 524505 607003 524571 607006
rect 583520 604210 584960 604300
rect 583342 604150 584960 604210
rect 538262 603334 547890 603394
rect 524505 603258 524571 603261
rect 524505 603256 538138 603258
rect 524505 603200 524510 603256
rect 524566 603200 538138 603256
rect 524505 603198 538138 603200
rect 524505 603195 524571 603198
rect 538078 603122 538138 603198
rect 538262 603122 538322 603334
rect 547830 603258 547890 603334
rect 557582 603334 567210 603394
rect 547830 603198 557458 603258
rect 538078 603062 538322 603122
rect 557398 603122 557458 603198
rect 557582 603122 557642 603334
rect 567150 603258 567210 603334
rect 567150 603198 576778 603258
rect 557398 603062 557642 603122
rect 576718 603122 576778 603198
rect 583342 603122 583402 604150
rect 583520 604060 584960 604150
rect 576718 603062 583402 603122
rect -960 596050 480 596140
rect 3969 596050 4035 596053
rect -960 596048 4035 596050
rect -960 595992 3974 596048
rect 4030 595992 4035 596048
rect -960 595990 4035 595992
rect -960 595900 480 595990
rect 3969 595987 4035 595990
rect 579981 592514 580047 592517
rect 583520 592514 584960 592604
rect 579981 592512 584960 592514
rect 579981 592456 579986 592512
rect 580042 592456 584960 592512
rect 579981 592454 584960 592456
rect 579981 592451 580047 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 579797 580818 579863 580821
rect 583520 580818 584960 580908
rect 579797 580816 584960 580818
rect 579797 580760 579802 580816
rect 579858 580760 584960 580816
rect 579797 580758 584960 580760
rect 579797 580755 579863 580758
rect 583520 580668 584960 580758
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3233 567354 3299 567357
rect -960 567352 3299 567354
rect -960 567296 3238 567352
rect 3294 567296 3299 567352
rect -960 567294 3299 567296
rect -960 567204 480 567294
rect 3233 567291 3299 567294
rect 521878 563212 521884 563276
rect 521948 563212 521954 563276
rect 521510 562668 521516 562732
rect 521580 562730 521586 562732
rect 521886 562730 521946 563212
rect 521580 562670 521946 562730
rect 521580 562668 521586 562670
rect 583520 557290 584960 557380
rect 583342 557230 584960 557290
rect 521510 556548 521516 556612
rect 521580 556548 521586 556612
rect 521518 556474 521578 556548
rect 521518 556414 528570 556474
rect 528510 556338 528570 556414
rect 538262 556414 547890 556474
rect 528510 556278 538138 556338
rect 538078 556202 538138 556278
rect 538262 556202 538322 556414
rect 547830 556338 547890 556414
rect 557582 556414 567210 556474
rect 547830 556278 557458 556338
rect 538078 556142 538322 556202
rect 557398 556202 557458 556278
rect 557582 556202 557642 556414
rect 567150 556338 567210 556414
rect 567150 556278 576778 556338
rect 557398 556142 557642 556202
rect 576718 556202 576778 556278
rect 583342 556202 583402 557230
rect 583520 557140 584960 557230
rect 576718 556142 583402 556202
rect -960 553074 480 553164
rect 2773 553074 2839 553077
rect -960 553072 2839 553074
rect -960 553016 2778 553072
rect 2834 553016 2839 553072
rect -960 553014 2839 553016
rect -960 552924 480 553014
rect 2773 553011 2839 553014
rect 579981 545594 580047 545597
rect 583520 545594 584960 545684
rect 579981 545592 584960 545594
rect 579981 545536 579986 545592
rect 580042 545536 584960 545592
rect 579981 545534 584960 545536
rect 579981 545531 580047 545534
rect 583520 545444 584960 545534
rect -960 538658 480 538748
rect 3049 538658 3115 538661
rect -960 538656 3115 538658
rect -960 538600 3054 538656
rect 3110 538600 3115 538656
rect -960 538598 3115 538600
rect -960 538508 480 538598
rect 3049 538595 3115 538598
rect 579797 533898 579863 533901
rect 583520 533898 584960 533988
rect 579797 533896 584960 533898
rect 579797 533840 579802 533896
rect 579858 533840 584960 533896
rect 579797 533838 584960 533840
rect 579797 533835 579863 533838
rect 583520 533748 584960 533838
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3325 509962 3391 509965
rect -960 509960 3391 509962
rect -960 509904 3330 509960
rect 3386 509904 3391 509960
rect -960 509902 3391 509904
rect -960 509812 480 509902
rect 3325 509899 3391 509902
rect 580809 498674 580875 498677
rect 583520 498674 584960 498764
rect 580809 498672 584960 498674
rect 580809 498616 580814 498672
rect 580870 498616 584960 498672
rect 580809 498614 584960 498616
rect 580809 498611 580875 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3325 495546 3391 495549
rect -960 495544 3391 495546
rect -960 495488 3330 495544
rect 3386 495488 3391 495544
rect -960 495486 3391 495488
rect -960 495396 480 495486
rect 3325 495483 3391 495486
rect 579613 486842 579679 486845
rect 583520 486842 584960 486932
rect 579613 486840 584960 486842
rect 579613 486784 579618 486840
rect 579674 486784 584960 486840
rect 579613 486782 584960 486784
rect 579613 486779 579679 486782
rect 583520 486692 584960 486782
rect -960 481130 480 481220
rect 3325 481130 3391 481133
rect -960 481128 3391 481130
rect -960 481072 3330 481128
rect 3386 481072 3391 481128
rect -960 481070 3391 481072
rect -960 480980 480 481070
rect 3325 481067 3391 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 583520 463450 584960 463540
rect 583342 463390 584960 463450
rect 539542 462708 539548 462772
rect 539612 462770 539618 462772
rect 549161 462770 549227 462773
rect 539612 462768 549227 462770
rect 539612 462712 549166 462768
rect 549222 462712 549227 462768
rect 539612 462710 549227 462712
rect 539612 462708 539618 462710
rect 549161 462707 549227 462710
rect 526437 462634 526503 462637
rect 533981 462634 534047 462637
rect 526437 462632 534047 462634
rect 526437 462576 526442 462632
rect 526498 462576 533986 462632
rect 534042 462576 534047 462632
rect 526437 462574 534047 462576
rect 526437 462571 526503 462574
rect 533981 462571 534047 462574
rect 560201 462634 560267 462637
rect 560201 462632 567210 462634
rect 560201 462576 560206 462632
rect 560262 462576 567210 462632
rect 560201 462574 567210 462576
rect 560201 462571 560267 462574
rect 534165 462498 534231 462501
rect 539542 462498 539548 462500
rect 534165 462496 539548 462498
rect 534165 462440 534170 462496
rect 534226 462440 539548 462496
rect 534165 462438 539548 462440
rect 534165 462435 534231 462438
rect 539542 462436 539548 462438
rect 539612 462436 539618 462500
rect 553301 462498 553367 462501
rect 550590 462496 553367 462498
rect 550590 462440 553306 462496
rect 553362 462440 553367 462496
rect 550590 462438 553367 462440
rect 567150 462498 567210 462574
rect 583342 462498 583402 463390
rect 583520 463300 584960 463390
rect 567150 462438 576778 462498
rect 521510 462300 521516 462364
rect 521580 462362 521586 462364
rect 549161 462362 549227 462365
rect 550590 462362 550650 462438
rect 553301 462435 553367 462438
rect 521580 462302 521762 462362
rect 521580 462300 521586 462302
rect 521702 462090 521762 462302
rect 549161 462360 550650 462362
rect 549161 462304 549166 462360
rect 549222 462304 550650 462360
rect 549161 462302 550650 462304
rect 576718 462362 576778 462438
rect 576902 462438 583402 462498
rect 576902 462362 576962 462438
rect 576718 462302 576962 462362
rect 549161 462299 549227 462302
rect 526437 462090 526503 462093
rect 521702 462088 526503 462090
rect 521702 462032 526442 462088
rect 526498 462032 526503 462088
rect 521702 462030 526503 462032
rect 526437 462027 526503 462030
rect -960 452434 480 452524
rect 3325 452434 3391 452437
rect -960 452432 3391 452434
rect -960 452376 3330 452432
rect 3386 452376 3391 452432
rect -960 452374 3391 452376
rect -960 452284 480 452374
rect 3325 452371 3391 452374
rect 579981 451754 580047 451757
rect 583520 451754 584960 451844
rect 579981 451752 584960 451754
rect 579981 451696 579986 451752
rect 580042 451696 584960 451752
rect 579981 451694 584960 451696
rect 579981 451691 580047 451694
rect 583520 451604 584960 451694
rect 579613 439922 579679 439925
rect 583520 439922 584960 440012
rect 579613 439920 584960 439922
rect 579613 439864 579618 439920
rect 579674 439864 584960 439920
rect 579613 439862 584960 439864
rect 579613 439859 579679 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3877 438018 3943 438021
rect -960 438016 3943 438018
rect -960 437960 3882 438016
rect 3938 437960 3943 438016
rect -960 437958 3943 437960
rect -960 437868 480 437958
rect 3877 437955 3943 437958
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3325 423738 3391 423741
rect -960 423736 3391 423738
rect -960 423680 3330 423736
rect 3386 423680 3391 423736
rect -960 423678 3391 423680
rect -960 423588 480 423678
rect 3325 423675 3391 423678
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 579981 404834 580047 404837
rect 583520 404834 584960 404924
rect 579981 404832 584960 404834
rect 579981 404776 579986 404832
rect 580042 404776 584960 404832
rect 579981 404774 584960 404776
rect 579981 404771 580047 404774
rect 583520 404684 584960 404774
rect -960 395042 480 395132
rect 3049 395042 3115 395045
rect -960 395040 3115 395042
rect -960 394984 3054 395040
rect 3110 394984 3115 395040
rect -960 394982 3115 394984
rect -960 394892 480 394982
rect 3049 394979 3115 394982
rect 579613 393002 579679 393005
rect 583520 393002 584960 393092
rect 579613 393000 584960 393002
rect 579613 392944 579618 393000
rect 579674 392944 584960 393000
rect 579613 392942 584960 392944
rect 579613 392939 579679 392942
rect 583520 392852 584960 392942
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3785 380626 3851 380629
rect -960 380624 3851 380626
rect -960 380568 3790 380624
rect 3846 380568 3851 380624
rect -960 380566 3851 380568
rect -960 380476 480 380566
rect 3785 380563 3851 380566
rect 580165 369610 580231 369613
rect 583520 369610 584960 369700
rect 580165 369608 584960 369610
rect 580165 369552 580170 369608
rect 580226 369552 584960 369608
rect 580165 369550 584960 369552
rect 580165 369547 580231 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 3141 366210 3207 366213
rect -960 366208 3207 366210
rect -960 366152 3146 366208
rect 3202 366152 3207 366208
rect -960 366150 3207 366152
rect -960 366060 480 366150
rect 3141 366147 3207 366150
rect 579981 357914 580047 357917
rect 583520 357914 584960 358004
rect 579981 357912 584960 357914
rect 579981 357856 579986 357912
rect 580042 357856 584960 357912
rect 579981 357854 584960 357856
rect 579981 357851 580047 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 579613 346082 579679 346085
rect 583520 346082 584960 346172
rect 579613 346080 584960 346082
rect 579613 346024 579618 346080
rect 579674 346024 584960 346080
rect 579613 346022 584960 346024
rect 579613 346019 579679 346022
rect 583520 345932 584960 346022
rect -960 337514 480 337604
rect 3141 337514 3207 337517
rect -960 337512 3207 337514
rect -960 337456 3146 337512
rect 3202 337456 3207 337512
rect -960 337454 3207 337456
rect -960 337364 480 337454
rect 3141 337451 3207 337454
rect 583520 334236 584960 334476
rect -960 323098 480 323188
rect 3601 323098 3667 323101
rect -960 323096 3667 323098
rect -960 323040 3606 323096
rect 3662 323040 3667 323096
rect -960 323038 3667 323040
rect -960 322948 480 323038
rect 3601 323035 3667 323038
rect 580717 322690 580783 322693
rect 583520 322690 584960 322780
rect 580717 322688 584960 322690
rect 580717 322632 580722 322688
rect 580778 322632 584960 322688
rect 580717 322630 584960 322632
rect 580717 322627 580783 322630
rect 583520 322540 584960 322630
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 580165 299162 580231 299165
rect 583520 299162 584960 299252
rect 580165 299160 584960 299162
rect 580165 299104 580170 299160
rect 580226 299104 584960 299160
rect 580165 299102 584960 299104
rect 580165 299099 580231 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 3601 294402 3667 294405
rect -960 294400 3667 294402
rect -960 294344 3606 294400
rect 3662 294344 3667 294400
rect -960 294342 3667 294344
rect -960 294252 480 294342
rect 3601 294339 3667 294342
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 3233 280122 3299 280125
rect -960 280120 3299 280122
rect -960 280064 3238 280120
rect 3294 280064 3299 280120
rect -960 280062 3299 280064
rect -960 279972 480 280062
rect 3233 280059 3299 280062
rect 583520 275770 584960 275860
rect 583342 275710 584960 275770
rect 539542 275028 539548 275092
rect 539612 275090 539618 275092
rect 549161 275090 549227 275093
rect 539612 275088 549227 275090
rect 539612 275032 549166 275088
rect 549222 275032 549227 275088
rect 539612 275030 549227 275032
rect 539612 275028 539618 275030
rect 549161 275027 549227 275030
rect 526437 274954 526503 274957
rect 533981 274954 534047 274957
rect 526437 274952 534047 274954
rect 526437 274896 526442 274952
rect 526498 274896 533986 274952
rect 534042 274896 534047 274952
rect 526437 274894 534047 274896
rect 526437 274891 526503 274894
rect 533981 274891 534047 274894
rect 560201 274954 560267 274957
rect 560201 274952 567210 274954
rect 560201 274896 560206 274952
rect 560262 274896 567210 274952
rect 560201 274894 567210 274896
rect 560201 274891 560267 274894
rect 534165 274818 534231 274821
rect 539542 274818 539548 274820
rect 534165 274816 539548 274818
rect 534165 274760 534170 274816
rect 534226 274760 539548 274816
rect 534165 274758 539548 274760
rect 534165 274755 534231 274758
rect 539542 274756 539548 274758
rect 539612 274756 539618 274820
rect 553301 274818 553367 274821
rect 550590 274816 553367 274818
rect 550590 274760 553306 274816
rect 553362 274760 553367 274816
rect 550590 274758 553367 274760
rect 567150 274818 567210 274894
rect 583342 274818 583402 275710
rect 583520 275620 584960 275710
rect 567150 274758 576778 274818
rect 521510 274620 521516 274684
rect 521580 274682 521586 274684
rect 549161 274682 549227 274685
rect 550590 274682 550650 274758
rect 553301 274755 553367 274758
rect 521580 274622 521762 274682
rect 521580 274620 521586 274622
rect 521702 274410 521762 274622
rect 549161 274680 550650 274682
rect 549161 274624 549166 274680
rect 549222 274624 550650 274680
rect 549161 274622 550650 274624
rect 576718 274682 576778 274758
rect 576902 274758 583402 274818
rect 576902 274682 576962 274758
rect 576718 274622 576962 274682
rect 549161 274619 549227 274622
rect 526437 274410 526503 274413
rect 521702 274408 526503 274410
rect 521702 274352 526442 274408
rect 526498 274352 526503 274408
rect 521702 274350 526503 274352
rect 526437 274347 526503 274350
rect -960 265706 480 265796
rect 2773 265706 2839 265709
rect -960 265704 2839 265706
rect -960 265648 2778 265704
rect 2834 265648 2839 265704
rect -960 265646 2839 265648
rect -960 265556 480 265646
rect 2773 265643 2839 265646
rect 580625 263938 580691 263941
rect 583520 263938 584960 264028
rect 580625 263936 584960 263938
rect 580625 263880 580630 263936
rect 580686 263880 584960 263936
rect 580625 263878 584960 263880
rect 580625 263875 580691 263878
rect 583520 263788 584960 263878
rect 579705 252242 579771 252245
rect 583520 252242 584960 252332
rect 579705 252240 584960 252242
rect 579705 252184 579710 252240
rect 579766 252184 584960 252240
rect 579705 252182 584960 252184
rect 579705 252179 579771 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3141 251290 3207 251293
rect -960 251288 3207 251290
rect -960 251232 3146 251288
rect 3202 251232 3207 251288
rect -960 251230 3207 251232
rect -960 251140 480 251230
rect 3141 251227 3207 251230
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 3141 237010 3207 237013
rect -960 237008 3207 237010
rect -960 236952 3146 237008
rect 3202 236952 3207 237008
rect -960 236950 3207 236952
rect -960 236860 480 236950
rect 3141 236947 3207 236950
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 3693 222594 3759 222597
rect -960 222592 3759 222594
rect -960 222536 3698 222592
rect 3754 222536 3759 222592
rect -960 222534 3759 222536
rect -960 222444 480 222534
rect 3693 222531 3759 222534
rect 580533 217018 580599 217021
rect 583520 217018 584960 217108
rect 580533 217016 584960 217018
rect 580533 216960 580538 217016
rect 580594 216960 584960 217016
rect 580533 216958 584960 216960
rect 580533 216955 580599 216958
rect 583520 216868 584960 216958
rect -960 208178 480 208268
rect 3325 208178 3391 208181
rect -960 208176 3391 208178
rect -960 208120 3330 208176
rect 3386 208120 3391 208176
rect -960 208118 3391 208120
rect -960 208028 480 208118
rect 3325 208115 3391 208118
rect 580165 205322 580231 205325
rect 583520 205322 584960 205412
rect 580165 205320 584960 205322
rect 580165 205264 580170 205320
rect 580226 205264 584960 205320
rect 580165 205262 584960 205264
rect 580165 205259 580231 205262
rect 583520 205172 584960 205262
rect -960 193898 480 193988
rect 3049 193898 3115 193901
rect -960 193896 3115 193898
rect -960 193840 3054 193896
rect 3110 193840 3115 193896
rect -960 193838 3115 193840
rect -960 193748 480 193838
rect 3049 193835 3115 193838
rect 583520 193476 584960 193716
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 2773 179482 2839 179485
rect -960 179480 2839 179482
rect -960 179424 2778 179480
rect 2834 179424 2839 179480
rect -960 179422 2839 179424
rect -960 179332 480 179422
rect 2773 179419 2839 179422
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 3141 165066 3207 165069
rect -960 165064 3207 165066
rect -960 165008 3146 165064
rect 3202 165008 3207 165064
rect -960 165006 3207 165008
rect -960 164916 480 165006
rect 3141 165003 3207 165006
rect 580165 158402 580231 158405
rect 583520 158402 584960 158492
rect 580165 158400 584960 158402
rect 580165 158344 580170 158400
rect 580226 158344 584960 158400
rect 580165 158342 584960 158344
rect 580165 158339 580231 158342
rect 583520 158252 584960 158342
rect -960 150786 480 150876
rect 3325 150786 3391 150789
rect -960 150784 3391 150786
rect -960 150728 3330 150784
rect 3386 150728 3391 150784
rect -960 150726 3391 150728
rect -960 150636 480 150726
rect 3325 150723 3391 150726
rect 583520 146556 584960 146796
rect -960 136370 480 136460
rect 3509 136370 3575 136373
rect -960 136368 3575 136370
rect -960 136312 3514 136368
rect 3570 136312 3575 136368
rect -960 136310 3575 136312
rect -960 136220 480 136310
rect 3509 136307 3575 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 580441 123178 580507 123181
rect 583520 123178 584960 123268
rect 580441 123176 584960 123178
rect 580441 123120 580446 123176
rect 580502 123120 584960 123176
rect 580441 123118 584960 123120
rect 580441 123115 580507 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 2957 122090 3023 122093
rect -960 122088 3023 122090
rect -960 122032 2962 122088
rect 3018 122032 3023 122088
rect -960 122030 3023 122032
rect -960 121940 480 122030
rect 2957 122027 3023 122030
rect 579613 111482 579679 111485
rect 583520 111482 584960 111572
rect 579613 111480 584960 111482
rect 579613 111424 579618 111480
rect 579674 111424 584960 111480
rect 579613 111422 584960 111424
rect 579613 111419 579679 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3233 107674 3299 107677
rect -960 107672 3299 107674
rect -960 107616 3238 107672
rect 3294 107616 3299 107672
rect -960 107614 3299 107616
rect -960 107524 480 107614
rect 3233 107611 3299 107614
rect 583520 99636 584960 99876
rect -960 93258 480 93348
rect 2773 93258 2839 93261
rect -960 93256 2839 93258
rect -960 93200 2778 93256
rect 2834 93200 2839 93256
rect -960 93198 2839 93200
rect -960 93108 480 93198
rect 2773 93195 2839 93198
rect 583520 87954 584960 88044
rect 583342 87894 584960 87954
rect 539542 87348 539548 87412
rect 539612 87410 539618 87412
rect 549161 87410 549227 87413
rect 539612 87408 549227 87410
rect 539612 87352 549166 87408
rect 549222 87352 549227 87408
rect 539612 87350 549227 87352
rect 539612 87348 539618 87350
rect 549161 87347 549227 87350
rect 533981 87274 534047 87277
rect 524462 87272 534047 87274
rect 524462 87216 533986 87272
rect 534042 87216 534047 87272
rect 524462 87214 534047 87216
rect 521510 86940 521516 87004
rect 521580 87002 521586 87004
rect 524462 87002 524522 87214
rect 533981 87211 534047 87214
rect 560201 87274 560267 87277
rect 560201 87272 567210 87274
rect 560201 87216 560206 87272
rect 560262 87216 567210 87272
rect 560201 87214 567210 87216
rect 560201 87211 560267 87214
rect 534165 87138 534231 87141
rect 539542 87138 539548 87140
rect 534165 87136 539548 87138
rect 534165 87080 534170 87136
rect 534226 87080 539548 87136
rect 534165 87078 539548 87080
rect 534165 87075 534231 87078
rect 539542 87076 539548 87078
rect 539612 87076 539618 87140
rect 553301 87138 553367 87141
rect 550590 87136 553367 87138
rect 550590 87080 553306 87136
rect 553362 87080 553367 87136
rect 550590 87078 553367 87080
rect 567150 87138 567210 87214
rect 583342 87138 583402 87894
rect 583520 87804 584960 87894
rect 567150 87078 576778 87138
rect 521580 86942 524522 87002
rect 549161 87002 549227 87005
rect 550590 87002 550650 87078
rect 553301 87075 553367 87078
rect 549161 87000 550650 87002
rect 549161 86944 549166 87000
rect 549222 86944 550650 87000
rect 549161 86942 550650 86944
rect 576718 87002 576778 87078
rect 576902 87078 583402 87138
rect 576902 87002 576962 87078
rect 576718 86942 576962 87002
rect 521580 86940 521586 86942
rect 549161 86939 549227 86942
rect -960 78978 480 79068
rect 3049 78978 3115 78981
rect -960 78976 3115 78978
rect -960 78920 3054 78976
rect 3110 78920 3115 78976
rect -960 78918 3115 78920
rect -960 78828 480 78918
rect 3049 78915 3115 78918
rect 580349 76258 580415 76261
rect 583520 76258 584960 76348
rect 580349 76256 584960 76258
rect 580349 76200 580354 76256
rect 580410 76200 584960 76256
rect 580349 76198 584960 76200
rect 580349 76195 580415 76198
rect 583520 76108 584960 76198
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 580165 64562 580231 64565
rect 583520 64562 584960 64652
rect 580165 64560 584960 64562
rect 580165 64504 580170 64560
rect 580226 64504 584960 64560
rect 580165 64502 584960 64504
rect 580165 64499 580231 64502
rect 583520 64412 584960 64502
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 522246 44644 522252 44708
rect 522316 44706 522322 44708
rect 524689 44706 524755 44709
rect 522316 44704 524755 44706
rect 522316 44648 524694 44704
rect 524750 44648 524755 44704
rect 522316 44646 524755 44648
rect 522316 44644 522322 44646
rect 524689 44643 524755 44646
rect 44081 42122 44147 42125
rect 79225 42122 79291 42125
rect 44081 42120 79291 42122
rect 44081 42064 44086 42120
rect 44142 42064 79230 42120
rect 79286 42064 79291 42120
rect 44081 42062 79291 42064
rect 44081 42059 44147 42062
rect 79225 42059 79291 42062
rect 100661 42122 100727 42125
rect 126237 42122 126303 42125
rect 100661 42120 126303 42122
rect 100661 42064 100666 42120
rect 100722 42064 126242 42120
rect 126298 42064 126303 42120
rect 100661 42062 126303 42064
rect 100661 42059 100727 42062
rect 126237 42059 126303 42062
rect 583520 41034 584960 41124
rect 583342 40974 584960 41034
rect 531262 40700 531268 40764
rect 531332 40762 531338 40764
rect 540881 40762 540947 40765
rect 531332 40760 540947 40762
rect 531332 40704 540886 40760
rect 540942 40704 540947 40760
rect 531332 40702 540947 40704
rect 531332 40700 531338 40702
rect 540881 40699 540947 40702
rect 524689 40490 524755 40493
rect 531262 40490 531268 40492
rect 524689 40488 531268 40490
rect 524689 40432 524694 40488
rect 524750 40432 531268 40488
rect 524689 40430 531268 40432
rect 524689 40427 524755 40430
rect 531262 40428 531268 40430
rect 531332 40428 531338 40492
rect 565077 40490 565143 40493
rect 560342 40488 565143 40490
rect 560342 40432 565082 40488
rect 565138 40432 565143 40488
rect 560342 40430 565143 40432
rect 540881 40354 540947 40357
rect 540881 40352 543842 40354
rect 540881 40296 540886 40352
rect 540942 40296 543842 40352
rect 540881 40294 543842 40296
rect 540881 40291 540947 40294
rect 543782 40082 543842 40294
rect 560201 40218 560267 40221
rect 560342 40218 560402 40430
rect 565077 40427 565143 40430
rect 572621 40218 572687 40221
rect 583342 40218 583402 40974
rect 583520 40884 584960 40974
rect 560201 40216 560402 40218
rect 560201 40160 560206 40216
rect 560262 40160 560402 40216
rect 560201 40158 560402 40160
rect 569910 40216 572687 40218
rect 569910 40160 572626 40216
rect 572682 40160 572687 40216
rect 569910 40158 572687 40160
rect 560201 40155 560267 40158
rect 550582 40082 550588 40084
rect 543782 40022 550588 40082
rect 550582 40020 550588 40022
rect 550652 40020 550658 40084
rect 565077 40082 565143 40085
rect 569910 40082 569970 40158
rect 572621 40155 572687 40158
rect 576902 40158 583402 40218
rect 565077 40080 569970 40082
rect 565077 40024 565082 40080
rect 565138 40024 569970 40080
rect 565077 40022 569970 40024
rect 572713 40082 572779 40085
rect 576902 40082 576962 40158
rect 572713 40080 576962 40082
rect 572713 40024 572718 40080
rect 572774 40024 576962 40080
rect 572713 40022 576962 40024
rect 565077 40019 565143 40022
rect 572713 40019 572779 40022
rect 550582 39748 550588 39812
rect 550652 39810 550658 39812
rect 560201 39810 560267 39813
rect 550652 39808 560267 39810
rect 550652 39752 560206 39808
rect 560262 39752 560267 39808
rect 550652 39750 560267 39752
rect 550652 39748 550658 39750
rect 560201 39747 560267 39750
rect 74349 38858 74415 38861
rect 73294 38856 74415 38858
rect 73294 38800 74354 38856
rect 74410 38800 74415 38856
rect 73294 38798 74415 38800
rect 73294 38722 73354 38798
rect 74349 38795 74415 38798
rect 73429 38722 73495 38725
rect 73294 38720 73495 38722
rect 73294 38664 73434 38720
rect 73490 38664 73495 38720
rect 73294 38662 73495 38664
rect 73429 38659 73495 38662
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 580257 29338 580323 29341
rect 583520 29338 584960 29428
rect 580257 29336 584960 29338
rect 580257 29280 580262 29336
rect 580318 29280 584960 29336
rect 580257 29278 584960 29280
rect 580257 29275 580323 29278
rect 118141 29202 118207 29205
rect 117270 29200 118207 29202
rect 117270 29144 118146 29200
rect 118202 29144 118207 29200
rect 583520 29188 584960 29278
rect 117270 29142 118207 29144
rect 117270 29066 117330 29142
rect 118141 29139 118207 29142
rect 117405 29066 117471 29069
rect 117270 29064 117471 29066
rect 117270 29008 117410 29064
rect 117466 29008 117471 29064
rect 117270 29006 117471 29008
rect 117405 29003 117471 29006
rect 121085 27842 121151 27845
rect 120030 27840 121151 27842
rect 120030 27784 121090 27840
rect 121146 27784 121151 27840
rect 120030 27782 121151 27784
rect 120030 27706 120090 27782
rect 121085 27779 121151 27782
rect 120165 27706 120231 27709
rect 120030 27704 120231 27706
rect 120030 27648 120170 27704
rect 120226 27648 120231 27704
rect 120030 27646 120231 27648
rect 120165 27643 120231 27646
rect 518014 21994 518020 21996
rect 614 21934 518020 21994
rect -960 21450 480 21540
rect 614 21450 674 21934
rect 518014 21932 518020 21934
rect 518084 21932 518090 21996
rect -960 21390 674 21450
rect -960 21300 480 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect 31477 9754 31543 9757
rect 31661 9754 31727 9757
rect 31477 9752 31727 9754
rect 31477 9696 31482 9752
rect 31538 9696 31666 9752
rect 31722 9696 31727 9752
rect 31477 9694 31727 9696
rect 31477 9691 31543 9694
rect 31661 9691 31727 9694
rect 108757 9754 108823 9757
rect 108941 9754 109007 9757
rect 108757 9752 109007 9754
rect 108757 9696 108762 9752
rect 108818 9696 108946 9752
rect 109002 9696 109007 9752
rect 108757 9694 109007 9696
rect 108757 9691 108823 9694
rect 108941 9691 109007 9694
rect 3417 8258 3483 8261
rect 516358 8258 516364 8260
rect 3417 8256 516364 8258
rect 3417 8200 3422 8256
rect 3478 8200 516364 8256
rect 3417 8198 516364 8200
rect 3417 8195 3483 8198
rect 516358 8196 516364 8198
rect 516428 8196 516434 8260
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
rect 442901 3362 442967 3365
rect 484577 3362 484643 3365
rect 442901 3360 484643 3362
rect 442901 3304 442906 3360
rect 442962 3304 484582 3360
rect 484638 3304 484643 3360
rect 442901 3302 484643 3304
rect 442901 3299 442967 3302
rect 484577 3299 484643 3302
rect 547229 3362 547295 3365
rect 582189 3362 582255 3365
rect 547229 3360 582255 3362
rect 547229 3304 547234 3360
rect 547290 3304 582194 3360
rect 582250 3304 582255 3360
rect 547229 3302 582255 3304
rect 547229 3299 547295 3302
rect 582189 3299 582255 3302
rect 441429 3090 441495 3093
rect 447041 3090 447107 3093
rect 441429 3088 447107 3090
rect 441429 3032 441434 3088
rect 441490 3032 447046 3088
rect 447102 3032 447107 3088
rect 441429 3030 447107 3032
rect 441429 3027 441495 3030
rect 447041 3027 447107 3030
<< via3 >>
rect 521516 646716 521580 646780
rect 520596 646580 520660 646644
rect 125732 646444 125796 646508
rect 521148 646444 521212 646508
rect 520964 646308 521028 646372
rect 520780 646172 520844 646236
rect 471284 645900 471348 645964
rect 125732 643784 125796 643788
rect 125732 643728 125782 643784
rect 125782 643728 125796 643784
rect 125732 643724 125796 643728
rect 50844 643316 50908 643380
rect 75316 643376 75380 643380
rect 75316 643320 75330 643376
rect 75330 643320 75380 643376
rect 75316 643316 75380 643320
rect 100524 643376 100588 643380
rect 100524 643320 100538 643376
rect 100538 643320 100588 643376
rect 100524 643316 100588 643320
rect 205404 643376 205468 643380
rect 205404 643320 205454 643376
rect 205454 643320 205468 643376
rect 205404 643316 205468 643320
rect 218468 643376 218532 643380
rect 218468 643320 218482 643376
rect 218482 643320 218532 643376
rect 218468 643316 218532 643320
rect 369348 643376 369412 643380
rect 369348 643320 369398 643376
rect 369398 643320 369412 643376
rect 369348 643316 369412 643320
rect 390508 643376 390572 643380
rect 390508 643320 390558 643376
rect 390558 643320 390572 643376
rect 390508 643316 390572 643320
rect 394740 643376 394804 643380
rect 394740 643320 394790 643376
rect 394790 643320 394804 643376
rect 394740 643316 394804 643320
rect 453620 643376 453684 643380
rect 453620 643320 453670 643376
rect 453670 643320 453684 643376
rect 453620 643316 453684 643320
rect 516364 643316 516428 643380
rect 518020 643316 518084 643380
rect 240916 643044 240980 643108
rect 253796 643044 253860 643108
rect 264468 643044 264532 643108
rect 273116 643044 273180 643108
rect 282868 643044 282932 643108
rect 311756 643044 311820 643108
rect 335308 643044 335372 643108
rect 349660 643044 349724 643108
rect 350764 643044 350828 643108
rect 369716 643044 369780 643108
rect 100524 642772 100588 642836
rect 75316 642636 75380 642700
rect 453620 642500 453684 642564
rect 471284 642364 471348 642428
rect 390508 642228 390572 642292
rect 369348 642092 369412 642156
rect 379652 642092 379716 642156
rect 391244 642092 391308 642156
rect 218468 641956 218532 642020
rect 75868 641820 75932 641884
rect 85436 641820 85500 641884
rect 95188 641820 95252 641884
rect 104756 641820 104820 641884
rect 153148 641820 153212 641884
rect 162532 641820 162596 641884
rect 164188 641820 164252 641884
rect 178724 641820 178788 641884
rect 186268 641820 186332 641884
rect 195836 641820 195900 641884
rect 205404 641820 205468 641884
rect 394740 641684 394804 641748
rect 398788 641684 398852 641748
rect 410564 641684 410628 641748
rect 418108 641684 418172 641748
rect 427676 641684 427740 641748
rect 442948 641684 443012 641748
rect 452516 641684 452580 641748
rect 462452 641684 462516 641748
rect 471836 641684 471900 641748
rect 481588 641684 481652 641748
rect 491156 641684 491220 641748
rect 500908 641684 500972 641748
rect 519492 641684 519556 641748
rect 520596 641684 520660 641748
rect 521332 641684 521396 641748
rect 521516 636788 521580 636852
rect 521516 636516 521580 636580
rect 521516 628764 521580 628828
rect 521516 627948 521580 628012
rect 521516 616796 521580 616860
rect 521516 610132 521580 610196
rect 521516 607004 521580 607068
rect 521884 563212 521948 563276
rect 521516 562668 521580 562732
rect 521516 556548 521580 556612
rect 539548 462708 539612 462772
rect 539548 462436 539612 462500
rect 521516 462300 521580 462364
rect 539548 275028 539612 275092
rect 539548 274756 539612 274820
rect 521516 274620 521580 274684
rect 539548 87348 539612 87412
rect 521516 86940 521580 87004
rect 539548 87076 539612 87140
rect 522252 44644 522316 44708
rect 531268 40700 531332 40764
rect 531268 40428 531332 40492
rect 550588 40020 550652 40084
rect 550588 39748 550652 39812
rect 518020 21932 518084 21996
rect 516364 8196 516428 8260
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 50843 643380 50909 643381
rect 50843 643316 50844 643380
rect 50908 643316 50909 643380
rect 50843 643315 50909 643316
rect 50846 641698 50906 643315
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 75315 643380 75381 643381
rect 75315 643316 75316 643380
rect 75380 643316 75381 643380
rect 75315 643315 75381 643316
rect 75318 642701 75378 643315
rect 75315 642700 75381 642701
rect 75315 642636 75316 642700
rect 75380 642636 75381 642700
rect 75315 642635 75381 642636
rect 75867 641884 75933 641885
rect 75867 641820 75868 641884
rect 75932 641820 75933 641884
rect 75867 641819 75933 641820
rect 75870 641698 75930 641819
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 85435 641884 85501 641885
rect 85435 641820 85436 641884
rect 85500 641820 85501 641884
rect 85435 641819 85501 641820
rect 85438 641698 85498 641819
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 95187 641884 95253 641885
rect 95187 641820 95188 641884
rect 95252 641820 95253 641884
rect 95187 641819 95253 641820
rect 95190 641698 95250 641819
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 639654 98604 675098
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 100523 643380 100589 643381
rect 100523 643316 100524 643380
rect 100588 643316 100589 643380
rect 100523 643315 100589 643316
rect 100526 642837 100586 643315
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 100523 642836 100589 642837
rect 100523 642772 100524 642836
rect 100588 642772 100589 642836
rect 100523 642771 100589 642772
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 104755 641884 104821 641885
rect 104755 641820 104756 641884
rect 104820 641820 104821 641884
rect 104755 641819 104821 641820
rect 104758 641698 104818 641819
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 125731 646508 125797 646509
rect 125731 646444 125732 646508
rect 125796 646444 125797 646508
rect 125731 646443 125797 646444
rect 125734 643789 125794 646443
rect 125731 643788 125797 643789
rect 125731 643724 125732 643788
rect 125796 643724 125797 643788
rect 125731 643723 125797 643724
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 136002 641550 136502 641610
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 153147 641884 153213 641885
rect 153147 641820 153148 641884
rect 153212 641820 153213 641884
rect 153147 641819 153213 641820
rect 153150 641698 153210 641819
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 625254 156204 660698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162531 641884 162597 641885
rect 162531 641820 162532 641884
rect 162596 641820 162597 641884
rect 162531 641819 162597 641820
rect 162534 641698 162594 641819
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 632454 163404 667898
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 164187 641884 164253 641885
rect 164187 641820 164188 641884
rect 164252 641820 164253 641884
rect 164187 641819 164253 641820
rect 164190 641698 164250 641819
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 178723 641884 178789 641885
rect 178723 641820 178724 641884
rect 178788 641820 178789 641884
rect 178723 641819 178789 641820
rect 178726 641698 178786 641819
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 186267 641884 186333 641885
rect 186267 641820 186268 641884
rect 186332 641820 186333 641884
rect 186267 641819 186333 641820
rect 186270 641698 186330 641819
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 195835 641884 195901 641885
rect 195835 641820 195836 641884
rect 195900 641820 195901 641884
rect 195835 641819 195901 641820
rect 195838 641698 195898 641819
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 205403 643380 205469 643381
rect 205403 643316 205404 643380
rect 205468 643316 205469 643380
rect 205403 643315 205469 643316
rect 205406 641885 205466 643315
rect 205403 641884 205469 641885
rect 205403 641820 205404 641884
rect 205468 641820 205469 641884
rect 205403 641819 205469 641820
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 218467 643380 218533 643381
rect 218467 643316 218468 643380
rect 218532 643316 218533 643380
rect 218467 643315 218533 643316
rect 218470 642021 218530 643315
rect 218467 642020 218533 642021
rect 218467 641956 218468 642020
rect 218532 641956 218533 642020
rect 218467 641955 218533 641956
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 240915 643108 240981 643109
rect 240915 643044 240916 643108
rect 240980 643044 240981 643108
rect 240915 643043 240981 643044
rect 240918 641698 240978 643043
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 387654 242604 423098
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 253795 643108 253861 643109
rect 253795 643044 253796 643108
rect 253860 643044 253861 643108
rect 253795 643043 253861 643044
rect 253798 641698 253858 643043
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 264467 643108 264533 643109
rect 264467 643044 264468 643108
rect 264532 643044 264533 643108
rect 264467 643043 264533 643044
rect 264470 641698 264530 643043
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 632454 271404 667898
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 273115 643108 273181 643109
rect 273115 643044 273116 643108
rect 273180 643044 273181 643108
rect 273115 643043 273181 643044
rect 273118 641698 273178 643043
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 282867 643108 282933 643109
rect 282867 643044 282868 643108
rect 282932 643044 282933 643108
rect 282867 643043 282933 643044
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 282870 641698 282930 643043
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 311755 643108 311821 643109
rect 311755 643044 311756 643108
rect 311820 643044 311821 643108
rect 311755 643043 311821 643044
rect 311758 641698 311818 643043
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335307 643108 335373 643109
rect 335307 643044 335308 643108
rect 335372 643044 335373 643108
rect 335307 643043 335373 643044
rect 335310 641698 335370 643043
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 349659 643108 349725 643109
rect 349659 643044 349660 643108
rect 349724 643044 349725 643108
rect 349659 643043 349725 643044
rect 349662 641698 349722 643043
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 639654 350604 675098
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 350763 643108 350829 643109
rect 350763 643044 350764 643108
rect 350828 643044 350829 643108
rect 350763 643043 350829 643044
rect 350766 641698 350826 643043
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 369347 643380 369413 643381
rect 369347 643316 369348 643380
rect 369412 643316 369413 643380
rect 369347 643315 369413 643316
rect 369350 642157 369410 643315
rect 369715 643108 369781 643109
rect 369715 643044 369716 643108
rect 369780 643044 369781 643108
rect 369715 643043 369781 643044
rect 369347 642156 369413 642157
rect 369347 642092 369348 642156
rect 369412 642092 369413 642156
rect 369347 642091 369413 642092
rect 369718 641698 369778 643043
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 379651 642156 379717 642157
rect 379651 642092 379652 642156
rect 379716 642092 379717 642156
rect 379651 642091 379717 642092
rect 379654 641698 379714 642091
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 390507 643380 390573 643381
rect 390507 643316 390508 643380
rect 390572 643316 390573 643380
rect 390507 643315 390573 643316
rect 394739 643380 394805 643381
rect 394739 643316 394740 643380
rect 394804 643316 394805 643380
rect 394739 643315 394805 643316
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 390510 642293 390570 643315
rect 390507 642292 390573 642293
rect 390507 642228 390508 642292
rect 390572 642228 390573 642292
rect 390507 642227 390573 642228
rect 391243 642156 391309 642157
rect 391243 642092 391244 642156
rect 391308 642092 391309 642156
rect 391243 642091 391309 642092
rect 391246 641698 391306 642091
rect 394742 641749 394802 643315
rect 394739 641748 394805 641749
rect 394739 641684 394740 641748
rect 394804 641684 394805 641748
rect 394739 641683 394805 641684
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 614454 397404 649898
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 398787 641748 398853 641749
rect 398787 641698 398788 641748
rect 398852 641698 398853 641748
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 410563 641748 410629 641749
rect 410563 641698 410564 641748
rect 410628 641698 410629 641748
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 632454 415404 667898
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418107 641748 418173 641749
rect 418107 641698 418108 641748
rect 418172 641698 418173 641748
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 427675 641748 427741 641749
rect 427675 641698 427676 641748
rect 427740 641698 427741 641748
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 442947 641748 443013 641749
rect 442947 641698 442948 641748
rect 443012 641698 443013 641748
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 453619 643380 453685 643381
rect 453619 643316 453620 643380
rect 453684 643316 453685 643380
rect 453619 643315 453685 643316
rect 453622 642565 453682 643315
rect 453619 642564 453685 642565
rect 453619 642500 453620 642564
rect 453684 642500 453685 642564
rect 453619 642499 453685 642500
rect 452515 641748 452581 641749
rect 452515 641698 452516 641748
rect 452580 641698 452581 641748
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 462451 641748 462517 641749
rect 462451 641698 462452 641748
rect 462516 641698 462517 641748
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 468804 614454 469404 649898
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 471283 645964 471349 645965
rect 471283 645900 471284 645964
rect 471348 645900 471349 645964
rect 471283 645899 471349 645900
rect 471286 642429 471346 645899
rect 471283 642428 471349 642429
rect 471283 642364 471284 642428
rect 471348 642364 471349 642428
rect 471283 642363 471349 642364
rect 471835 641748 471901 641749
rect 471835 641698 471836 641748
rect 471900 641698 471901 641748
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 481587 641748 481653 641749
rect 481587 641698 481588 641748
rect 481652 641698 481653 641748
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 491155 641748 491221 641749
rect 491155 641698 491156 641748
rect 491220 641698 491221 641748
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 500907 641748 500973 641749
rect 500907 641698 500908 641748
rect 500972 641698 500973 641748
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 521515 646780 521581 646781
rect 521515 646716 521516 646780
rect 521580 646716 521581 646780
rect 521515 646715 521581 646716
rect 520595 646644 520661 646645
rect 520595 646580 520596 646644
rect 520660 646580 520661 646644
rect 520595 646579 520661 646580
rect 516363 643380 516429 643381
rect 516363 643316 516364 643380
rect 516428 643316 516429 643380
rect 516363 643315 516429 643316
rect 518019 643380 518085 643381
rect 518019 643316 518020 643380
rect 518084 643316 518085 643380
rect 518019 643315 518085 643316
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 516366 8261 516426 643315
rect 518022 21997 518082 643315
rect 520598 641749 520658 646579
rect 521147 646508 521213 646509
rect 521147 646444 521148 646508
rect 521212 646444 521213 646508
rect 521147 646443 521213 646444
rect 520963 646372 521029 646373
rect 520963 646308 520964 646372
rect 521028 646308 521029 646372
rect 520963 646307 521029 646308
rect 520779 646236 520845 646237
rect 520779 646172 520780 646236
rect 520844 646172 520845 646236
rect 520779 646171 520845 646172
rect 519491 641748 519557 641749
rect 519491 641698 519492 641748
rect 519556 641698 519557 641748
rect 520595 641748 520661 641749
rect 520595 641684 520596 641748
rect 520660 641684 520661 641748
rect 520595 641683 520661 641684
rect 520782 611690 520842 646171
rect 520230 611630 520842 611690
rect 520230 610330 520290 611630
rect 520230 610270 520842 610330
rect 520782 88770 520842 610270
rect 520966 279170 521026 646307
rect 521150 464810 521210 646443
rect 521331 641748 521397 641749
rect 521331 641684 521332 641748
rect 521396 641684 521397 641748
rect 521331 641683 521397 641684
rect 521334 606930 521394 641683
rect 521518 636853 521578 646715
rect 521515 636852 521581 636853
rect 521515 636788 521516 636852
rect 521580 636788 521581 636852
rect 521515 636787 521581 636788
rect 521515 636580 521581 636581
rect 521515 636516 521516 636580
rect 521580 636516 521581 636580
rect 521515 636515 521581 636516
rect 521518 628829 521578 636515
rect 521515 628828 521581 628829
rect 521515 628764 521516 628828
rect 521580 628764 521581 628828
rect 521515 628763 521581 628764
rect 521515 628012 521581 628013
rect 521515 627948 521516 628012
rect 521580 627948 521581 628012
rect 521515 627947 521581 627948
rect 521518 616861 521578 627947
rect 521515 616860 521581 616861
rect 521515 616796 521516 616860
rect 521580 616796 521581 616860
rect 521515 616795 521581 616796
rect 521515 610196 521581 610197
rect 521515 610132 521516 610196
rect 521580 610132 521581 610196
rect 521515 610131 521581 610132
rect 521518 607069 521578 610131
rect 521515 607068 521581 607069
rect 521515 607004 521516 607068
rect 521580 607004 521581 607068
rect 521515 607003 521581 607004
rect 521334 606870 521762 606930
rect 521702 591290 521762 606870
rect 521518 591230 521762 591290
rect 521518 583130 521578 591230
rect 521518 583070 521762 583130
rect 521702 574970 521762 583070
rect 521702 574910 522130 574970
rect 522070 570210 522130 574910
rect 521886 570150 522130 570210
rect 521886 563277 521946 570150
rect 521883 563276 521949 563277
rect 521883 563212 521884 563276
rect 521948 563212 521949 563276
rect 521883 563211 521949 563212
rect 521515 562732 521581 562733
rect 521515 562730 521516 562732
rect 521334 562670 521516 562730
rect 521334 556610 521394 562670
rect 521515 562668 521516 562670
rect 521580 562668 521581 562732
rect 521515 562667 521581 562668
rect 521515 556612 521581 556613
rect 521515 556610 521516 556612
rect 521334 556550 521516 556610
rect 521515 556548 521516 556550
rect 521580 556548 521581 556612
rect 521515 556547 521581 556548
rect 521150 464750 521394 464810
rect 521334 462090 521394 464750
rect 521515 462364 521581 462365
rect 521515 462300 521516 462364
rect 521580 462300 521581 462364
rect 521515 462299 521581 462300
rect 521518 462090 521578 462299
rect 521334 462030 521578 462090
rect 520966 279110 521394 279170
rect 521334 274410 521394 279110
rect 521515 274684 521581 274685
rect 521515 274620 521516 274684
rect 521580 274620 521581 274684
rect 521515 274619 521581 274620
rect 521518 274410 521578 274619
rect 521334 274350 521578 274410
rect 520782 88710 521394 88770
rect 521334 86730 521394 88710
rect 521515 87004 521581 87005
rect 521515 86940 521516 87004
rect 521580 86940 521581 87004
rect 521515 86939 521581 86940
rect 521518 86730 521578 86939
rect 521334 86670 521578 86730
rect 522254 44709 522314 641462
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522251 44708 522317 44709
rect 522251 44644 522252 44708
rect 522316 44644 522317 44708
rect 522251 44643 522317 44644
rect 518019 21996 518085 21997
rect 518019 21932 518020 21996
rect 518084 21932 518085 21996
rect 518019 21931 518085 21932
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 516363 8260 516429 8261
rect 516363 8196 516364 8260
rect 516428 8196 516429 8260
rect 516363 8195 516429 8196
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 539547 462772 539613 462773
rect 539547 462708 539548 462772
rect 539612 462708 539613 462772
rect 539547 462707 539613 462708
rect 533604 427254 534204 462698
rect 539550 462501 539610 462707
rect 539547 462500 539613 462501
rect 539547 462436 539548 462500
rect 539612 462436 539613 462500
rect 539547 462435 539613 462436
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 539547 275092 539613 275093
rect 539547 275028 539548 275092
rect 539612 275028 539613 275092
rect 539547 275027 539613 275028
rect 539550 274821 539610 275027
rect 539547 274820 539613 274821
rect 539547 274756 539548 274820
rect 539612 274756 539613 274820
rect 539547 274755 539613 274756
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 539547 87412 539613 87413
rect 539547 87348 539548 87412
rect 539612 87348 539613 87412
rect 539547 87347 539613 87348
rect 539550 87141 539610 87347
rect 539547 87140 539613 87141
rect 539547 87076 539548 87140
rect 539612 87076 539613 87140
rect 539547 87075 539613 87076
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 531267 40764 531333 40765
rect 531267 40700 531268 40764
rect 531332 40700 531333 40764
rect 531267 40699 531333 40700
rect 531270 40493 531330 40699
rect 531267 40492 531333 40493
rect 531267 40428 531268 40492
rect 531332 40428 531333 40492
rect 531267 40427 531333 40428
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 550587 40084 550653 40085
rect 550587 40020 550588 40084
rect 550652 40020 550653 40084
rect 550587 40019 550653 40020
rect 550590 39813 550650 40019
rect 550587 39812 550653 39813
rect 550587 39748 550588 39812
rect 550652 39748 550653 39812
rect 550587 39747 550653 39748
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 50758 641462 50994 641698
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 75782 641462 76018 641698
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 85350 641462 85586 641698
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 95102 641462 95338 641698
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 101786 642698 102022 642934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 104670 641462 104906 641698
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 135766 641462 136002 641698
rect 136502 641462 136738 641698
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 153062 641462 153298 641698
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162446 641462 162682 641698
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 164102 641462 164338 641698
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 178638 641462 178874 641698
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 186182 641462 186418 641698
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 195750 641462 195986 641698
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 240830 641462 241066 641698
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 253710 641462 253946 641698
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 264382 641462 264618 641698
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 273030 641462 273266 641698
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 281786 642698 282022 642934
rect 282782 641462 283018 641698
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 311670 641462 311906 641698
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335222 641462 335458 641698
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 349574 641462 349810 641698
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 350678 641462 350914 641698
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 369630 641462 369866 641698
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 379566 641462 379802 641698
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 391158 641462 391394 641698
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 398702 641684 398788 641698
rect 398788 641684 398852 641698
rect 398852 641684 398938 641698
rect 398702 641462 398938 641684
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 410478 641684 410564 641698
rect 410564 641684 410628 641698
rect 410628 641684 410714 641698
rect 410478 641462 410714 641684
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418022 641684 418108 641698
rect 418108 641684 418172 641698
rect 418172 641684 418258 641698
rect 418022 641462 418258 641684
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 427590 641684 427676 641698
rect 427676 641684 427740 641698
rect 427740 641684 427826 641698
rect 427590 641462 427826 641684
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 442862 641684 442948 641698
rect 442948 641684 443012 641698
rect 443012 641684 443098 641698
rect 442862 641462 443098 641684
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 452430 641684 452516 641698
rect 452516 641684 452580 641698
rect 452580 641684 452666 641698
rect 452430 641462 452666 641684
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 462366 641684 462452 641698
rect 462452 641684 462516 641698
rect 462516 641684 462602 641698
rect 462366 641462 462602 641684
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 471750 641684 471836 641698
rect 471836 641684 471900 641698
rect 471900 641684 471986 641698
rect 471750 641462 471986 641684
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 481502 641684 481588 641698
rect 481588 641684 481652 641698
rect 481652 641684 481738 641698
rect 481502 641462 481738 641684
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 491070 641684 491156 641698
rect 491156 641684 491220 641698
rect 491220 641684 491306 641698
rect 491070 641462 491306 641684
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 500822 641684 500908 641698
rect 500908 641684 500972 641698
rect 500972 641684 501058 641698
rect 500822 641462 501058 641684
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 519406 641684 519492 641698
rect 519492 641684 519556 641698
rect 519556 641684 519642 641698
rect 519406 641462 519642 641684
rect 522166 641462 522402 641698
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect 50716 641698 65020 641740
rect 50716 641462 50758 641698
rect 50994 641462 65020 641698
rect 50716 641420 65020 641462
rect 64700 640380 65020 641420
rect 67460 641698 76060 641740
rect 67460 641462 75782 641698
rect 76018 641462 76060 641698
rect 67460 641420 76060 641462
rect 85308 641698 85628 641740
rect 85308 641462 85350 641698
rect 85586 641462 85628 641698
rect 67460 640380 67780 641420
rect 64700 640060 67780 640380
rect 85308 640380 85628 641462
rect 86780 641698 95380 641740
rect 86780 641462 95102 641698
rect 95338 641462 95380 641698
rect 86780 641420 95380 641462
rect 104628 641698 104948 641740
rect 104628 641462 104670 641698
rect 104906 641462 104948 641698
rect 86780 640380 87100 641420
rect 85308 640060 87100 640380
rect 104628 640380 104948 641462
rect 106100 641420 117276 641740
rect 106100 640380 106420 641420
rect 116956 641060 117276 641420
rect 125420 641698 136044 641740
rect 125420 641462 135766 641698
rect 136002 641462 136044 641698
rect 125420 641420 136044 641462
rect 136460 641698 143588 641740
rect 136460 641462 136502 641698
rect 136738 641462 143588 641698
rect 136460 641420 143588 641462
rect 116956 640740 124268 641060
rect 104628 640060 106420 640380
rect 123948 640380 124268 640740
rect 125420 640380 125740 641420
rect 123948 640060 125740 640380
rect 143268 640380 143588 641420
rect 144740 641698 153340 641740
rect 144740 641462 153062 641698
rect 153298 641462 153340 641698
rect 144740 641420 153340 641462
rect 162404 641698 164380 642012
rect 162404 641462 162446 641698
rect 162682 641692 164102 641698
rect 162682 641462 162724 641692
rect 162404 641420 162724 641462
rect 164060 641462 164102 641692
rect 164338 641462 164380 641698
rect 164060 641420 164380 641462
rect 178596 641698 186460 641740
rect 178596 641462 178638 641698
rect 178874 641462 186182 641698
rect 186418 641462 186460 641698
rect 178596 641420 186460 641462
rect 195708 641698 196028 641740
rect 195708 641462 195750 641698
rect 195986 641462 196028 641698
rect 144740 640380 145060 641420
rect 195708 641060 196028 641462
rect 201412 641420 210012 641740
rect 195708 640740 200260 641060
rect 143268 640060 145060 640380
rect 199940 640380 200260 640740
rect 201412 640380 201732 641420
rect 199940 640060 201732 640380
rect 209692 640380 210012 641420
rect 212636 641420 220868 641740
rect 212636 640380 212956 641420
rect 209692 640060 212956 640380
rect 220548 640380 220868 641420
rect 226804 641698 241108 641740
rect 226804 641462 240830 641698
rect 241066 641462 241108 641698
rect 226804 641420 241108 641462
rect 253668 641698 264660 641740
rect 253668 641462 253710 641698
rect 253946 641462 264382 641698
rect 264618 641462 264660 641698
rect 253668 641420 264660 641462
rect 272988 641698 283060 641740
rect 272988 641462 273030 641698
rect 273266 641462 282782 641698
rect 283018 641462 283060 641698
rect 272988 641420 283060 641462
rect 311628 641698 311948 641740
rect 311628 641462 311670 641698
rect 311906 641462 311948 641698
rect 226804 640380 227124 641420
rect 253668 640740 254172 641420
rect 272988 640740 273492 641420
rect 311628 641060 311948 641462
rect 318620 641420 325932 641740
rect 311628 640740 316180 641060
rect 220548 640060 227124 640380
rect 315860 640380 316180 640740
rect 318620 640380 318940 641420
rect 325612 641060 325932 641420
rect 335180 641698 335500 641740
rect 335180 641462 335222 641698
rect 335458 641462 335500 641698
rect 335180 641060 335500 641462
rect 325612 640740 335500 641060
rect 349532 641698 349852 641740
rect 349532 641462 349574 641698
rect 349810 641462 349852 641698
rect 349532 641060 349852 641462
rect 350452 641698 350956 641740
rect 350452 641462 350678 641698
rect 350914 641462 350956 641698
rect 350452 641420 350956 641462
rect 369588 641698 379844 641740
rect 369588 641462 369630 641698
rect 369866 641462 379566 641698
rect 379802 641462 379844 641698
rect 369588 641420 379844 641462
rect 391116 641698 398980 641740
rect 391116 641462 391158 641698
rect 391394 641462 398702 641698
rect 398938 641462 398980 641698
rect 391116 641420 398980 641462
rect 410436 641698 418300 641740
rect 410436 641462 410478 641698
rect 410714 641462 418022 641698
rect 418258 641462 418300 641698
rect 410436 641420 418300 641462
rect 427548 641698 427868 641740
rect 427548 641462 427590 641698
rect 427826 641462 427868 641698
rect 350452 641060 350772 641420
rect 349532 640740 350772 641060
rect 369588 640740 370092 641420
rect 427548 641060 427868 641462
rect 434540 641698 443140 641740
rect 434540 641462 442862 641698
rect 443098 641462 443140 641698
rect 434540 641420 443140 641462
rect 452388 641698 452708 641740
rect 452388 641462 452430 641698
rect 452666 641462 452708 641698
rect 427548 640740 432100 641060
rect 315860 640060 318940 640380
rect 431780 640380 432100 640740
rect 434540 640380 434860 641420
rect 431780 640060 434860 640380
rect 452388 640380 452708 641462
rect 453860 641698 462644 641740
rect 453860 641462 462366 641698
rect 462602 641462 462644 641698
rect 453860 641420 462644 641462
rect 471708 641698 472028 641740
rect 471708 641462 471750 641698
rect 471986 641462 472028 641698
rect 453860 640380 454180 641420
rect 452388 640060 454180 640380
rect 471708 640380 472028 641462
rect 473180 641698 481780 641740
rect 473180 641462 481502 641698
rect 481738 641462 481780 641698
rect 473180 641420 481780 641462
rect 491028 641698 491348 641740
rect 491028 641462 491070 641698
rect 491306 641462 491348 641698
rect 473180 640380 473500 641420
rect 471708 640060 473500 640380
rect 491028 640380 491348 641462
rect 492500 641698 501100 641740
rect 492500 641462 500822 641698
rect 501058 641462 501100 641698
rect 492500 641420 501100 641462
rect 519364 641698 522444 641740
rect 519364 641462 519406 641698
rect 519642 641462 522166 641698
rect 522402 641462 522444 641698
rect 519364 641420 522444 641462
rect 492500 640380 492820 641420
rect 491028 640060 492820 640380
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use user_proj_example  mprj
timestamp 1607540551
transform 1 0 44000 0 1 44000
box 0 0 479012 600000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
