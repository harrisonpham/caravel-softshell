VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 2395.060 BY 3000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.840 2996.000 8.120 3000.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 638.960 2996.000 639.240 3000.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 702.440 2996.000 702.720 3000.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 765.460 2996.000 765.740 3000.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 828.480 2996.000 828.760 3000.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 891.960 2996.000 892.240 3000.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 954.980 2996.000 955.260 3000.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1018.000 2996.000 1018.280 3000.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1081.020 2996.000 1081.300 3000.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.500 2996.000 1144.780 3000.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1207.520 2996.000 1207.800 3000.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.860 2996.000 71.140 3000.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1270.540 2996.000 1270.820 3000.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1334.020 2996.000 1334.300 3000.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1397.040 2996.000 1397.320 3000.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1460.060 2996.000 1460.340 3000.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1523.080 2996.000 1523.360 3000.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1586.560 2996.000 1586.840 3000.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.580 2996.000 1649.860 3000.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1712.600 2996.000 1712.880 3000.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1776.080 2996.000 1776.360 3000.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.100 2996.000 1839.380 3000.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.880 2996.000 134.160 3000.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1902.120 2996.000 1902.400 3000.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.140 2996.000 1965.420 3000.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2028.620 2996.000 2028.900 3000.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2091.640 2996.000 2091.920 3000.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2154.660 2996.000 2154.940 3000.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2218.140 2996.000 2218.420 3000.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2281.160 2996.000 2281.440 3000.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2344.180 2996.000 2344.460 3000.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 196.900 2996.000 197.180 3000.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 260.380 2996.000 260.660 3000.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.400 2996.000 323.680 3000.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 386.420 2996.000 386.700 3000.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 449.900 2996.000 450.180 3000.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 512.920 2996.000 513.200 3000.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 575.940 2996.000 576.220 3000.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.540 2996.000 28.820 3000.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 660.120 2996.000 660.400 3000.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 723.140 2996.000 723.420 3000.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 786.620 2996.000 786.900 3000.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 849.640 2996.000 849.920 3000.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 912.660 2996.000 912.940 3000.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 976.140 2996.000 976.420 3000.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1039.160 2996.000 1039.440 3000.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.180 2996.000 1102.460 3000.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1165.200 2996.000 1165.480 3000.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1228.680 2996.000 1228.960 3000.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.020 2996.000 92.300 3000.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1291.700 2996.000 1291.980 3000.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1354.720 2996.000 1355.000 3000.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1418.200 2996.000 1418.480 3000.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1481.220 2996.000 1481.500 3000.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1544.240 2996.000 1544.520 3000.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1607.720 2996.000 1608.000 3000.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1670.740 2996.000 1671.020 3000.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1733.760 2996.000 1734.040 3000.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1796.780 2996.000 1797.060 3000.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1860.260 2996.000 1860.540 3000.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 155.040 2996.000 155.320 3000.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.280 2996.000 1923.560 3000.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1986.300 2996.000 1986.580 3000.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2049.780 2996.000 2050.060 3000.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2112.800 2996.000 2113.080 3000.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2175.820 2996.000 2176.100 3000.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2238.840 2996.000 2239.120 3000.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2302.320 2996.000 2302.600 3000.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2365.340 2996.000 2365.620 3000.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 218.060 2996.000 218.340 3000.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 281.080 2996.000 281.360 3000.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 344.560 2996.000 344.840 3000.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 407.580 2996.000 407.860 3000.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 470.600 2996.000 470.880 3000.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 534.080 2996.000 534.360 3000.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 597.100 2996.000 597.380 3000.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.700 2996.000 49.980 3000.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 681.280 2996.000 681.560 3000.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 744.300 2996.000 744.580 3000.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 807.780 2996.000 808.060 3000.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.800 2996.000 871.080 3000.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 933.820 2996.000 934.100 3000.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 996.840 2996.000 997.120 3000.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1060.320 2996.000 1060.600 3000.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1123.340 2996.000 1123.620 3000.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1186.360 2996.000 1186.640 3000.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1249.840 2996.000 1250.120 3000.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.720 2996.000 113.000 3000.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1312.860 2996.000 1313.140 3000.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1375.880 2996.000 1376.160 3000.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1438.900 2996.000 1439.180 3000.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1502.380 2996.000 1502.660 3000.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1565.400 2996.000 1565.680 3000.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1628.420 2996.000 1628.700 3000.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.900 2996.000 1692.180 3000.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1754.920 2996.000 1755.200 3000.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1817.940 2996.000 1818.220 3000.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1880.960 2996.000 1881.240 3000.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 176.200 2996.000 176.480 3000.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1944.440 2996.000 1944.720 3000.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2007.460 2996.000 2007.740 3000.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2070.480 2996.000 2070.760 3000.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2133.960 2996.000 2134.240 3000.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2196.980 2996.000 2197.260 3000.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2260.000 2996.000 2260.280 3000.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2323.020 2996.000 2323.300 3000.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2386.500 2996.000 2386.780 3000.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 239.220 2996.000 239.500 3000.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 302.240 2996.000 302.520 3000.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 365.260 2996.000 365.540 3000.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 428.740 2996.000 429.020 3000.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 491.760 2996.000 492.040 3000.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 554.780 2996.000 555.060 3000.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 618.260 2996.000 618.540 3000.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 518.900 0.000 519.180 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.140 0.000 1988.420 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2002.860 0.000 2003.140 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2017.580 0.000 2017.860 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2032.300 0.000 2032.580 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2047.020 0.000 2047.300 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2061.740 0.000 2062.020 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2076.460 0.000 2076.740 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2091.180 0.000 2091.460 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2105.900 0.000 2106.180 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2120.620 0.000 2120.900 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 665.640 0.000 665.920 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2135.340 0.000 2135.620 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2150.060 0.000 2150.340 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2164.320 0.000 2164.600 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2179.040 0.000 2179.320 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2193.760 0.000 2194.040 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2208.480 0.000 2208.760 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2223.200 0.000 2223.480 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2237.920 0.000 2238.200 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2252.640 0.000 2252.920 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2267.360 0.000 2267.640 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.360 0.000 680.640 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2282.080 0.000 2282.360 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2296.800 0.000 2297.080 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2311.520 0.000 2311.800 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2326.240 0.000 2326.520 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2340.960 0.000 2341.240 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2355.680 0.000 2355.960 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2370.400 0.000 2370.680 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2385.120 0.000 2385.400 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 695.080 0.000 695.360 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 709.800 0.000 710.080 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 724.520 0.000 724.800 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 739.240 0.000 739.520 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 753.960 0.000 754.240 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 768.680 0.000 768.960 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.400 0.000 783.680 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 798.120 0.000 798.400 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 533.620 0.000 533.900 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 812.840 0.000 813.120 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 827.560 0.000 827.840 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 842.280 0.000 842.560 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 857.000 0.000 857.280 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 871.720 0.000 872.000 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 886.440 0.000 886.720 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 901.160 0.000 901.440 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 915.420 0.000 915.700 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.140 0.000 930.420 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 944.860 0.000 945.140 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 548.340 0.000 548.620 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 959.580 0.000 959.860 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 974.300 0.000 974.580 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.020 0.000 989.300 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1003.740 0.000 1004.020 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1018.460 0.000 1018.740 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1033.180 0.000 1033.460 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1047.900 0.000 1048.180 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1062.620 0.000 1062.900 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1077.340 0.000 1077.620 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1092.060 0.000 1092.340 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 563.060 0.000 563.340 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1106.780 0.000 1107.060 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1121.500 0.000 1121.780 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1136.220 0.000 1136.500 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.940 0.000 1151.220 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1165.200 0.000 1165.480 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.920 0.000 1180.200 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1194.640 0.000 1194.920 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1209.360 0.000 1209.640 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1224.080 0.000 1224.360 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1238.800 0.000 1239.080 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 577.780 0.000 578.060 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1253.520 0.000 1253.800 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1268.240 0.000 1268.520 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1282.960 0.000 1283.240 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1297.680 0.000 1297.960 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1312.400 0.000 1312.680 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1327.120 0.000 1327.400 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1341.840 0.000 1342.120 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1356.560 0.000 1356.840 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1371.280 0.000 1371.560 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1386.000 0.000 1386.280 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 592.500 0.000 592.780 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.720 0.000 1401.000 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1414.980 0.000 1415.260 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.700 0.000 1429.980 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1444.420 0.000 1444.700 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1459.140 0.000 1459.420 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1473.860 0.000 1474.140 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1488.580 0.000 1488.860 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1503.300 0.000 1503.580 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.020 0.000 1518.300 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1532.740 0.000 1533.020 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 607.220 0.000 607.500 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1547.460 0.000 1547.740 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1562.180 0.000 1562.460 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1576.900 0.000 1577.180 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1591.620 0.000 1591.900 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1606.340 0.000 1606.620 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1621.060 0.000 1621.340 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1635.780 0.000 1636.060 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1650.500 0.000 1650.780 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1664.760 0.000 1665.040 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.480 0.000 1679.760 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 621.940 0.000 622.220 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1694.200 0.000 1694.480 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1708.920 0.000 1709.200 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1723.640 0.000 1723.920 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1738.360 0.000 1738.640 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1753.080 0.000 1753.360 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1767.800 0.000 1768.080 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1782.520 0.000 1782.800 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1797.240 0.000 1797.520 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1811.960 0.000 1812.240 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1826.680 0.000 1826.960 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 636.660 0.000 636.940 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1841.400 0.000 1841.680 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1856.120 0.000 1856.400 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1870.840 0.000 1871.120 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1885.560 0.000 1885.840 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1900.280 0.000 1900.560 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1914.540 0.000 1914.820 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.260 0.000 1929.540 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1943.980 0.000 1944.260 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1958.700 0.000 1958.980 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1973.420 0.000 1973.700 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 651.380 0.000 651.660 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 523.960 0.000 524.240 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1993.200 0.000 1993.480 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2007.920 0.000 2008.200 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2022.640 0.000 2022.920 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2037.360 0.000 2037.640 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2052.080 0.000 2052.360 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.800 0.000 2067.080 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2081.060 0.000 2081.340 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2095.780 0.000 2096.060 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2110.500 0.000 2110.780 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2125.220 0.000 2125.500 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 670.700 0.000 670.980 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2139.940 0.000 2140.220 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2154.660 0.000 2154.940 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2169.380 0.000 2169.660 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2184.100 0.000 2184.380 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2198.820 0.000 2199.100 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2213.540 0.000 2213.820 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2228.260 0.000 2228.540 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2242.980 0.000 2243.260 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2257.700 0.000 2257.980 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2272.420 0.000 2272.700 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 685.420 0.000 685.700 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2287.140 0.000 2287.420 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2301.860 0.000 2302.140 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.580 0.000 2316.860 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2330.840 0.000 2331.120 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2345.560 0.000 2345.840 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2360.280 0.000 2360.560 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2375.000 0.000 2375.280 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2389.720 0.000 2390.000 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 700.140 0.000 700.420 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 714.860 0.000 715.140 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 729.580 0.000 729.860 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 744.300 0.000 744.580 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 759.020 0.000 759.300 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 773.740 0.000 774.020 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 788.460 0.000 788.740 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 803.180 0.000 803.460 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 538.680 0.000 538.960 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.900 0.000 818.180 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 832.160 0.000 832.440 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 846.880 0.000 847.160 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 861.600 0.000 861.880 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 876.320 0.000 876.600 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 891.040 0.000 891.320 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 905.760 0.000 906.040 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 920.480 0.000 920.760 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 935.200 0.000 935.480 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 949.920 0.000 950.200 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 553.400 0.000 553.680 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 964.640 0.000 964.920 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 979.360 0.000 979.640 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 994.080 0.000 994.360 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1008.800 0.000 1009.080 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1023.520 0.000 1023.800 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1038.240 0.000 1038.520 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1052.960 0.000 1053.240 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.680 0.000 1067.960 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1081.940 0.000 1082.220 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1096.660 0.000 1096.940 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 568.120 0.000 568.400 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1111.380 0.000 1111.660 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1126.100 0.000 1126.380 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1140.820 0.000 1141.100 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1155.540 0.000 1155.820 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1170.260 0.000 1170.540 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1184.980 0.000 1185.260 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1199.700 0.000 1199.980 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1214.420 0.000 1214.700 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1229.140 0.000 1229.420 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1243.860 0.000 1244.140 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 582.380 0.000 582.660 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1258.580 0.000 1258.860 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1273.300 0.000 1273.580 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1288.020 0.000 1288.300 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1302.740 0.000 1303.020 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1317.460 0.000 1317.740 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1331.720 0.000 1332.000 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1346.440 0.000 1346.720 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1361.160 0.000 1361.440 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1375.880 0.000 1376.160 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1390.600 0.000 1390.880 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 597.100 0.000 597.380 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1405.320 0.000 1405.600 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1420.040 0.000 1420.320 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1434.760 0.000 1435.040 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1449.480 0.000 1449.760 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1464.200 0.000 1464.480 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1478.920 0.000 1479.200 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1493.640 0.000 1493.920 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1508.360 0.000 1508.640 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1523.080 0.000 1523.360 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1537.800 0.000 1538.080 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 611.820 0.000 612.100 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1552.520 0.000 1552.800 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1567.240 0.000 1567.520 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1581.500 0.000 1581.780 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1596.220 0.000 1596.500 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1610.940 0.000 1611.220 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1625.660 0.000 1625.940 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1640.380 0.000 1640.660 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1655.100 0.000 1655.380 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1669.820 0.000 1670.100 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1684.540 0.000 1684.820 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 626.540 0.000 626.820 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1699.260 0.000 1699.540 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1713.980 0.000 1714.260 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1728.700 0.000 1728.980 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.420 0.000 1743.700 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1758.140 0.000 1758.420 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1772.860 0.000 1773.140 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1787.580 0.000 1787.860 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1802.300 0.000 1802.580 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1817.020 0.000 1817.300 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1831.280 0.000 1831.560 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 641.260 0.000 641.540 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1846.000 0.000 1846.280 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1860.720 0.000 1861.000 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1875.440 0.000 1875.720 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1890.160 0.000 1890.440 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1904.880 0.000 1905.160 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1919.600 0.000 1919.880 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1934.320 0.000 1934.600 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1949.040 0.000 1949.320 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1963.760 0.000 1964.040 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1978.480 0.000 1978.760 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 655.980 0.000 656.260 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 528.560 0.000 528.840 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1997.800 0.000 1998.080 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2012.520 0.000 2012.800 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2027.240 0.000 2027.520 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2041.960 0.000 2042.240 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2056.680 0.000 2056.960 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2071.400 0.000 2071.680 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2086.120 0.000 2086.400 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2100.840 0.000 2101.120 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2115.560 0.000 2115.840 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2130.280 0.000 2130.560 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 675.760 0.000 676.040 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2145.000 0.000 2145.280 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2159.720 0.000 2160.000 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2174.440 0.000 2174.720 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2189.160 0.000 2189.440 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2203.880 0.000 2204.160 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2218.600 0.000 2218.880 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2233.320 0.000 2233.600 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2247.580 0.000 2247.860 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2262.300 0.000 2262.580 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2277.020 0.000 2277.300 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 690.480 0.000 690.760 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2291.740 0.000 2292.020 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2306.460 0.000 2306.740 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2321.180 0.000 2321.460 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2335.900 0.000 2336.180 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2350.620 0.000 2350.900 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2365.340 0.000 2365.620 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2380.060 0.000 2380.340 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2394.780 0.000 2395.060 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 705.200 0.000 705.480 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 719.920 0.000 720.200 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.640 0.000 734.920 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 748.900 0.000 749.180 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 763.620 0.000 763.900 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 778.340 0.000 778.620 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.060 0.000 793.340 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 807.780 0.000 808.060 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.280 0.000 543.560 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 822.500 0.000 822.780 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 837.220 0.000 837.500 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.940 0.000 852.220 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 866.660 0.000 866.940 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 881.380 0.000 881.660 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 896.100 0.000 896.380 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 910.820 0.000 911.100 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 925.540 0.000 925.820 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 940.260 0.000 940.540 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 954.980 0.000 955.260 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 558.000 0.000 558.280 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 969.700 0.000 969.980 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 984.420 0.000 984.700 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 998.680 0.000 998.960 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1013.400 0.000 1013.680 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1028.120 0.000 1028.400 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1042.840 0.000 1043.120 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1057.560 0.000 1057.840 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1072.280 0.000 1072.560 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1087.000 0.000 1087.280 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1101.720 0.000 1102.000 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 572.720 0.000 573.000 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1116.440 0.000 1116.720 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1131.160 0.000 1131.440 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1145.880 0.000 1146.160 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1160.600 0.000 1160.880 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.320 0.000 1175.600 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1190.040 0.000 1190.320 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1204.760 0.000 1205.040 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1219.480 0.000 1219.760 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1234.200 0.000 1234.480 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1248.460 0.000 1248.740 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.440 0.000 587.720 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1263.180 0.000 1263.460 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1277.900 0.000 1278.180 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1292.620 0.000 1292.900 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1307.340 0.000 1307.620 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.060 0.000 1322.340 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1336.780 0.000 1337.060 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1351.500 0.000 1351.780 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1366.220 0.000 1366.500 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1380.940 0.000 1381.220 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1395.660 0.000 1395.940 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 602.160 0.000 602.440 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1410.380 0.000 1410.660 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1425.100 0.000 1425.380 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1439.820 0.000 1440.100 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1454.540 0.000 1454.820 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1469.260 0.000 1469.540 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.980 0.000 1484.260 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1498.240 0.000 1498.520 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1512.960 0.000 1513.240 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1527.680 0.000 1527.960 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.400 0.000 1542.680 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 616.880 0.000 617.160 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1557.120 0.000 1557.400 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1571.840 0.000 1572.120 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1586.560 0.000 1586.840 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1601.280 0.000 1601.560 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1616.000 0.000 1616.280 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1630.720 0.000 1631.000 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1645.440 0.000 1645.720 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1660.160 0.000 1660.440 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1674.880 0.000 1675.160 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1689.600 0.000 1689.880 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 631.600 0.000 631.880 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1704.320 0.000 1704.600 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1719.040 0.000 1719.320 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.760 0.000 1734.040 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1748.020 0.000 1748.300 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1762.740 0.000 1763.020 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1777.460 0.000 1777.740 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.180 0.000 1792.460 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1806.900 0.000 1807.180 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1821.620 0.000 1821.900 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1836.340 0.000 1836.620 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 646.320 0.000 646.600 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1851.060 0.000 1851.340 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1865.780 0.000 1866.060 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1880.500 0.000 1880.780 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1895.220 0.000 1895.500 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1909.940 0.000 1910.220 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1924.660 0.000 1924.940 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1939.380 0.000 1939.660 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1954.100 0.000 1954.380 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1968.820 0.000 1969.100 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.540 0.000 1983.820 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 661.040 0.000 661.320 4.000 ;
    END
  END la_oen[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.020 0.000 0.300 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.620 0.000 4.900 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 9.680 0.000 9.960 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.000 0.000 29.280 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 195.520 0.000 195.800 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.240 0.000 210.520 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.960 0.000 225.240 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 239.680 0.000 239.960 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.400 0.000 254.680 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 269.120 0.000 269.400 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 283.840 0.000 284.120 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 298.560 0.000 298.840 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 313.280 0.000 313.560 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 328.000 0.000 328.280 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.780 0.000 49.060 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 342.720 0.000 343.000 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.440 0.000 357.720 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 372.160 0.000 372.440 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 386.880 0.000 387.160 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.600 0.000 401.880 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 415.860 0.000 416.140 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 430.580 0.000 430.860 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 445.300 0.000 445.580 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.020 0.000 460.300 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 474.740 0.000 475.020 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.560 0.000 68.840 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 489.460 0.000 489.740 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 504.180 0.000 504.460 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.880 0.000 88.160 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 107.660 0.000 107.940 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 122.380 0.000 122.660 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.100 0.000 137.380 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.820 0.000 152.100 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.080 0.000 166.360 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.800 0.000 181.080 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.280 0.000 14.560 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.060 0.000 34.340 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 200.580 0.000 200.860 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 215.300 0.000 215.580 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 230.020 0.000 230.300 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 244.740 0.000 245.020 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 259.460 0.000 259.740 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 274.180 0.000 274.460 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.900 0.000 289.180 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 303.620 0.000 303.900 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 318.340 0.000 318.620 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 332.600 0.000 332.880 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.840 0.000 54.120 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.320 0.000 347.600 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 362.040 0.000 362.320 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 376.760 0.000 377.040 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 391.480 0.000 391.760 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 406.200 0.000 406.480 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 420.920 0.000 421.200 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 435.640 0.000 435.920 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 450.360 0.000 450.640 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 465.080 0.000 465.360 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 479.800 0.000 480.080 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.160 0.000 73.440 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 494.520 0.000 494.800 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 509.240 0.000 509.520 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.940 0.000 93.220 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.260 0.000 112.540 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.980 0.000 127.260 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.700 0.000 141.980 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 156.420 0.000 156.700 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 171.140 0.000 171.420 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.860 0.000 186.140 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.120 0.000 39.400 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 205.640 0.000 205.920 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 220.360 0.000 220.640 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 235.080 0.000 235.360 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 249.340 0.000 249.620 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 264.060 0.000 264.340 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 278.780 0.000 279.060 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 293.500 0.000 293.780 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 308.220 0.000 308.500 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 322.940 0.000 323.220 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 337.660 0.000 337.940 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.440 0.000 58.720 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 352.380 0.000 352.660 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 367.100 0.000 367.380 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 381.820 0.000 382.100 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 396.540 0.000 396.820 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 411.260 0.000 411.540 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 425.980 0.000 426.260 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 440.700 0.000 440.980 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 455.420 0.000 455.700 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 470.140 0.000 470.420 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.860 0.000 485.140 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.220 0.000 78.500 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 499.120 0.000 499.400 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 513.840 0.000 514.120 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.540 0.000 97.820 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.320 0.000 117.600 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.040 0.000 132.320 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 146.760 0.000 147.040 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 161.480 0.000 161.760 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 176.200 0.000 176.480 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.920 0.000 191.200 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.720 0.000 44.000 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.500 0.000 63.780 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.820 0.000 83.100 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 102.600 0.000 102.880 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.340 0.000 19.620 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.400 0.000 24.680 4.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.670 10.640 20.270 2986.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.470 10.640 97.070 2986.800 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 3.150 10.795 2391.930 2986.645 ;
      LAYER met1 ;
        RECT 0.000 4.460 2391.930 2992.300 ;
      LAYER met2 ;
        RECT 0.030 2995.720 7.560 2996.000 ;
        RECT 8.400 2995.720 28.260 2996.000 ;
        RECT 29.100 2995.720 49.420 2996.000 ;
        RECT 50.260 2995.720 70.580 2996.000 ;
        RECT 71.420 2995.720 91.740 2996.000 ;
        RECT 92.580 2995.720 112.440 2996.000 ;
        RECT 113.280 2995.720 133.600 2996.000 ;
        RECT 134.440 2995.720 154.760 2996.000 ;
        RECT 155.600 2995.720 175.920 2996.000 ;
        RECT 176.760 2995.720 196.620 2996.000 ;
        RECT 197.460 2995.720 217.780 2996.000 ;
        RECT 218.620 2995.720 238.940 2996.000 ;
        RECT 239.780 2995.720 260.100 2996.000 ;
        RECT 260.940 2995.720 280.800 2996.000 ;
        RECT 281.640 2995.720 301.960 2996.000 ;
        RECT 302.800 2995.720 323.120 2996.000 ;
        RECT 323.960 2995.720 344.280 2996.000 ;
        RECT 345.120 2995.720 364.980 2996.000 ;
        RECT 365.820 2995.720 386.140 2996.000 ;
        RECT 386.980 2995.720 407.300 2996.000 ;
        RECT 408.140 2995.720 428.460 2996.000 ;
        RECT 429.300 2995.720 449.620 2996.000 ;
        RECT 450.460 2995.720 470.320 2996.000 ;
        RECT 471.160 2995.720 491.480 2996.000 ;
        RECT 492.320 2995.720 512.640 2996.000 ;
        RECT 513.480 2995.720 533.800 2996.000 ;
        RECT 534.640 2995.720 554.500 2996.000 ;
        RECT 555.340 2995.720 575.660 2996.000 ;
        RECT 576.500 2995.720 596.820 2996.000 ;
        RECT 597.660 2995.720 617.980 2996.000 ;
        RECT 618.820 2995.720 638.680 2996.000 ;
        RECT 639.520 2995.720 659.840 2996.000 ;
        RECT 660.680 2995.720 681.000 2996.000 ;
        RECT 681.840 2995.720 702.160 2996.000 ;
        RECT 703.000 2995.720 722.860 2996.000 ;
        RECT 723.700 2995.720 744.020 2996.000 ;
        RECT 744.860 2995.720 765.180 2996.000 ;
        RECT 766.020 2995.720 786.340 2996.000 ;
        RECT 787.180 2995.720 807.500 2996.000 ;
        RECT 808.340 2995.720 828.200 2996.000 ;
        RECT 829.040 2995.720 849.360 2996.000 ;
        RECT 850.200 2995.720 870.520 2996.000 ;
        RECT 871.360 2995.720 891.680 2996.000 ;
        RECT 892.520 2995.720 912.380 2996.000 ;
        RECT 913.220 2995.720 933.540 2996.000 ;
        RECT 934.380 2995.720 954.700 2996.000 ;
        RECT 955.540 2995.720 975.860 2996.000 ;
        RECT 976.700 2995.720 996.560 2996.000 ;
        RECT 997.400 2995.720 1017.720 2996.000 ;
        RECT 1018.560 2995.720 1038.880 2996.000 ;
        RECT 1039.720 2995.720 1060.040 2996.000 ;
        RECT 1060.880 2995.720 1080.740 2996.000 ;
        RECT 1081.580 2995.720 1101.900 2996.000 ;
        RECT 1102.740 2995.720 1123.060 2996.000 ;
        RECT 1123.900 2995.720 1144.220 2996.000 ;
        RECT 1145.060 2995.720 1164.920 2996.000 ;
        RECT 1165.760 2995.720 1186.080 2996.000 ;
        RECT 1186.920 2995.720 1207.240 2996.000 ;
        RECT 1208.080 2995.720 1228.400 2996.000 ;
        RECT 1229.240 2995.720 1249.560 2996.000 ;
        RECT 1250.400 2995.720 1270.260 2996.000 ;
        RECT 1271.100 2995.720 1291.420 2996.000 ;
        RECT 1292.260 2995.720 1312.580 2996.000 ;
        RECT 1313.420 2995.720 1333.740 2996.000 ;
        RECT 1334.580 2995.720 1354.440 2996.000 ;
        RECT 1355.280 2995.720 1375.600 2996.000 ;
        RECT 1376.440 2995.720 1396.760 2996.000 ;
        RECT 1397.600 2995.720 1417.920 2996.000 ;
        RECT 1418.760 2995.720 1438.620 2996.000 ;
        RECT 1439.460 2995.720 1459.780 2996.000 ;
        RECT 1460.620 2995.720 1480.940 2996.000 ;
        RECT 1481.780 2995.720 1502.100 2996.000 ;
        RECT 1502.940 2995.720 1522.800 2996.000 ;
        RECT 1523.640 2995.720 1543.960 2996.000 ;
        RECT 1544.800 2995.720 1565.120 2996.000 ;
        RECT 1565.960 2995.720 1586.280 2996.000 ;
        RECT 1587.120 2995.720 1607.440 2996.000 ;
        RECT 1608.280 2995.720 1628.140 2996.000 ;
        RECT 1628.980 2995.720 1649.300 2996.000 ;
        RECT 1650.140 2995.720 1670.460 2996.000 ;
        RECT 1671.300 2995.720 1691.620 2996.000 ;
        RECT 1692.460 2995.720 1712.320 2996.000 ;
        RECT 1713.160 2995.720 1733.480 2996.000 ;
        RECT 1734.320 2995.720 1754.640 2996.000 ;
        RECT 1755.480 2995.720 1775.800 2996.000 ;
        RECT 1776.640 2995.720 1796.500 2996.000 ;
        RECT 1797.340 2995.720 1817.660 2996.000 ;
        RECT 1818.500 2995.720 1838.820 2996.000 ;
        RECT 1839.660 2995.720 1859.980 2996.000 ;
        RECT 1860.820 2995.720 1880.680 2996.000 ;
        RECT 1881.520 2995.720 1901.840 2996.000 ;
        RECT 1902.680 2995.720 1923.000 2996.000 ;
        RECT 1923.840 2995.720 1944.160 2996.000 ;
        RECT 1945.000 2995.720 1964.860 2996.000 ;
        RECT 1965.700 2995.720 1986.020 2996.000 ;
        RECT 1986.860 2995.720 2007.180 2996.000 ;
        RECT 2008.020 2995.720 2028.340 2996.000 ;
        RECT 2029.180 2995.720 2049.500 2996.000 ;
        RECT 2050.340 2995.720 2070.200 2996.000 ;
        RECT 2071.040 2995.720 2091.360 2996.000 ;
        RECT 2092.200 2995.720 2112.520 2996.000 ;
        RECT 2113.360 2995.720 2133.680 2996.000 ;
        RECT 2134.520 2995.720 2154.380 2996.000 ;
        RECT 2155.220 2995.720 2175.540 2996.000 ;
        RECT 2176.380 2995.720 2196.700 2996.000 ;
        RECT 2197.540 2995.720 2217.860 2996.000 ;
        RECT 2218.700 2995.720 2238.560 2996.000 ;
        RECT 2239.400 2995.720 2259.720 2996.000 ;
        RECT 2260.560 2995.720 2280.880 2996.000 ;
        RECT 2281.720 2995.720 2302.040 2996.000 ;
        RECT 2302.880 2995.720 2322.740 2996.000 ;
        RECT 2323.580 2995.720 2343.900 2996.000 ;
        RECT 2344.740 2995.720 2365.060 2996.000 ;
        RECT 2365.900 2995.720 2386.220 2996.000 ;
        RECT 2387.060 2995.720 2389.990 2996.000 ;
        RECT 0.030 4.280 2389.990 2995.720 ;
        RECT 0.580 4.000 4.340 4.280 ;
        RECT 5.180 4.000 9.400 4.280 ;
        RECT 10.240 4.000 14.000 4.280 ;
        RECT 14.840 4.000 19.060 4.280 ;
        RECT 19.900 4.000 24.120 4.280 ;
        RECT 24.960 4.000 28.720 4.280 ;
        RECT 29.560 4.000 33.780 4.280 ;
        RECT 34.620 4.000 38.840 4.280 ;
        RECT 39.680 4.000 43.440 4.280 ;
        RECT 44.280 4.000 48.500 4.280 ;
        RECT 49.340 4.000 53.560 4.280 ;
        RECT 54.400 4.000 58.160 4.280 ;
        RECT 59.000 4.000 63.220 4.280 ;
        RECT 64.060 4.000 68.280 4.280 ;
        RECT 69.120 4.000 72.880 4.280 ;
        RECT 73.720 4.000 77.940 4.280 ;
        RECT 78.780 4.000 82.540 4.280 ;
        RECT 83.380 4.000 87.600 4.280 ;
        RECT 88.440 4.000 92.660 4.280 ;
        RECT 93.500 4.000 97.260 4.280 ;
        RECT 98.100 4.000 102.320 4.280 ;
        RECT 103.160 4.000 107.380 4.280 ;
        RECT 108.220 4.000 111.980 4.280 ;
        RECT 112.820 4.000 117.040 4.280 ;
        RECT 117.880 4.000 122.100 4.280 ;
        RECT 122.940 4.000 126.700 4.280 ;
        RECT 127.540 4.000 131.760 4.280 ;
        RECT 132.600 4.000 136.820 4.280 ;
        RECT 137.660 4.000 141.420 4.280 ;
        RECT 142.260 4.000 146.480 4.280 ;
        RECT 147.320 4.000 151.540 4.280 ;
        RECT 152.380 4.000 156.140 4.280 ;
        RECT 156.980 4.000 161.200 4.280 ;
        RECT 162.040 4.000 165.800 4.280 ;
        RECT 166.640 4.000 170.860 4.280 ;
        RECT 171.700 4.000 175.920 4.280 ;
        RECT 176.760 4.000 180.520 4.280 ;
        RECT 181.360 4.000 185.580 4.280 ;
        RECT 186.420 4.000 190.640 4.280 ;
        RECT 191.480 4.000 195.240 4.280 ;
        RECT 196.080 4.000 200.300 4.280 ;
        RECT 201.140 4.000 205.360 4.280 ;
        RECT 206.200 4.000 209.960 4.280 ;
        RECT 210.800 4.000 215.020 4.280 ;
        RECT 215.860 4.000 220.080 4.280 ;
        RECT 220.920 4.000 224.680 4.280 ;
        RECT 225.520 4.000 229.740 4.280 ;
        RECT 230.580 4.000 234.800 4.280 ;
        RECT 235.640 4.000 239.400 4.280 ;
        RECT 240.240 4.000 244.460 4.280 ;
        RECT 245.300 4.000 249.060 4.280 ;
        RECT 249.900 4.000 254.120 4.280 ;
        RECT 254.960 4.000 259.180 4.280 ;
        RECT 260.020 4.000 263.780 4.280 ;
        RECT 264.620 4.000 268.840 4.280 ;
        RECT 269.680 4.000 273.900 4.280 ;
        RECT 274.740 4.000 278.500 4.280 ;
        RECT 279.340 4.000 283.560 4.280 ;
        RECT 284.400 4.000 288.620 4.280 ;
        RECT 289.460 4.000 293.220 4.280 ;
        RECT 294.060 4.000 298.280 4.280 ;
        RECT 299.120 4.000 303.340 4.280 ;
        RECT 304.180 4.000 307.940 4.280 ;
        RECT 308.780 4.000 313.000 4.280 ;
        RECT 313.840 4.000 318.060 4.280 ;
        RECT 318.900 4.000 322.660 4.280 ;
        RECT 323.500 4.000 327.720 4.280 ;
        RECT 328.560 4.000 332.320 4.280 ;
        RECT 333.160 4.000 337.380 4.280 ;
        RECT 338.220 4.000 342.440 4.280 ;
        RECT 343.280 4.000 347.040 4.280 ;
        RECT 347.880 4.000 352.100 4.280 ;
        RECT 352.940 4.000 357.160 4.280 ;
        RECT 358.000 4.000 361.760 4.280 ;
        RECT 362.600 4.000 366.820 4.280 ;
        RECT 367.660 4.000 371.880 4.280 ;
        RECT 372.720 4.000 376.480 4.280 ;
        RECT 377.320 4.000 381.540 4.280 ;
        RECT 382.380 4.000 386.600 4.280 ;
        RECT 387.440 4.000 391.200 4.280 ;
        RECT 392.040 4.000 396.260 4.280 ;
        RECT 397.100 4.000 401.320 4.280 ;
        RECT 402.160 4.000 405.920 4.280 ;
        RECT 406.760 4.000 410.980 4.280 ;
        RECT 411.820 4.000 415.580 4.280 ;
        RECT 416.420 4.000 420.640 4.280 ;
        RECT 421.480 4.000 425.700 4.280 ;
        RECT 426.540 4.000 430.300 4.280 ;
        RECT 431.140 4.000 435.360 4.280 ;
        RECT 436.200 4.000 440.420 4.280 ;
        RECT 441.260 4.000 445.020 4.280 ;
        RECT 445.860 4.000 450.080 4.280 ;
        RECT 450.920 4.000 455.140 4.280 ;
        RECT 455.980 4.000 459.740 4.280 ;
        RECT 460.580 4.000 464.800 4.280 ;
        RECT 465.640 4.000 469.860 4.280 ;
        RECT 470.700 4.000 474.460 4.280 ;
        RECT 475.300 4.000 479.520 4.280 ;
        RECT 480.360 4.000 484.580 4.280 ;
        RECT 485.420 4.000 489.180 4.280 ;
        RECT 490.020 4.000 494.240 4.280 ;
        RECT 495.080 4.000 498.840 4.280 ;
        RECT 499.680 4.000 503.900 4.280 ;
        RECT 504.740 4.000 508.960 4.280 ;
        RECT 509.800 4.000 513.560 4.280 ;
        RECT 514.400 4.000 518.620 4.280 ;
        RECT 519.460 4.000 523.680 4.280 ;
        RECT 524.520 4.000 528.280 4.280 ;
        RECT 529.120 4.000 533.340 4.280 ;
        RECT 534.180 4.000 538.400 4.280 ;
        RECT 539.240 4.000 543.000 4.280 ;
        RECT 543.840 4.000 548.060 4.280 ;
        RECT 548.900 4.000 553.120 4.280 ;
        RECT 553.960 4.000 557.720 4.280 ;
        RECT 558.560 4.000 562.780 4.280 ;
        RECT 563.620 4.000 567.840 4.280 ;
        RECT 568.680 4.000 572.440 4.280 ;
        RECT 573.280 4.000 577.500 4.280 ;
        RECT 578.340 4.000 582.100 4.280 ;
        RECT 582.940 4.000 587.160 4.280 ;
        RECT 588.000 4.000 592.220 4.280 ;
        RECT 593.060 4.000 596.820 4.280 ;
        RECT 597.660 4.000 601.880 4.280 ;
        RECT 602.720 4.000 606.940 4.280 ;
        RECT 607.780 4.000 611.540 4.280 ;
        RECT 612.380 4.000 616.600 4.280 ;
        RECT 617.440 4.000 621.660 4.280 ;
        RECT 622.500 4.000 626.260 4.280 ;
        RECT 627.100 4.000 631.320 4.280 ;
        RECT 632.160 4.000 636.380 4.280 ;
        RECT 637.220 4.000 640.980 4.280 ;
        RECT 641.820 4.000 646.040 4.280 ;
        RECT 646.880 4.000 651.100 4.280 ;
        RECT 651.940 4.000 655.700 4.280 ;
        RECT 656.540 4.000 660.760 4.280 ;
        RECT 661.600 4.000 665.360 4.280 ;
        RECT 666.200 4.000 670.420 4.280 ;
        RECT 671.260 4.000 675.480 4.280 ;
        RECT 676.320 4.000 680.080 4.280 ;
        RECT 680.920 4.000 685.140 4.280 ;
        RECT 685.980 4.000 690.200 4.280 ;
        RECT 691.040 4.000 694.800 4.280 ;
        RECT 695.640 4.000 699.860 4.280 ;
        RECT 700.700 4.000 704.920 4.280 ;
        RECT 705.760 4.000 709.520 4.280 ;
        RECT 710.360 4.000 714.580 4.280 ;
        RECT 715.420 4.000 719.640 4.280 ;
        RECT 720.480 4.000 724.240 4.280 ;
        RECT 725.080 4.000 729.300 4.280 ;
        RECT 730.140 4.000 734.360 4.280 ;
        RECT 735.200 4.000 738.960 4.280 ;
        RECT 739.800 4.000 744.020 4.280 ;
        RECT 744.860 4.000 748.620 4.280 ;
        RECT 749.460 4.000 753.680 4.280 ;
        RECT 754.520 4.000 758.740 4.280 ;
        RECT 759.580 4.000 763.340 4.280 ;
        RECT 764.180 4.000 768.400 4.280 ;
        RECT 769.240 4.000 773.460 4.280 ;
        RECT 774.300 4.000 778.060 4.280 ;
        RECT 778.900 4.000 783.120 4.280 ;
        RECT 783.960 4.000 788.180 4.280 ;
        RECT 789.020 4.000 792.780 4.280 ;
        RECT 793.620 4.000 797.840 4.280 ;
        RECT 798.680 4.000 802.900 4.280 ;
        RECT 803.740 4.000 807.500 4.280 ;
        RECT 808.340 4.000 812.560 4.280 ;
        RECT 813.400 4.000 817.620 4.280 ;
        RECT 818.460 4.000 822.220 4.280 ;
        RECT 823.060 4.000 827.280 4.280 ;
        RECT 828.120 4.000 831.880 4.280 ;
        RECT 832.720 4.000 836.940 4.280 ;
        RECT 837.780 4.000 842.000 4.280 ;
        RECT 842.840 4.000 846.600 4.280 ;
        RECT 847.440 4.000 851.660 4.280 ;
        RECT 852.500 4.000 856.720 4.280 ;
        RECT 857.560 4.000 861.320 4.280 ;
        RECT 862.160 4.000 866.380 4.280 ;
        RECT 867.220 4.000 871.440 4.280 ;
        RECT 872.280 4.000 876.040 4.280 ;
        RECT 876.880 4.000 881.100 4.280 ;
        RECT 881.940 4.000 886.160 4.280 ;
        RECT 887.000 4.000 890.760 4.280 ;
        RECT 891.600 4.000 895.820 4.280 ;
        RECT 896.660 4.000 900.880 4.280 ;
        RECT 901.720 4.000 905.480 4.280 ;
        RECT 906.320 4.000 910.540 4.280 ;
        RECT 911.380 4.000 915.140 4.280 ;
        RECT 915.980 4.000 920.200 4.280 ;
        RECT 921.040 4.000 925.260 4.280 ;
        RECT 926.100 4.000 929.860 4.280 ;
        RECT 930.700 4.000 934.920 4.280 ;
        RECT 935.760 4.000 939.980 4.280 ;
        RECT 940.820 4.000 944.580 4.280 ;
        RECT 945.420 4.000 949.640 4.280 ;
        RECT 950.480 4.000 954.700 4.280 ;
        RECT 955.540 4.000 959.300 4.280 ;
        RECT 960.140 4.000 964.360 4.280 ;
        RECT 965.200 4.000 969.420 4.280 ;
        RECT 970.260 4.000 974.020 4.280 ;
        RECT 974.860 4.000 979.080 4.280 ;
        RECT 979.920 4.000 984.140 4.280 ;
        RECT 984.980 4.000 988.740 4.280 ;
        RECT 989.580 4.000 993.800 4.280 ;
        RECT 994.640 4.000 998.400 4.280 ;
        RECT 999.240 4.000 1003.460 4.280 ;
        RECT 1004.300 4.000 1008.520 4.280 ;
        RECT 1009.360 4.000 1013.120 4.280 ;
        RECT 1013.960 4.000 1018.180 4.280 ;
        RECT 1019.020 4.000 1023.240 4.280 ;
        RECT 1024.080 4.000 1027.840 4.280 ;
        RECT 1028.680 4.000 1032.900 4.280 ;
        RECT 1033.740 4.000 1037.960 4.280 ;
        RECT 1038.800 4.000 1042.560 4.280 ;
        RECT 1043.400 4.000 1047.620 4.280 ;
        RECT 1048.460 4.000 1052.680 4.280 ;
        RECT 1053.520 4.000 1057.280 4.280 ;
        RECT 1058.120 4.000 1062.340 4.280 ;
        RECT 1063.180 4.000 1067.400 4.280 ;
        RECT 1068.240 4.000 1072.000 4.280 ;
        RECT 1072.840 4.000 1077.060 4.280 ;
        RECT 1077.900 4.000 1081.660 4.280 ;
        RECT 1082.500 4.000 1086.720 4.280 ;
        RECT 1087.560 4.000 1091.780 4.280 ;
        RECT 1092.620 4.000 1096.380 4.280 ;
        RECT 1097.220 4.000 1101.440 4.280 ;
        RECT 1102.280 4.000 1106.500 4.280 ;
        RECT 1107.340 4.000 1111.100 4.280 ;
        RECT 1111.940 4.000 1116.160 4.280 ;
        RECT 1117.000 4.000 1121.220 4.280 ;
        RECT 1122.060 4.000 1125.820 4.280 ;
        RECT 1126.660 4.000 1130.880 4.280 ;
        RECT 1131.720 4.000 1135.940 4.280 ;
        RECT 1136.780 4.000 1140.540 4.280 ;
        RECT 1141.380 4.000 1145.600 4.280 ;
        RECT 1146.440 4.000 1150.660 4.280 ;
        RECT 1151.500 4.000 1155.260 4.280 ;
        RECT 1156.100 4.000 1160.320 4.280 ;
        RECT 1161.160 4.000 1164.920 4.280 ;
        RECT 1165.760 4.000 1169.980 4.280 ;
        RECT 1170.820 4.000 1175.040 4.280 ;
        RECT 1175.880 4.000 1179.640 4.280 ;
        RECT 1180.480 4.000 1184.700 4.280 ;
        RECT 1185.540 4.000 1189.760 4.280 ;
        RECT 1190.600 4.000 1194.360 4.280 ;
        RECT 1195.200 4.000 1199.420 4.280 ;
        RECT 1200.260 4.000 1204.480 4.280 ;
        RECT 1205.320 4.000 1209.080 4.280 ;
        RECT 1209.920 4.000 1214.140 4.280 ;
        RECT 1214.980 4.000 1219.200 4.280 ;
        RECT 1220.040 4.000 1223.800 4.280 ;
        RECT 1224.640 4.000 1228.860 4.280 ;
        RECT 1229.700 4.000 1233.920 4.280 ;
        RECT 1234.760 4.000 1238.520 4.280 ;
        RECT 1239.360 4.000 1243.580 4.280 ;
        RECT 1244.420 4.000 1248.180 4.280 ;
        RECT 1249.020 4.000 1253.240 4.280 ;
        RECT 1254.080 4.000 1258.300 4.280 ;
        RECT 1259.140 4.000 1262.900 4.280 ;
        RECT 1263.740 4.000 1267.960 4.280 ;
        RECT 1268.800 4.000 1273.020 4.280 ;
        RECT 1273.860 4.000 1277.620 4.280 ;
        RECT 1278.460 4.000 1282.680 4.280 ;
        RECT 1283.520 4.000 1287.740 4.280 ;
        RECT 1288.580 4.000 1292.340 4.280 ;
        RECT 1293.180 4.000 1297.400 4.280 ;
        RECT 1298.240 4.000 1302.460 4.280 ;
        RECT 1303.300 4.000 1307.060 4.280 ;
        RECT 1307.900 4.000 1312.120 4.280 ;
        RECT 1312.960 4.000 1317.180 4.280 ;
        RECT 1318.020 4.000 1321.780 4.280 ;
        RECT 1322.620 4.000 1326.840 4.280 ;
        RECT 1327.680 4.000 1331.440 4.280 ;
        RECT 1332.280 4.000 1336.500 4.280 ;
        RECT 1337.340 4.000 1341.560 4.280 ;
        RECT 1342.400 4.000 1346.160 4.280 ;
        RECT 1347.000 4.000 1351.220 4.280 ;
        RECT 1352.060 4.000 1356.280 4.280 ;
        RECT 1357.120 4.000 1360.880 4.280 ;
        RECT 1361.720 4.000 1365.940 4.280 ;
        RECT 1366.780 4.000 1371.000 4.280 ;
        RECT 1371.840 4.000 1375.600 4.280 ;
        RECT 1376.440 4.000 1380.660 4.280 ;
        RECT 1381.500 4.000 1385.720 4.280 ;
        RECT 1386.560 4.000 1390.320 4.280 ;
        RECT 1391.160 4.000 1395.380 4.280 ;
        RECT 1396.220 4.000 1400.440 4.280 ;
        RECT 1401.280 4.000 1405.040 4.280 ;
        RECT 1405.880 4.000 1410.100 4.280 ;
        RECT 1410.940 4.000 1414.700 4.280 ;
        RECT 1415.540 4.000 1419.760 4.280 ;
        RECT 1420.600 4.000 1424.820 4.280 ;
        RECT 1425.660 4.000 1429.420 4.280 ;
        RECT 1430.260 4.000 1434.480 4.280 ;
        RECT 1435.320 4.000 1439.540 4.280 ;
        RECT 1440.380 4.000 1444.140 4.280 ;
        RECT 1444.980 4.000 1449.200 4.280 ;
        RECT 1450.040 4.000 1454.260 4.280 ;
        RECT 1455.100 4.000 1458.860 4.280 ;
        RECT 1459.700 4.000 1463.920 4.280 ;
        RECT 1464.760 4.000 1468.980 4.280 ;
        RECT 1469.820 4.000 1473.580 4.280 ;
        RECT 1474.420 4.000 1478.640 4.280 ;
        RECT 1479.480 4.000 1483.700 4.280 ;
        RECT 1484.540 4.000 1488.300 4.280 ;
        RECT 1489.140 4.000 1493.360 4.280 ;
        RECT 1494.200 4.000 1497.960 4.280 ;
        RECT 1498.800 4.000 1503.020 4.280 ;
        RECT 1503.860 4.000 1508.080 4.280 ;
        RECT 1508.920 4.000 1512.680 4.280 ;
        RECT 1513.520 4.000 1517.740 4.280 ;
        RECT 1518.580 4.000 1522.800 4.280 ;
        RECT 1523.640 4.000 1527.400 4.280 ;
        RECT 1528.240 4.000 1532.460 4.280 ;
        RECT 1533.300 4.000 1537.520 4.280 ;
        RECT 1538.360 4.000 1542.120 4.280 ;
        RECT 1542.960 4.000 1547.180 4.280 ;
        RECT 1548.020 4.000 1552.240 4.280 ;
        RECT 1553.080 4.000 1556.840 4.280 ;
        RECT 1557.680 4.000 1561.900 4.280 ;
        RECT 1562.740 4.000 1566.960 4.280 ;
        RECT 1567.800 4.000 1571.560 4.280 ;
        RECT 1572.400 4.000 1576.620 4.280 ;
        RECT 1577.460 4.000 1581.220 4.280 ;
        RECT 1582.060 4.000 1586.280 4.280 ;
        RECT 1587.120 4.000 1591.340 4.280 ;
        RECT 1592.180 4.000 1595.940 4.280 ;
        RECT 1596.780 4.000 1601.000 4.280 ;
        RECT 1601.840 4.000 1606.060 4.280 ;
        RECT 1606.900 4.000 1610.660 4.280 ;
        RECT 1611.500 4.000 1615.720 4.280 ;
        RECT 1616.560 4.000 1620.780 4.280 ;
        RECT 1621.620 4.000 1625.380 4.280 ;
        RECT 1626.220 4.000 1630.440 4.280 ;
        RECT 1631.280 4.000 1635.500 4.280 ;
        RECT 1636.340 4.000 1640.100 4.280 ;
        RECT 1640.940 4.000 1645.160 4.280 ;
        RECT 1646.000 4.000 1650.220 4.280 ;
        RECT 1651.060 4.000 1654.820 4.280 ;
        RECT 1655.660 4.000 1659.880 4.280 ;
        RECT 1660.720 4.000 1664.480 4.280 ;
        RECT 1665.320 4.000 1669.540 4.280 ;
        RECT 1670.380 4.000 1674.600 4.280 ;
        RECT 1675.440 4.000 1679.200 4.280 ;
        RECT 1680.040 4.000 1684.260 4.280 ;
        RECT 1685.100 4.000 1689.320 4.280 ;
        RECT 1690.160 4.000 1693.920 4.280 ;
        RECT 1694.760 4.000 1698.980 4.280 ;
        RECT 1699.820 4.000 1704.040 4.280 ;
        RECT 1704.880 4.000 1708.640 4.280 ;
        RECT 1709.480 4.000 1713.700 4.280 ;
        RECT 1714.540 4.000 1718.760 4.280 ;
        RECT 1719.600 4.000 1723.360 4.280 ;
        RECT 1724.200 4.000 1728.420 4.280 ;
        RECT 1729.260 4.000 1733.480 4.280 ;
        RECT 1734.320 4.000 1738.080 4.280 ;
        RECT 1738.920 4.000 1743.140 4.280 ;
        RECT 1743.980 4.000 1747.740 4.280 ;
        RECT 1748.580 4.000 1752.800 4.280 ;
        RECT 1753.640 4.000 1757.860 4.280 ;
        RECT 1758.700 4.000 1762.460 4.280 ;
        RECT 1763.300 4.000 1767.520 4.280 ;
        RECT 1768.360 4.000 1772.580 4.280 ;
        RECT 1773.420 4.000 1777.180 4.280 ;
        RECT 1778.020 4.000 1782.240 4.280 ;
        RECT 1783.080 4.000 1787.300 4.280 ;
        RECT 1788.140 4.000 1791.900 4.280 ;
        RECT 1792.740 4.000 1796.960 4.280 ;
        RECT 1797.800 4.000 1802.020 4.280 ;
        RECT 1802.860 4.000 1806.620 4.280 ;
        RECT 1807.460 4.000 1811.680 4.280 ;
        RECT 1812.520 4.000 1816.740 4.280 ;
        RECT 1817.580 4.000 1821.340 4.280 ;
        RECT 1822.180 4.000 1826.400 4.280 ;
        RECT 1827.240 4.000 1831.000 4.280 ;
        RECT 1831.840 4.000 1836.060 4.280 ;
        RECT 1836.900 4.000 1841.120 4.280 ;
        RECT 1841.960 4.000 1845.720 4.280 ;
        RECT 1846.560 4.000 1850.780 4.280 ;
        RECT 1851.620 4.000 1855.840 4.280 ;
        RECT 1856.680 4.000 1860.440 4.280 ;
        RECT 1861.280 4.000 1865.500 4.280 ;
        RECT 1866.340 4.000 1870.560 4.280 ;
        RECT 1871.400 4.000 1875.160 4.280 ;
        RECT 1876.000 4.000 1880.220 4.280 ;
        RECT 1881.060 4.000 1885.280 4.280 ;
        RECT 1886.120 4.000 1889.880 4.280 ;
        RECT 1890.720 4.000 1894.940 4.280 ;
        RECT 1895.780 4.000 1900.000 4.280 ;
        RECT 1900.840 4.000 1904.600 4.280 ;
        RECT 1905.440 4.000 1909.660 4.280 ;
        RECT 1910.500 4.000 1914.260 4.280 ;
        RECT 1915.100 4.000 1919.320 4.280 ;
        RECT 1920.160 4.000 1924.380 4.280 ;
        RECT 1925.220 4.000 1928.980 4.280 ;
        RECT 1929.820 4.000 1934.040 4.280 ;
        RECT 1934.880 4.000 1939.100 4.280 ;
        RECT 1939.940 4.000 1943.700 4.280 ;
        RECT 1944.540 4.000 1948.760 4.280 ;
        RECT 1949.600 4.000 1953.820 4.280 ;
        RECT 1954.660 4.000 1958.420 4.280 ;
        RECT 1959.260 4.000 1963.480 4.280 ;
        RECT 1964.320 4.000 1968.540 4.280 ;
        RECT 1969.380 4.000 1973.140 4.280 ;
        RECT 1973.980 4.000 1978.200 4.280 ;
        RECT 1979.040 4.000 1983.260 4.280 ;
        RECT 1984.100 4.000 1987.860 4.280 ;
        RECT 1988.700 4.000 1992.920 4.280 ;
        RECT 1993.760 4.000 1997.520 4.280 ;
        RECT 1998.360 4.000 2002.580 4.280 ;
        RECT 2003.420 4.000 2007.640 4.280 ;
        RECT 2008.480 4.000 2012.240 4.280 ;
        RECT 2013.080 4.000 2017.300 4.280 ;
        RECT 2018.140 4.000 2022.360 4.280 ;
        RECT 2023.200 4.000 2026.960 4.280 ;
        RECT 2027.800 4.000 2032.020 4.280 ;
        RECT 2032.860 4.000 2037.080 4.280 ;
        RECT 2037.920 4.000 2041.680 4.280 ;
        RECT 2042.520 4.000 2046.740 4.280 ;
        RECT 2047.580 4.000 2051.800 4.280 ;
        RECT 2052.640 4.000 2056.400 4.280 ;
        RECT 2057.240 4.000 2061.460 4.280 ;
        RECT 2062.300 4.000 2066.520 4.280 ;
        RECT 2067.360 4.000 2071.120 4.280 ;
        RECT 2071.960 4.000 2076.180 4.280 ;
        RECT 2077.020 4.000 2080.780 4.280 ;
        RECT 2081.620 4.000 2085.840 4.280 ;
        RECT 2086.680 4.000 2090.900 4.280 ;
        RECT 2091.740 4.000 2095.500 4.280 ;
        RECT 2096.340 4.000 2100.560 4.280 ;
        RECT 2101.400 4.000 2105.620 4.280 ;
        RECT 2106.460 4.000 2110.220 4.280 ;
        RECT 2111.060 4.000 2115.280 4.280 ;
        RECT 2116.120 4.000 2120.340 4.280 ;
        RECT 2121.180 4.000 2124.940 4.280 ;
        RECT 2125.780 4.000 2130.000 4.280 ;
        RECT 2130.840 4.000 2135.060 4.280 ;
        RECT 2135.900 4.000 2139.660 4.280 ;
        RECT 2140.500 4.000 2144.720 4.280 ;
        RECT 2145.560 4.000 2149.780 4.280 ;
        RECT 2150.620 4.000 2154.380 4.280 ;
        RECT 2155.220 4.000 2159.440 4.280 ;
        RECT 2160.280 4.000 2164.040 4.280 ;
        RECT 2164.880 4.000 2169.100 4.280 ;
        RECT 2169.940 4.000 2174.160 4.280 ;
        RECT 2175.000 4.000 2178.760 4.280 ;
        RECT 2179.600 4.000 2183.820 4.280 ;
        RECT 2184.660 4.000 2188.880 4.280 ;
        RECT 2189.720 4.000 2193.480 4.280 ;
        RECT 2194.320 4.000 2198.540 4.280 ;
        RECT 2199.380 4.000 2203.600 4.280 ;
        RECT 2204.440 4.000 2208.200 4.280 ;
        RECT 2209.040 4.000 2213.260 4.280 ;
        RECT 2214.100 4.000 2218.320 4.280 ;
        RECT 2219.160 4.000 2222.920 4.280 ;
        RECT 2223.760 4.000 2227.980 4.280 ;
        RECT 2228.820 4.000 2233.040 4.280 ;
        RECT 2233.880 4.000 2237.640 4.280 ;
        RECT 2238.480 4.000 2242.700 4.280 ;
        RECT 2243.540 4.000 2247.300 4.280 ;
        RECT 2248.140 4.000 2252.360 4.280 ;
        RECT 2253.200 4.000 2257.420 4.280 ;
        RECT 2258.260 4.000 2262.020 4.280 ;
        RECT 2262.860 4.000 2267.080 4.280 ;
        RECT 2267.920 4.000 2272.140 4.280 ;
        RECT 2272.980 4.000 2276.740 4.280 ;
        RECT 2277.580 4.000 2281.800 4.280 ;
        RECT 2282.640 4.000 2286.860 4.280 ;
        RECT 2287.700 4.000 2291.460 4.280 ;
        RECT 2292.300 4.000 2296.520 4.280 ;
        RECT 2297.360 4.000 2301.580 4.280 ;
        RECT 2302.420 4.000 2306.180 4.280 ;
        RECT 2307.020 4.000 2311.240 4.280 ;
        RECT 2312.080 4.000 2316.300 4.280 ;
        RECT 2317.140 4.000 2320.900 4.280 ;
        RECT 2321.740 4.000 2325.960 4.280 ;
        RECT 2326.800 4.000 2330.560 4.280 ;
        RECT 2331.400 4.000 2335.620 4.280 ;
        RECT 2336.460 4.000 2340.680 4.280 ;
        RECT 2341.520 4.000 2345.280 4.280 ;
        RECT 2346.120 4.000 2350.340 4.280 ;
        RECT 2351.180 4.000 2355.400 4.280 ;
        RECT 2356.240 4.000 2360.000 4.280 ;
        RECT 2360.840 4.000 2365.060 4.280 ;
        RECT 2365.900 4.000 2370.120 4.280 ;
        RECT 2370.960 4.000 2374.720 4.280 ;
        RECT 2375.560 4.000 2379.780 4.280 ;
        RECT 2380.620 4.000 2384.840 4.280 ;
        RECT 2385.680 4.000 2389.440 4.280 ;
      LAYER met3 ;
        RECT 8.735 4.255 2386.805 2987.745 ;
      LAYER met4 ;
        RECT 20.925 2987.200 2376.455 2987.745 ;
        RECT 20.925 10.640 95.070 2987.200 ;
        RECT 97.470 10.640 2376.455 2987.200 ;
  END
END user_proj_example
END LIBRARY

