magic
tech sky130A
magscale 1 2
timestamp 1607720773
<< locali >>
rect 297925 699635 297959 699805
rect 300041 699567 300075 699805
rect 305101 699567 305135 699873
rect 494069 666587 494103 676141
rect 116593 658631 116627 659277
rect 125057 658767 125091 659277
rect 129289 658835 129323 659277
rect 137569 658971 137603 659277
rect 179705 659243 179739 659345
rect 368581 659175 368615 659617
rect 369133 659175 369167 659617
rect 381277 659107 381311 659617
rect 381645 659107 381679 659617
rect 385325 659039 385359 659617
rect 410717 658903 410751 659617
rect 423229 658699 423263 659617
rect 469597 658563 469631 659617
rect 77953 57443 77987 57613
rect 81633 57443 81667 57613
rect 83565 57511 83599 57613
rect 94605 57511 94639 57613
rect 64923 57341 65015 57375
rect 64981 57239 65015 57341
rect 65165 57341 65625 57375
rect 64889 57171 64923 57205
rect 65165 57171 65199 57341
rect 64889 57137 65199 57171
rect 62957 56763 62991 56865
rect 69581 56627 69615 56661
rect 69581 56593 69765 56627
rect 79149 56559 79183 57409
rect 82553 57239 82587 57341
rect 119813 57239 119847 57341
rect 119997 57307 120031 57545
rect 91661 56967 91695 57137
rect 99389 56627 99423 56933
rect 102057 56763 102091 57069
rect 115121 56967 115155 57205
rect 120089 57171 120123 57545
rect 122573 57443 122607 57545
rect 129657 57307 129691 57477
rect 124539 57273 124781 57307
rect 119905 57137 120123 57171
rect 119905 57035 119939 57137
rect 102609 56763 102643 56933
rect 102701 56695 102735 56933
rect 115029 56695 115063 56933
rect 128829 56627 128863 56797
rect 130577 56559 130611 57545
rect 132233 57239 132267 57409
rect 100861 48331 100895 52309
rect 121561 48331 121595 51561
rect 132509 48331 132543 57477
rect 141985 57171 142019 57545
rect 147689 56831 147723 57477
rect 151737 57171 151771 57545
rect 156061 57171 156095 57749
rect 191205 57715 191239 57817
rect 191113 57579 191147 57681
rect 176669 57375 176703 57545
rect 185593 57375 185627 57477
rect 169401 56899 169435 57273
rect 142663 56661 142813 56695
rect 171149 56559 171183 56661
rect 173081 56627 173115 57341
rect 185501 56695 185535 57341
rect 191021 57035 191055 57545
rect 191297 57171 191331 57817
rect 195897 57035 195931 57477
rect 195989 48331 196023 57137
rect 211905 56763 211939 57477
rect 212825 57035 212859 57749
rect 215769 57715 215803 57885
rect 224141 57783 224175 57953
rect 224233 57783 224267 57885
rect 215861 56627 215895 57681
rect 224233 56695 224267 57273
rect 538781 57171 538815 57477
rect 334173 48331 334207 55573
rect 98561 46971 98595 48297
rect 336749 46971 336783 56457
rect 101045 31671 101079 38573
rect 128645 27727 128679 37213
rect 145021 29019 145055 35717
rect 192033 29019 192067 38573
rect 195897 29019 195931 38573
rect 338129 37315 338163 46869
rect 336749 27659 336783 37213
rect 121653 18003 121687 27557
rect 128921 19227 128955 27557
rect 192217 9707 192251 19261
rect 212549 18003 212583 27557
rect 22017 3859 22051 4097
rect 26157 3655 26191 3893
rect 35909 3723 35943 4029
rect 45477 3723 45511 4029
rect 36001 3179 36035 3621
rect 45385 3179 45419 3621
rect 45661 3315 45695 4029
rect 55229 3723 55263 4233
rect 59921 3519 59955 4165
rect 64797 3723 64831 4233
rect 96663 4165 96755 4199
rect 96721 4131 96755 4165
rect 75285 3723 75319 4097
rect 106289 4131 106323 6341
rect 84117 3791 84151 4097
rect 88993 3859 89027 4029
rect 64889 3451 64923 3689
rect 68201 3621 68385 3655
rect 68201 3519 68235 3621
rect 64889 3417 65165 3451
rect 69673 3111 69707 3689
rect 71881 3451 71915 3553
rect 71823 3417 71915 3451
rect 82829 3383 82863 3553
rect 104173 3383 104207 3485
rect 148701 3451 148735 3893
rect 156705 3587 156739 3961
rect 161489 3587 161523 3961
rect 166273 3315 166307 3689
rect 169125 3587 169159 3893
rect 191113 3587 191147 3893
rect 143273 595 143307 2805
rect 195621 595 195655 9605
rect 200773 3927 200807 4029
rect 212457 595 212491 9605
rect 333989 8347 334023 17901
rect 336749 9571 336783 17901
rect 338129 9707 338163 27557
rect 431233 3791 431267 4097
rect 433165 2839 433199 3757
rect 213469 595 213503 2805
rect 445493 2839 445527 3553
rect 446689 3179 446723 3689
rect 453773 3111 453807 3757
rect 455981 3315 456015 3553
rect 456073 3519 456107 3893
rect 456165 3519 456199 3825
rect 456257 3723 456291 4165
rect 457361 3383 457395 3689
rect 462145 3383 462179 3825
rect 465733 3485 465917 3519
rect 445585 2839 445619 3009
rect 455889 2907 455923 3281
rect 455889 2873 456165 2907
rect 460857 2839 460891 3349
rect 465733 3179 465767 3485
rect 465825 3179 465859 3417
rect 471805 3247 471839 3757
rect 476129 3451 476163 3757
rect 532893 3587 532927 3961
rect 532985 3859 533019 3961
rect 533353 3723 533387 3825
rect 533445 3723 533479 4029
rect 469321 2975 469355 3213
rect 549821 3043 549855 3349
rect 510905 2839 510939 3009
rect 552673 2975 552707 3145
rect 333621 595 333655 2805
<< viali >>
rect 305101 699873 305135 699907
rect 297925 699805 297959 699839
rect 297925 699601 297959 699635
rect 300041 699805 300075 699839
rect 300041 699533 300075 699567
rect 305101 699533 305135 699567
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 368581 659617 368615 659651
rect 179705 659345 179739 659379
rect 116593 659277 116627 659311
rect 125057 659277 125091 659311
rect 129289 659277 129323 659311
rect 137569 659277 137603 659311
rect 179705 659209 179739 659243
rect 368581 659141 368615 659175
rect 369133 659617 369167 659651
rect 369133 659141 369167 659175
rect 381277 659617 381311 659651
rect 381277 659073 381311 659107
rect 381645 659617 381679 659651
rect 381645 659073 381679 659107
rect 385325 659617 385359 659651
rect 385325 659005 385359 659039
rect 410717 659617 410751 659651
rect 137569 658937 137603 658971
rect 410717 658869 410751 658903
rect 423229 659617 423263 659651
rect 129289 658801 129323 658835
rect 125057 658733 125091 658767
rect 423229 658665 423263 658699
rect 469597 659617 469631 659651
rect 116593 658597 116627 658631
rect 469597 658529 469631 658563
rect 224141 57953 224175 57987
rect 215769 57885 215803 57919
rect 191205 57817 191239 57851
rect 156061 57749 156095 57783
rect 77953 57613 77987 57647
rect 81633 57613 81667 57647
rect 83565 57613 83599 57647
rect 83565 57477 83599 57511
rect 94605 57613 94639 57647
rect 94605 57477 94639 57511
rect 119997 57545 120031 57579
rect 77953 57409 77987 57443
rect 79149 57409 79183 57443
rect 81633 57409 81667 57443
rect 64889 57341 64923 57375
rect 64889 57205 64923 57239
rect 64981 57205 65015 57239
rect 65625 57341 65659 57375
rect 62957 56865 62991 56899
rect 62957 56729 62991 56763
rect 69581 56661 69615 56695
rect 69765 56593 69799 56627
rect 82553 57341 82587 57375
rect 119813 57341 119847 57375
rect 119997 57273 120031 57307
rect 120089 57545 120123 57579
rect 82553 57205 82587 57239
rect 115121 57205 115155 57239
rect 119813 57205 119847 57239
rect 91661 57137 91695 57171
rect 102057 57069 102091 57103
rect 91661 56933 91695 56967
rect 99389 56933 99423 56967
rect 122573 57545 122607 57579
rect 130577 57545 130611 57579
rect 122573 57409 122607 57443
rect 129657 57477 129691 57511
rect 124505 57273 124539 57307
rect 124781 57273 124815 57307
rect 129657 57273 129691 57307
rect 119905 57001 119939 57035
rect 102057 56729 102091 56763
rect 102609 56933 102643 56967
rect 102609 56729 102643 56763
rect 102701 56933 102735 56967
rect 102701 56661 102735 56695
rect 115029 56933 115063 56967
rect 115121 56933 115155 56967
rect 115029 56661 115063 56695
rect 128829 56797 128863 56831
rect 99389 56593 99423 56627
rect 128829 56593 128863 56627
rect 79149 56525 79183 56559
rect 141985 57545 142019 57579
rect 132509 57477 132543 57511
rect 132233 57409 132267 57443
rect 132233 57205 132267 57239
rect 130577 56525 130611 56559
rect 100861 52309 100895 52343
rect 98561 48297 98595 48331
rect 100861 48297 100895 48331
rect 121561 51561 121595 51595
rect 121561 48297 121595 48331
rect 151737 57545 151771 57579
rect 141985 57137 142019 57171
rect 147689 57477 147723 57511
rect 151737 57137 151771 57171
rect 191113 57681 191147 57715
rect 191205 57681 191239 57715
rect 191297 57817 191331 57851
rect 176669 57545 176703 57579
rect 191021 57545 191055 57579
rect 191113 57545 191147 57579
rect 185593 57477 185627 57511
rect 173081 57341 173115 57375
rect 176669 57341 176703 57375
rect 185501 57341 185535 57375
rect 185593 57341 185627 57375
rect 156061 57137 156095 57171
rect 169401 57273 169435 57307
rect 169401 56865 169435 56899
rect 147689 56797 147723 56831
rect 142629 56661 142663 56695
rect 142813 56661 142847 56695
rect 171149 56661 171183 56695
rect 212825 57749 212859 57783
rect 191297 57137 191331 57171
rect 195897 57477 195931 57511
rect 191021 57001 191055 57035
rect 211905 57477 211939 57511
rect 195897 57001 195931 57035
rect 195989 57137 196023 57171
rect 185501 56661 185535 56695
rect 173081 56593 173115 56627
rect 171149 56525 171183 56559
rect 132509 48297 132543 48331
rect 224141 57749 224175 57783
rect 224233 57885 224267 57919
rect 224233 57749 224267 57783
rect 215769 57681 215803 57715
rect 215861 57681 215895 57715
rect 212825 57001 212859 57035
rect 211905 56729 211939 56763
rect 538781 57477 538815 57511
rect 224233 57273 224267 57307
rect 538781 57137 538815 57171
rect 224233 56661 224267 56695
rect 215861 56593 215895 56627
rect 336749 56457 336783 56491
rect 195989 48297 196023 48331
rect 334173 55573 334207 55607
rect 334173 48297 334207 48331
rect 98561 46937 98595 46971
rect 336749 46937 336783 46971
rect 338129 46869 338163 46903
rect 101045 38573 101079 38607
rect 192033 38573 192067 38607
rect 101045 31637 101079 31671
rect 128645 37213 128679 37247
rect 145021 35717 145055 35751
rect 145021 28985 145055 29019
rect 192033 28985 192067 29019
rect 195897 38573 195931 38607
rect 338129 37281 338163 37315
rect 195897 28985 195931 29019
rect 336749 37213 336783 37247
rect 128645 27693 128679 27727
rect 336749 27625 336783 27659
rect 121653 27557 121687 27591
rect 128921 27557 128955 27591
rect 212549 27557 212583 27591
rect 128921 19193 128955 19227
rect 192217 19261 192251 19295
rect 121653 17969 121687 18003
rect 212549 17969 212583 18003
rect 338129 27557 338163 27591
rect 192217 9673 192251 9707
rect 333989 17901 334023 17935
rect 195621 9605 195655 9639
rect 106289 6341 106323 6375
rect 55229 4233 55263 4267
rect 22017 4097 22051 4131
rect 35909 4029 35943 4063
rect 22017 3825 22051 3859
rect 26157 3893 26191 3927
rect 35909 3689 35943 3723
rect 45477 4029 45511 4063
rect 45477 3689 45511 3723
rect 45661 4029 45695 4063
rect 26157 3621 26191 3655
rect 36001 3621 36035 3655
rect 36001 3145 36035 3179
rect 45385 3621 45419 3655
rect 64797 4233 64831 4267
rect 55229 3689 55263 3723
rect 59921 4165 59955 4199
rect 96629 4165 96663 4199
rect 75285 4097 75319 4131
rect 84117 4097 84151 4131
rect 96721 4097 96755 4131
rect 106289 4097 106323 4131
rect 88993 4029 89027 4063
rect 156705 3961 156739 3995
rect 88993 3825 89027 3859
rect 148701 3893 148735 3927
rect 84117 3757 84151 3791
rect 64797 3689 64831 3723
rect 64889 3689 64923 3723
rect 59921 3485 59955 3519
rect 69673 3689 69707 3723
rect 75285 3689 75319 3723
rect 68385 3621 68419 3655
rect 68201 3485 68235 3519
rect 65165 3417 65199 3451
rect 45661 3281 45695 3315
rect 45385 3145 45419 3179
rect 71881 3553 71915 3587
rect 71789 3417 71823 3451
rect 82829 3553 82863 3587
rect 82829 3349 82863 3383
rect 104173 3485 104207 3519
rect 156705 3553 156739 3587
rect 161489 3961 161523 3995
rect 169125 3893 169159 3927
rect 161489 3553 161523 3587
rect 166273 3689 166307 3723
rect 148701 3417 148735 3451
rect 104173 3349 104207 3383
rect 169125 3553 169159 3587
rect 191113 3893 191147 3927
rect 191113 3553 191147 3587
rect 166273 3281 166307 3315
rect 69673 3077 69707 3111
rect 143273 2805 143307 2839
rect 143273 561 143307 595
rect 212457 9605 212491 9639
rect 200773 4029 200807 4063
rect 200773 3893 200807 3927
rect 195621 561 195655 595
rect 336749 17901 336783 17935
rect 338129 9673 338163 9707
rect 336749 9537 336783 9571
rect 333989 8313 334023 8347
rect 456257 4165 456291 4199
rect 431233 4097 431267 4131
rect 456073 3893 456107 3927
rect 431233 3757 431267 3791
rect 433165 3757 433199 3791
rect 453773 3757 453807 3791
rect 446689 3689 446723 3723
rect 212457 561 212491 595
rect 213469 2805 213503 2839
rect 213469 561 213503 595
rect 333621 2805 333655 2839
rect 433165 2805 433199 2839
rect 445493 3553 445527 3587
rect 446689 3145 446723 3179
rect 455981 3553 456015 3587
rect 456073 3485 456107 3519
rect 456165 3825 456199 3859
rect 533445 4029 533479 4063
rect 532893 3961 532927 3995
rect 462145 3825 462179 3859
rect 456257 3689 456291 3723
rect 457361 3689 457395 3723
rect 456165 3485 456199 3519
rect 471805 3757 471839 3791
rect 457361 3349 457395 3383
rect 460857 3349 460891 3383
rect 462145 3349 462179 3383
rect 465917 3485 465951 3519
rect 453773 3077 453807 3111
rect 455889 3281 455923 3315
rect 455981 3281 456015 3315
rect 445493 2805 445527 2839
rect 445585 3009 445619 3043
rect 456165 2873 456199 2907
rect 445585 2805 445619 2839
rect 465733 3145 465767 3179
rect 465825 3417 465859 3451
rect 476129 3757 476163 3791
rect 532985 3961 533019 3995
rect 532985 3825 533019 3859
rect 533353 3825 533387 3859
rect 533353 3689 533387 3723
rect 533445 3689 533479 3723
rect 532893 3553 532927 3587
rect 476129 3417 476163 3451
rect 465825 3145 465859 3179
rect 469321 3213 469355 3247
rect 471805 3213 471839 3247
rect 549821 3349 549855 3383
rect 469321 2941 469355 2975
rect 510905 3009 510939 3043
rect 549821 3009 549855 3043
rect 552673 3145 552707 3179
rect 460857 2805 460891 2839
rect 552673 2941 552707 2975
rect 510905 2805 510939 2839
rect 333621 561 333655 595
<< metal1 >>
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 333974 700992 333980 701004
rect 154172 700964 333980 700992
rect 154172 700952 154178 700964
rect 333974 700952 333980 700964
rect 334032 700952 334038 701004
rect 137830 700884 137836 700936
rect 137888 700924 137894 700936
rect 329834 700924 329840 700936
rect 137888 700896 329840 700924
rect 137888 700884 137894 700896
rect 329834 700884 329840 700896
rect 329892 700884 329898 700936
rect 269022 700816 269028 700868
rect 269080 700856 269086 700868
rect 462314 700856 462320 700868
rect 269080 700828 462320 700856
rect 269080 700816 269086 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 273162 700748 273168 700800
rect 273220 700788 273226 700800
rect 478506 700788 478512 700800
rect 273220 700760 478512 700788
rect 273220 700748 273226 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 105446 700680 105452 700732
rect 105504 700720 105510 700732
rect 338114 700720 338120 700732
rect 105504 700692 338120 700720
rect 105504 700680 105510 700692
rect 338114 700680 338120 700692
rect 338172 700680 338178 700732
rect 89162 700612 89168 700664
rect 89220 700652 89226 700664
rect 347866 700652 347872 700664
rect 89220 700624 347872 700652
rect 89220 700612 89226 700624
rect 347866 700612 347872 700624
rect 347924 700612 347930 700664
rect 72970 700544 72976 700596
rect 73028 700584 73034 700596
rect 343634 700584 343640 700596
rect 73028 700556 343640 700584
rect 73028 700544 73034 700556
rect 343634 700544 343640 700556
rect 343692 700544 343698 700596
rect 255222 700476 255228 700528
rect 255280 700516 255286 700528
rect 527174 700516 527180 700528
rect 255280 700488 527180 700516
rect 255280 700476 255286 700488
rect 527174 700476 527180 700488
rect 527232 700476 527238 700528
rect 259362 700408 259368 700460
rect 259420 700448 259426 700460
rect 543458 700448 543464 700460
rect 259420 700420 543464 700448
rect 259420 700408 259426 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 351914 700380 351920 700392
rect 40552 700352 351920 700380
rect 40552 700340 40558 700352
rect 351914 700340 351920 700352
rect 351972 700340 351978 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 360194 700312 360200 700324
rect 24360 700284 360200 700312
rect 24360 700272 24366 700284
rect 360194 700272 360200 700284
rect 360252 700272 360258 700324
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 325694 700244 325700 700256
rect 170364 700216 325700 700244
rect 170364 700204 170370 700216
rect 325694 700204 325700 700216
rect 325752 700204 325758 700256
rect 285582 700136 285588 700188
rect 285640 700176 285646 700188
rect 413646 700176 413652 700188
rect 285640 700148 413652 700176
rect 285640 700136 285646 700148
rect 413646 700136 413652 700148
rect 413704 700136 413710 700188
rect 281442 700068 281448 700120
rect 281500 700108 281506 700120
rect 397454 700108 397460 700120
rect 281500 700080 397460 700108
rect 281500 700068 281506 700080
rect 397454 700068 397460 700080
rect 397512 700068 397518 700120
rect 202782 700000 202788 700052
rect 202840 700040 202846 700052
rect 317414 700040 317420 700052
rect 202840 700012 317420 700040
rect 202840 700000 202846 700012
rect 317414 700000 317420 700012
rect 317472 700000 317478 700052
rect 218974 699932 218980 699984
rect 219032 699972 219038 699984
rect 321554 699972 321560 699984
rect 219032 699944 321560 699972
rect 219032 699932 219038 699944
rect 321554 699932 321560 699944
rect 321612 699932 321618 699984
rect 305089 699907 305147 699913
rect 305089 699873 305101 699907
rect 305135 699904 305147 699907
rect 348786 699904 348792 699916
rect 305135 699876 348792 699904
rect 305135 699873 305147 699876
rect 305089 699867 305147 699873
rect 348786 699864 348792 699876
rect 348844 699864 348850 699916
rect 267642 699796 267648 699848
rect 267700 699836 267706 699848
rect 297913 699839 297971 699845
rect 297913 699836 297925 699839
rect 267700 699808 297925 699836
rect 267700 699796 267706 699808
rect 297913 699805 297925 699808
rect 297959 699805 297971 699839
rect 297913 699799 297971 699805
rect 298002 699796 298008 699848
rect 298060 699836 298066 699848
rect 300029 699839 300087 699845
rect 300029 699836 300041 699839
rect 298060 699808 300041 699836
rect 298060 699796 298066 699808
rect 300029 699805 300041 699808
rect 300075 699805 300087 699839
rect 300029 699799 300087 699805
rect 300118 699796 300124 699848
rect 300176 699836 300182 699848
rect 300762 699836 300768 699848
rect 300176 699808 300768 699836
rect 300176 699796 300182 699808
rect 300762 699796 300768 699808
rect 300820 699796 300826 699848
rect 293862 699728 293868 699780
rect 293920 699768 293926 699780
rect 332502 699768 332508 699780
rect 293920 699740 332508 699768
rect 293920 699728 293926 699740
rect 332502 699728 332508 699740
rect 332560 699728 332566 699780
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 283834 699660 283840 699712
rect 283892 699700 283898 699712
rect 309134 699700 309140 699712
rect 283892 699672 309140 699700
rect 283892 699660 283898 699672
rect 309134 699660 309140 699672
rect 309192 699660 309198 699712
rect 297913 699635 297971 699641
rect 297913 699601 297925 699635
rect 297959 699632 297971 699635
rect 304994 699632 305000 699644
rect 297959 699604 305000 699632
rect 297959 699601 297971 699604
rect 297913 699595 297971 699601
rect 304994 699592 305000 699604
rect 305052 699592 305058 699644
rect 300029 699567 300087 699573
rect 300029 699533 300041 699567
rect 300075 699564 300087 699567
rect 305089 699567 305147 699573
rect 305089 699564 305101 699567
rect 300075 699536 305101 699564
rect 300075 699533 300087 699536
rect 300029 699527 300087 699533
rect 305089 699533 305101 699536
rect 305135 699533 305147 699567
rect 305089 699527 305147 699533
rect 242802 696940 242808 696992
rect 242860 696980 242866 696992
rect 580166 696980 580172 696992
rect 242860 696952 580172 696980
rect 242860 696940 242866 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 364334 692792 364340 692844
rect 364392 692832 364398 692844
rect 365070 692832 365076 692844
rect 364392 692804 365076 692832
rect 364392 692792 364398 692804
rect 365070 692792 365076 692804
rect 365128 692792 365134 692844
rect 246942 685856 246948 685908
rect 247000 685896 247006 685908
rect 580166 685896 580172 685908
rect 247000 685868 580172 685896
rect 247000 685856 247006 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 364334 683068 364340 683120
rect 364392 683108 364398 683120
rect 364610 683108 364616 683120
rect 364392 683080 364616 683108
rect 364392 683068 364398 683080
rect 364610 683068 364616 683080
rect 364668 683068 364674 683120
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 364426 681748 364432 681760
rect 3568 681720 364432 681748
rect 3568 681708 3574 681720
rect 364426 681708 364432 681720
rect 364484 681708 364490 681760
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 364334 673548 364340 673600
rect 364392 673588 364398 673600
rect 364610 673588 364616 673600
rect 364392 673560 364616 673588
rect 364392 673548 364398 673560
rect 364610 673548 364616 673560
rect 364668 673548 364674 673600
rect 238662 673480 238668 673532
rect 238720 673520 238726 673532
rect 580166 673520 580172 673532
rect 238720 673492 580172 673520
rect 238720 673480 238726 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 364334 668584 364340 668636
rect 364392 668624 364398 668636
rect 364518 668624 364524 668636
rect 364392 668596 364524 668624
rect 364392 668584 364398 668596
rect 364518 668584 364524 668596
rect 364576 668584 364582 668636
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 372614 667944 372620 667956
rect 3476 667916 372620 667944
rect 3476 667904 3482 667916
rect 372614 667904 372620 667916
rect 372672 667904 372678 667956
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 288894 663280 288900 663332
rect 288952 663320 288958 663332
rect 364518 663320 364524 663332
rect 288952 663292 364524 663320
rect 288952 663280 288958 663292
rect 364518 663280 364524 663292
rect 364576 663280 364582 663332
rect 235902 663212 235908 663264
rect 235960 663252 235966 663264
rect 314102 663252 314108 663264
rect 235960 663224 314108 663252
rect 235960 663212 235966 663224
rect 314102 663212 314108 663224
rect 314160 663212 314166 663264
rect 276198 663144 276204 663196
rect 276256 663184 276262 663196
rect 429286 663184 429292 663196
rect 276256 663156 429292 663184
rect 276256 663144 276262 663156
rect 429286 663144 429292 663156
rect 429344 663144 429350 663196
rect 263594 663076 263600 663128
rect 263652 663116 263658 663128
rect 494146 663116 494152 663128
rect 263652 663088 494152 663116
rect 263652 663076 263658 663088
rect 494146 663076 494152 663088
rect 494204 663076 494210 663128
rect 250990 663008 250996 663060
rect 251048 663048 251054 663060
rect 559006 663048 559012 663060
rect 251048 663020 559012 663048
rect 251048 663008 251054 663020
rect 559006 663008 559012 663020
rect 559064 663008 559070 663060
rect 300762 662804 300768 662856
rect 300820 662844 300826 662856
rect 301498 662844 301504 662856
rect 300820 662816 301504 662844
rect 300820 662804 300826 662816
rect 301498 662804 301504 662816
rect 301556 662804 301562 662856
rect 204622 662736 204628 662788
rect 204680 662776 204686 662788
rect 539870 662776 539876 662788
rect 204680 662748 539876 662776
rect 204680 662736 204686 662748
rect 539870 662736 539876 662748
rect 539928 662736 539934 662788
rect 192018 662668 192024 662720
rect 192076 662708 192082 662720
rect 539962 662708 539968 662720
rect 192076 662680 539968 662708
rect 192076 662668 192082 662680
rect 539962 662668 539968 662680
rect 540020 662668 540026 662720
rect 8846 662600 8852 662652
rect 8904 662640 8910 662652
rect 394142 662640 394148 662652
rect 8904 662612 394148 662640
rect 8904 662600 8910 662612
rect 394142 662600 394148 662612
rect 394200 662600 394206 662652
rect 9582 662532 9588 662584
rect 9640 662572 9646 662584
rect 406746 662572 406752 662584
rect 9640 662544 406752 662572
rect 9640 662532 9646 662544
rect 406746 662532 406752 662544
rect 406804 662532 406810 662584
rect 175182 662464 175188 662516
rect 175240 662504 175246 662516
rect 577498 662504 577504 662516
rect 175240 662476 577504 662504
rect 175240 662464 175246 662476
rect 577498 662464 577504 662476
rect 577556 662464 577562 662516
rect 9490 662396 9496 662448
rect 9548 662436 9554 662448
rect 432046 662436 432052 662448
rect 9548 662408 432052 662436
rect 9548 662396 9554 662408
rect 432046 662396 432052 662408
rect 432104 662396 432110 662448
rect 95234 662328 95240 662380
rect 95292 662368 95298 662380
rect 232590 662368 232596 662380
rect 95292 662340 232596 662368
rect 95292 662328 95298 662340
rect 232590 662328 232596 662340
rect 232648 662328 232654 662380
rect 233878 662328 233884 662380
rect 233936 662368 233942 662380
rect 398374 662368 398380 662380
rect 233936 662340 398380 662368
rect 233936 662328 233942 662340
rect 398374 662328 398380 662340
rect 398432 662328 398438 662380
rect 208854 662260 208860 662312
rect 208912 662300 208918 662312
rect 381630 662300 381636 662312
rect 208912 662272 381636 662300
rect 208912 662260 208918 662272
rect 381630 662260 381636 662272
rect 381688 662260 381694 662312
rect 230658 662192 230664 662244
rect 230716 662232 230722 662244
rect 419350 662232 419356 662244
rect 230716 662204 419356 662232
rect 230716 662192 230722 662204
rect 419350 662192 419356 662204
rect 419408 662192 419414 662244
rect 213822 662124 213828 662176
rect 213880 662164 213886 662176
rect 448882 662164 448888 662176
rect 213880 662136 448888 662164
rect 213880 662124 213886 662136
rect 448882 662124 448888 662136
rect 448940 662124 448946 662176
rect 112070 662056 112076 662108
rect 112128 662096 112134 662108
rect 369118 662096 369124 662108
rect 112128 662068 369124 662096
rect 112128 662056 112134 662068
rect 369118 662056 369124 662068
rect 369176 662056 369182 662108
rect 196250 661988 196256 662040
rect 196308 662028 196314 662040
rect 540054 662028 540060 662040
rect 196308 662000 540060 662028
rect 196308 661988 196314 662000
rect 540054 661988 540060 662000
rect 540112 661988 540118 662040
rect 107838 661920 107844 661972
rect 107896 661960 107902 661972
rect 169754 661960 169760 661972
rect 107896 661932 169760 661960
rect 107896 661920 107902 661932
rect 169754 661920 169760 661932
rect 169812 661920 169818 661972
rect 183646 661920 183652 661972
rect 183704 661960 183710 661972
rect 541710 661960 541716 661972
rect 183704 661932 541716 661960
rect 183704 661920 183710 661932
rect 541710 661920 541716 661932
rect 541768 661920 541774 661972
rect 91002 661852 91008 661904
rect 91060 661892 91066 661904
rect 165890 661892 165896 661904
rect 91060 661864 165896 661892
rect 91060 661852 91066 661864
rect 165890 661852 165896 661864
rect 165948 661852 165954 661904
rect 170950 661852 170956 661904
rect 171008 661892 171014 661904
rect 541618 661892 541624 661904
rect 171008 661864 541624 661892
rect 171008 661852 171014 661864
rect 541618 661852 541624 661864
rect 541676 661852 541682 661904
rect 166810 661784 166816 661836
rect 166868 661824 166874 661836
rect 540882 661824 540888 661836
rect 166868 661796 540888 661824
rect 166868 661784 166874 661796
rect 540882 661784 540888 661796
rect 540940 661784 540946 661836
rect 120442 661716 120448 661768
rect 120500 661756 120506 661768
rect 158714 661756 158720 661768
rect 120500 661728 158720 661756
rect 120500 661716 120506 661728
rect 158714 661716 158720 661728
rect 158772 661716 158778 661768
rect 162578 661716 162584 661768
rect 162636 661756 162642 661768
rect 538766 661756 538772 661768
rect 162636 661728 538772 661756
rect 162636 661716 162642 661728
rect 538766 661716 538772 661728
rect 538824 661716 538830 661768
rect 154114 661648 154120 661700
rect 154172 661688 154178 661700
rect 540790 661688 540796 661700
rect 154172 661660 540796 661688
rect 154172 661648 154178 661660
rect 540790 661648 540796 661660
rect 540848 661648 540854 661700
rect 82538 661580 82544 661632
rect 82596 661620 82602 661632
rect 155678 661620 155684 661632
rect 82596 661592 155684 661620
rect 82596 661580 82602 661592
rect 155678 661580 155684 661592
rect 155736 661580 155742 661632
rect 158346 661580 158352 661632
rect 158404 661620 158410 661632
rect 548518 661620 548524 661632
rect 158404 661592 548524 661620
rect 158404 661580 158410 661592
rect 548518 661580 548524 661592
rect 548576 661580 548582 661632
rect 53098 661512 53104 661564
rect 53156 661552 53162 661564
rect 444650 661552 444656 661564
rect 53156 661524 444656 661552
rect 53156 661512 53162 661524
rect 444650 661512 444656 661524
rect 444708 661512 444714 661564
rect 145742 661444 145748 661496
rect 145800 661484 145806 661496
rect 540606 661484 540612 661496
rect 145800 661456 540612 661484
rect 145800 661444 145806 661456
rect 540606 661444 540612 661456
rect 540664 661444 540670 661496
rect 141510 661376 141516 661428
rect 141568 661416 141574 661428
rect 540698 661416 540704 661428
rect 141568 661388 540704 661416
rect 141568 661376 141574 661388
rect 540698 661376 540704 661388
rect 540756 661376 540762 661428
rect 54478 661308 54484 661360
rect 54536 661348 54542 661360
rect 457254 661348 457260 661360
rect 54536 661320 457260 661348
rect 54536 661308 54542 661320
rect 457254 661308 457260 661320
rect 457312 661308 457318 661360
rect 457530 661308 457536 661360
rect 457588 661348 457594 661360
rect 495158 661348 495164 661360
rect 457588 661320 495164 661348
rect 457588 661308 457594 661320
rect 495158 661308 495164 661320
rect 495216 661308 495222 661360
rect 4062 661240 4068 661292
rect 4120 661280 4126 661292
rect 436186 661280 436192 661292
rect 4120 661252 436192 661280
rect 4120 661240 4126 661252
rect 436186 661240 436192 661252
rect 436244 661240 436250 661292
rect 448514 661240 448520 661292
rect 448572 661280 448578 661292
rect 528830 661280 528836 661292
rect 448572 661252 528836 661280
rect 448572 661240 448578 661252
rect 528830 661240 528836 661252
rect 528888 661240 528894 661292
rect 103606 661172 103612 661224
rect 103664 661212 103670 661224
rect 540238 661212 540244 661224
rect 103664 661184 540244 661212
rect 103664 661172 103670 661184
rect 540238 661172 540244 661184
rect 540296 661172 540302 661224
rect 9398 661104 9404 661156
rect 9456 661144 9462 661156
rect 461486 661144 461492 661156
rect 9456 661116 461492 661144
rect 9456 661104 9462 661116
rect 461486 661104 461492 661116
rect 461544 661104 461550 661156
rect 9122 661036 9128 661088
rect 9180 661076 9186 661088
rect 486786 661076 486792 661088
rect 9180 661048 486792 661076
rect 9180 661036 9186 661048
rect 486786 661036 486792 661048
rect 486844 661036 486850 661088
rect 3878 660968 3884 661020
rect 3936 661008 3942 661020
rect 213822 661008 213828 661020
rect 3936 660980 213828 661008
rect 3936 660968 3942 660980
rect 213822 660968 213828 660980
rect 213880 660968 213886 661020
rect 225690 660968 225696 661020
rect 225748 661008 225754 661020
rect 538398 661008 538404 661020
rect 225748 660980 538404 661008
rect 225748 660968 225754 660980
rect 538398 660968 538404 660980
rect 538456 660968 538462 661020
rect 213086 660900 213092 660952
rect 213144 660940 213150 660952
rect 538490 660940 538496 660952
rect 213144 660912 538496 660940
rect 213144 660900 213150 660912
rect 538490 660900 538496 660912
rect 538548 660900 538554 660952
rect 200482 660832 200488 660884
rect 200540 660872 200546 660884
rect 538582 660872 538588 660884
rect 200540 660844 538588 660872
rect 200540 660832 200546 660844
rect 538582 660832 538588 660844
rect 538640 660832 538646 660884
rect 187786 660764 187792 660816
rect 187844 660804 187850 660816
rect 538674 660804 538680 660816
rect 187844 660776 538680 660804
rect 187844 660764 187850 660776
rect 538674 660764 538680 660776
rect 538732 660764 538738 660816
rect 8202 660696 8208 660748
rect 8260 660736 8266 660748
rect 377306 660736 377312 660748
rect 8260 660708 377312 660736
rect 8260 660696 8266 660708
rect 377306 660696 377312 660708
rect 377364 660696 377370 660748
rect 8110 660628 8116 660680
rect 8168 660668 8174 660680
rect 389910 660668 389916 660680
rect 8168 660640 389916 660668
rect 8168 660628 8174 660640
rect 389910 660628 389916 660640
rect 389968 660628 389974 660680
rect 149974 660560 149980 660612
rect 150032 660600 150038 660612
rect 539502 660600 539508 660612
rect 150032 660572 539508 660600
rect 150032 660560 150038 660572
rect 539502 660560 539508 660572
rect 539560 660560 539566 660612
rect 8018 660492 8024 660544
rect 8076 660532 8082 660544
rect 402514 660532 402520 660544
rect 8076 660504 402520 660532
rect 8076 660492 8082 660504
rect 402514 660492 402520 660504
rect 402572 660492 402578 660544
rect 7926 660424 7932 660476
rect 7984 660464 7990 660476
rect 415210 660464 415216 660476
rect 7984 660436 415216 660464
rect 7984 660424 7990 660436
rect 415210 660424 415216 660436
rect 415268 660424 415274 660476
rect 169754 660356 169760 660408
rect 169812 660396 169818 660408
rect 580718 660396 580724 660408
rect 169812 660368 580724 660396
rect 169812 660356 169818 660368
rect 580718 660356 580724 660368
rect 580776 660356 580782 660408
rect 158714 660288 158720 660340
rect 158772 660328 158778 660340
rect 580902 660328 580908 660340
rect 158772 660300 580908 660328
rect 158772 660288 158778 660300
rect 580902 660288 580908 660300
rect 580960 660288 580966 660340
rect 133046 660220 133052 660272
rect 133104 660260 133110 660272
rect 540422 660260 540428 660272
rect 133104 660232 540428 660260
rect 133104 660220 133110 660232
rect 540422 660220 540428 660232
rect 540480 660220 540486 660272
rect 58710 660152 58716 660204
rect 58768 660192 58774 660204
rect 474090 660192 474096 660204
rect 58768 660164 474096 660192
rect 58768 660152 58774 660164
rect 474090 660152 474096 660164
rect 474148 660152 474154 660204
rect 7834 660084 7840 660136
rect 7892 660124 7898 660136
rect 427814 660124 427820 660136
rect 7892 660096 427820 660124
rect 7892 660084 7898 660096
rect 427814 660084 427820 660096
rect 427872 660084 427878 660136
rect 7742 660016 7748 660068
rect 7800 660056 7806 660068
rect 440234 660056 440240 660068
rect 7800 660028 440240 660056
rect 7800 660016 7806 660028
rect 440234 660016 440240 660028
rect 440292 660016 440298 660068
rect 99650 659948 99656 660000
rect 99708 659988 99714 660000
rect 539134 659988 539140 660000
rect 99708 659960 539140 659988
rect 99708 659948 99714 659960
rect 539134 659948 539140 659960
rect 539192 659948 539198 660000
rect 7650 659880 7656 659932
rect 7708 659920 7714 659932
rect 452654 659920 452660 659932
rect 7708 659892 452660 659920
rect 7708 659880 7714 659892
rect 452654 659880 452660 659892
rect 452712 659880 452718 659932
rect 7558 659812 7564 659864
rect 7616 659852 7622 659864
rect 465350 659852 465356 659864
rect 7616 659824 465356 659852
rect 7616 659812 7622 659824
rect 465350 659812 465356 659824
rect 465408 659812 465414 659864
rect 9214 659744 9220 659796
rect 9272 659784 9278 659796
rect 478046 659784 478052 659796
rect 9272 659756 478052 659784
rect 9272 659744 9278 659756
rect 478046 659744 478052 659756
rect 478104 659744 478110 659796
rect 6178 659676 6184 659728
rect 6236 659716 6242 659728
rect 490558 659716 490564 659728
rect 6236 659688 490564 659716
rect 6236 659676 6242 659688
rect 490558 659676 490564 659688
rect 490616 659676 490622 659728
rect 3326 659608 3332 659660
rect 3384 659648 3390 659660
rect 230658 659648 230664 659660
rect 3384 659620 230664 659648
rect 3384 659608 3390 659620
rect 230658 659608 230664 659620
rect 230716 659608 230722 659660
rect 368566 659648 368572 659660
rect 368527 659620 368572 659648
rect 368566 659608 368572 659620
rect 368624 659608 368630 659660
rect 369118 659648 369124 659660
rect 369079 659620 369124 659648
rect 369118 659608 369124 659620
rect 369176 659608 369182 659660
rect 381262 659648 381268 659660
rect 381223 659620 381268 659648
rect 381262 659608 381268 659620
rect 381320 659608 381326 659660
rect 381630 659648 381636 659660
rect 381591 659620 381636 659648
rect 381630 659608 381636 659620
rect 381688 659608 381694 659660
rect 385310 659648 385316 659660
rect 385271 659620 385316 659648
rect 385310 659608 385316 659620
rect 385368 659608 385374 659660
rect 410702 659648 410708 659660
rect 410663 659620 410708 659648
rect 410702 659608 410708 659620
rect 410760 659608 410766 659660
rect 423214 659648 423220 659660
rect 423175 659620 423220 659648
rect 423214 659608 423220 659620
rect 423272 659608 423278 659660
rect 469582 659648 469588 659660
rect 469543 659620 469588 659648
rect 469582 659608 469588 659620
rect 469640 659608 469646 659660
rect 3234 659540 3240 659592
rect 3292 659580 3298 659592
rect 233878 659580 233884 659592
rect 3292 659552 233884 659580
rect 3292 659540 3298 659552
rect 233878 659540 233884 659552
rect 233936 659540 233942 659592
rect 234522 659540 234528 659592
rect 234580 659580 234586 659592
rect 541894 659580 541900 659592
rect 234580 659552 541900 659580
rect 234580 659540 234586 659552
rect 541894 659540 541900 659552
rect 541952 659540 541958 659592
rect 230290 659472 230296 659524
rect 230348 659512 230354 659524
rect 539686 659512 539692 659524
rect 230348 659484 539692 659512
rect 230348 659472 230354 659484
rect 539686 659472 539692 659484
rect 539744 659472 539750 659524
rect 221826 659404 221832 659456
rect 221884 659444 221890 659456
rect 541802 659444 541808 659456
rect 221884 659416 541808 659444
rect 221884 659404 221890 659416
rect 541802 659404 541808 659416
rect 541860 659404 541866 659456
rect 179690 659376 179696 659388
rect 179651 659348 179696 659376
rect 179690 659336 179696 659348
rect 179748 659336 179754 659388
rect 217594 659336 217600 659388
rect 217652 659376 217658 659388
rect 539778 659376 539784 659388
rect 217652 659348 539784 659376
rect 217652 659336 217658 659348
rect 539778 659336 539784 659348
rect 539836 659336 539842 659388
rect 116578 659308 116584 659320
rect 116539 659280 116584 659308
rect 116578 659268 116584 659280
rect 116636 659268 116642 659320
rect 125042 659308 125048 659320
rect 125003 659280 125048 659308
rect 125042 659268 125048 659280
rect 125100 659268 125106 659320
rect 129274 659308 129280 659320
rect 129235 659280 129280 659308
rect 129274 659268 129280 659280
rect 129332 659268 129338 659320
rect 137554 659308 137560 659320
rect 137515 659280 137560 659308
rect 137554 659268 137560 659280
rect 137612 659268 137618 659320
rect 165890 659268 165896 659320
rect 165948 659308 165954 659320
rect 580626 659308 580632 659320
rect 165948 659280 580632 659308
rect 165948 659268 165954 659280
rect 580626 659268 580632 659280
rect 580684 659268 580690 659320
rect 179693 659243 179751 659249
rect 179693 659209 179705 659243
rect 179739 659240 179751 659243
rect 540146 659240 540152 659252
rect 179739 659212 540152 659240
rect 179739 659209 179751 659212
rect 179693 659203 179751 659209
rect 540146 659200 540152 659212
rect 540204 659200 540210 659252
rect 8662 659132 8668 659184
rect 8720 659172 8726 659184
rect 368569 659175 368627 659181
rect 368569 659172 368581 659175
rect 8720 659144 368581 659172
rect 8720 659132 8726 659144
rect 368569 659141 368581 659144
rect 368615 659141 368627 659175
rect 368569 659135 368627 659141
rect 369121 659175 369179 659181
rect 369121 659141 369133 659175
rect 369167 659172 369179 659175
rect 580810 659172 580816 659184
rect 369167 659144 580816 659172
rect 369167 659141 369179 659144
rect 369121 659135 369179 659141
rect 580810 659132 580816 659144
rect 580868 659132 580874 659184
rect 8754 659064 8760 659116
rect 8812 659104 8818 659116
rect 381265 659107 381323 659113
rect 381265 659104 381277 659107
rect 8812 659076 381277 659104
rect 8812 659064 8818 659076
rect 381265 659073 381277 659076
rect 381311 659073 381323 659107
rect 381265 659067 381323 659073
rect 381633 659107 381691 659113
rect 381633 659073 381645 659107
rect 381679 659104 381691 659107
rect 580166 659104 580172 659116
rect 381679 659076 580172 659104
rect 381679 659073 381691 659076
rect 381633 659067 381691 659073
rect 580166 659064 580172 659076
rect 580224 659064 580230 659116
rect 5074 658996 5080 659048
rect 5132 659036 5138 659048
rect 385313 659039 385371 659045
rect 385313 659036 385325 659039
rect 5132 659008 385325 659036
rect 5132 658996 5138 659008
rect 385313 659005 385325 659008
rect 385359 659005 385371 659039
rect 385313 658999 385371 659005
rect 137557 658971 137615 658977
rect 137557 658937 137569 658971
rect 137603 658968 137615 658971
rect 539410 658968 539416 658980
rect 137603 658940 539416 658968
rect 137603 658937 137615 658940
rect 137557 658931 137615 658937
rect 539410 658928 539416 658940
rect 539468 658928 539474 658980
rect 4982 658860 4988 658912
rect 5040 658900 5046 658912
rect 410705 658903 410763 658909
rect 410705 658900 410717 658903
rect 5040 658872 410717 658900
rect 5040 658860 5046 658872
rect 410705 658869 410717 658872
rect 410751 658869 410763 658903
rect 410705 658863 410763 658869
rect 129277 658835 129335 658841
rect 129277 658801 129289 658835
rect 129323 658832 129335 658835
rect 540514 658832 540520 658844
rect 129323 658804 540520 658832
rect 129323 658801 129335 658804
rect 129277 658795 129335 658801
rect 540514 658792 540520 658804
rect 540572 658792 540578 658844
rect 125045 658767 125103 658773
rect 125045 658733 125057 658767
rect 125091 658764 125103 658767
rect 539318 658764 539324 658776
rect 125091 658736 539324 658764
rect 125091 658733 125103 658736
rect 125045 658727 125103 658733
rect 539318 658724 539324 658736
rect 539376 658724 539382 658776
rect 4890 658656 4896 658708
rect 4948 658696 4954 658708
rect 423217 658699 423275 658705
rect 423217 658696 423229 658699
rect 4948 658668 423229 658696
rect 4948 658656 4954 658668
rect 423217 658665 423229 658668
rect 423263 658665 423275 658699
rect 423217 658659 423275 658665
rect 116581 658631 116639 658637
rect 116581 658597 116593 658631
rect 116627 658628 116639 658631
rect 540330 658628 540336 658640
rect 116627 658600 540336 658628
rect 116627 658597 116639 658600
rect 116581 658591 116639 658597
rect 540330 658588 540336 658600
rect 540388 658588 540394 658640
rect 9306 658520 9312 658572
rect 9364 658560 9370 658572
rect 469585 658563 469643 658569
rect 469585 658560 469597 658563
rect 9364 658532 469597 658560
rect 9364 658520 9370 658532
rect 469585 658529 469597 658532
rect 469631 658529 469643 658563
rect 469585 658523 469643 658529
rect 3142 653556 3148 653608
rect 3200 653596 3206 653608
rect 8662 653596 8668 653608
rect 3200 653568 8668 653596
rect 3200 653556 3206 653568
rect 8662 653556 8668 653568
rect 8720 653556 8726 653608
rect 539686 651312 539692 651364
rect 539744 651352 539750 651364
rect 580074 651352 580080 651364
rect 539744 651324 580080 651352
rect 539744 651312 539750 651324
rect 580074 651312 580080 651324
rect 580132 651312 580138 651364
rect 541894 640228 541900 640280
rect 541952 640268 541958 640280
rect 580074 640268 580080 640280
rect 541952 640240 580080 640268
rect 541952 640228 541958 640240
rect 580074 640228 580080 640240
rect 580132 640228 580138 640280
rect 539594 627852 539600 627904
rect 539652 627892 539658 627904
rect 580074 627892 580080 627904
rect 539652 627864 580080 627892
rect 539652 627852 539658 627864
rect 580074 627852 580080 627864
rect 580132 627852 580138 627904
rect 3142 624860 3148 624912
rect 3200 624900 3206 624912
rect 8202 624900 8208 624912
rect 3200 624872 8208 624900
rect 3200 624860 3206 624872
rect 8202 624860 8208 624872
rect 8260 624860 8266 624912
rect 2774 610444 2780 610496
rect 2832 610484 2838 610496
rect 5074 610484 5080 610496
rect 2832 610456 5080 610484
rect 2832 610444 2838 610456
rect 5074 610444 5080 610456
rect 5132 610444 5138 610496
rect 539778 604392 539784 604444
rect 539836 604432 539842 604444
rect 580074 604432 580080 604444
rect 539836 604404 580080 604432
rect 539836 604392 539842 604404
rect 580074 604392 580080 604404
rect 580132 604392 580138 604444
rect 3142 596028 3148 596080
rect 3200 596068 3206 596080
rect 8754 596068 8760 596080
rect 3200 596040 8760 596068
rect 3200 596028 3206 596040
rect 8754 596028 8760 596040
rect 8812 596028 8818 596080
rect 541802 593308 541808 593360
rect 541860 593348 541866 593360
rect 580074 593348 580080 593360
rect 541860 593320 580080 593348
rect 541860 593308 541866 593320
rect 580074 593308 580080 593320
rect 580132 593308 580138 593360
rect 538490 580932 538496 580984
rect 538548 580972 538554 580984
rect 580074 580972 580080 580984
rect 538548 580944 580080 580972
rect 538548 580932 538554 580944
rect 580074 580932 580080 580944
rect 580132 580932 580138 580984
rect 3142 567536 3148 567588
rect 3200 567576 3206 567588
rect 8110 567576 8116 567588
rect 3200 567548 8116 567576
rect 3200 567536 3206 567548
rect 8110 567536 8116 567548
rect 8168 567536 8174 567588
rect 539870 557472 539876 557524
rect 539928 557512 539934 557524
rect 580074 557512 580080 557524
rect 539928 557484 580080 557512
rect 539928 557472 539934 557484
rect 580074 557472 580080 557484
rect 580132 557472 580138 557524
rect 3234 538772 3240 538824
rect 3292 538812 3298 538824
rect 8846 538812 8852 538824
rect 3292 538784 8852 538812
rect 3292 538772 3298 538784
rect 8846 538772 8852 538784
rect 8904 538772 8910 538824
rect 538582 534012 538588 534064
rect 538640 534052 538646 534064
rect 580166 534052 580172 534064
rect 538640 534024 580172 534052
rect 538640 534012 538646 534024
rect 580166 534012 580172 534024
rect 580224 534012 580230 534064
rect 539962 510552 539968 510604
rect 540020 510592 540026 510604
rect 579798 510592 579804 510604
rect 540020 510564 579804 510592
rect 540020 510552 540026 510564
rect 579798 510552 579804 510564
rect 579856 510552 579862 510604
rect 3234 510008 3240 510060
rect 3292 510048 3298 510060
rect 8018 510048 8024 510060
rect 3292 510020 8024 510048
rect 3292 510008 3298 510020
rect 8018 510008 8024 510020
rect 8076 510008 8082 510060
rect 540054 499468 540060 499520
rect 540112 499508 540118 499520
rect 579982 499508 579988 499520
rect 540112 499480 579988 499508
rect 540112 499468 540118 499480
rect 579982 499468 579988 499480
rect 580040 499468 580046 499520
rect 2774 496680 2780 496732
rect 2832 496720 2838 496732
rect 4982 496720 4988 496732
rect 2832 496692 4988 496720
rect 2832 496680 2838 496692
rect 4982 496680 4988 496692
rect 5040 496680 5046 496732
rect 538674 487092 538680 487144
rect 538732 487132 538738 487144
rect 580166 487132 580172 487144
rect 538732 487104 580172 487132
rect 538732 487092 538738 487104
rect 580166 487092 580172 487104
rect 580224 487092 580230 487144
rect 3234 481176 3240 481228
rect 3292 481216 3298 481228
rect 9582 481216 9588 481228
rect 3292 481188 9588 481216
rect 3292 481176 3298 481188
rect 9582 481176 9588 481188
rect 9640 481176 9646 481228
rect 540146 463632 540152 463684
rect 540204 463672 540210 463684
rect 579798 463672 579804 463684
rect 540204 463644 579804 463672
rect 540204 463632 540210 463644
rect 579798 463632 579804 463644
rect 579856 463632 579862 463684
rect 541710 452548 541716 452600
rect 541768 452588 541774 452600
rect 579982 452588 579988 452600
rect 541768 452560 579988 452588
rect 541768 452548 541774 452560
rect 579982 452548 579988 452560
rect 580040 452548 580046 452600
rect 3234 452412 3240 452464
rect 3292 452452 3298 452464
rect 7926 452452 7932 452464
rect 3292 452424 7932 452452
rect 3292 452412 3298 452424
rect 7926 452412 7932 452424
rect 7984 452412 7990 452464
rect 577498 440172 577504 440224
rect 577556 440212 577562 440224
rect 579706 440212 579712 440224
rect 577556 440184 579712 440212
rect 577556 440172 577562 440184
rect 579706 440172 579712 440184
rect 579764 440172 579770 440224
rect 2774 438744 2780 438796
rect 2832 438784 2838 438796
rect 4890 438784 4896 438796
rect 2832 438756 4896 438784
rect 2832 438744 2838 438756
rect 4890 438744 4896 438756
rect 4948 438744 4954 438796
rect 540882 416712 540888 416764
rect 540940 416752 540946 416764
rect 579798 416752 579804 416764
rect 540940 416724 579804 416752
rect 540940 416712 540946 416724
rect 579798 416712 579804 416724
rect 579856 416712 579862 416764
rect 541618 405628 541624 405680
rect 541676 405668 541682 405680
rect 579982 405668 579988 405680
rect 541676 405640 579988 405668
rect 541676 405628 541682 405640
rect 579982 405628 579988 405640
rect 580040 405628 580046 405680
rect 3326 395224 3332 395276
rect 3384 395264 3390 395276
rect 7834 395264 7840 395276
rect 3384 395236 7840 395264
rect 3384 395224 3390 395236
rect 7834 395224 7840 395236
rect 7892 395224 7898 395276
rect 538766 393252 538772 393304
rect 538824 393292 538830 393304
rect 580166 393292 580172 393304
rect 538824 393264 580172 393292
rect 538824 393252 538830 393264
rect 580166 393252 580172 393264
rect 580224 393252 580230 393304
rect 540790 369792 540796 369844
rect 540848 369832 540854 369844
rect 579798 369832 579804 369844
rect 540848 369804 579804 369832
rect 540848 369792 540854 369804
rect 579798 369792 579804 369804
rect 579856 369792 579862 369844
rect 3142 366664 3148 366716
rect 3200 366704 3206 366716
rect 9490 366704 9496 366716
rect 3200 366676 9496 366704
rect 3200 366664 3206 366676
rect 9490 366664 9496 366676
rect 9548 366664 9554 366716
rect 548518 358708 548524 358760
rect 548576 358748 548582 358760
rect 579982 358748 579988 358760
rect 548576 358720 579988 358748
rect 548576 358708 548582 358720
rect 579982 358708 579988 358720
rect 580040 358708 580046 358760
rect 539502 346332 539508 346384
rect 539560 346372 539566 346384
rect 580166 346372 580172 346384
rect 539560 346344 580172 346372
rect 539560 346332 539566 346344
rect 580166 346332 580172 346344
rect 580224 346332 580230 346384
rect 3326 337492 3332 337544
rect 3384 337532 3390 337544
rect 7742 337532 7748 337544
rect 3384 337504 7748 337532
rect 3384 337492 3390 337504
rect 7742 337492 7748 337504
rect 7800 337492 7806 337544
rect 540698 322872 540704 322924
rect 540756 322912 540762 322924
rect 579798 322912 579804 322924
rect 540756 322884 579804 322912
rect 540756 322872 540762 322884
rect 579798 322872 579804 322884
rect 579856 322872 579862 322924
rect 540606 311788 540612 311840
rect 540664 311828 540670 311840
rect 579982 311828 579988 311840
rect 540664 311800 579988 311828
rect 540664 311788 540670 311800
rect 579982 311788 579988 311800
rect 580040 311788 580046 311840
rect 3050 309068 3056 309120
rect 3108 309108 3114 309120
rect 53098 309108 53104 309120
rect 3108 309080 53104 309108
rect 3108 309068 3114 309080
rect 53098 309068 53104 309080
rect 53156 309068 53162 309120
rect 539410 299412 539416 299464
rect 539468 299452 539474 299464
rect 580166 299452 580172 299464
rect 539468 299424 580172 299452
rect 539468 299412 539474 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 3142 294788 3148 294840
rect 3200 294828 3206 294840
rect 7650 294828 7656 294840
rect 3200 294800 7656 294828
rect 3200 294788 3206 294800
rect 7650 294788 7656 294800
rect 7708 294788 7714 294840
rect 3326 280100 3332 280152
rect 3384 280140 3390 280152
rect 9398 280140 9404 280152
rect 3384 280112 9404 280140
rect 3384 280100 3390 280112
rect 9398 280100 9404 280112
rect 9456 280100 9462 280152
rect 540514 275952 540520 276004
rect 540572 275992 540578 276004
rect 579798 275992 579804 276004
rect 540572 275964 579804 275992
rect 540572 275952 540578 275964
rect 579798 275952 579804 275964
rect 579856 275952 579862 276004
rect 3326 266296 3332 266348
rect 3384 266336 3390 266348
rect 54478 266336 54484 266348
rect 3384 266308 54484 266336
rect 3384 266296 3390 266308
rect 54478 266296 54484 266308
rect 54536 266296 54542 266348
rect 540422 264868 540428 264920
rect 540480 264908 540486 264920
rect 579982 264908 579988 264920
rect 540480 264880 579988 264908
rect 540480 264868 540486 264880
rect 579982 264868 579988 264880
rect 580040 264868 580046 264920
rect 539318 252492 539324 252544
rect 539376 252532 539382 252544
rect 580166 252532 580172 252544
rect 539376 252504 580172 252532
rect 539376 252492 539382 252504
rect 580166 252492 580172 252504
rect 580224 252492 580230 252544
rect 3326 252220 3332 252272
rect 3384 252260 3390 252272
rect 7558 252260 7564 252272
rect 3384 252232 7564 252260
rect 3384 252220 3390 252232
rect 7558 252220 7564 252232
rect 7616 252220 7622 252272
rect 3326 237328 3332 237380
rect 3384 237368 3390 237380
rect 58710 237368 58716 237380
rect 3384 237340 58716 237368
rect 3384 237328 3390 237340
rect 58710 237328 58716 237340
rect 58768 237328 58774 237380
rect 540330 229032 540336 229084
rect 540388 229072 540394 229084
rect 579798 229072 579804 229084
rect 540388 229044 579804 229072
rect 540388 229032 540394 229044
rect 579798 229032 579804 229044
rect 579856 229032 579862 229084
rect 3326 223048 3332 223100
rect 3384 223088 3390 223100
rect 9306 223088 9312 223100
rect 3384 223060 9312 223088
rect 3384 223048 3390 223060
rect 9306 223048 9312 223060
rect 9364 223048 9370 223100
rect 3326 208156 3332 208208
rect 3384 208196 3390 208208
rect 9214 208196 9220 208208
rect 3384 208168 9220 208196
rect 3384 208156 3390 208168
rect 9214 208156 9220 208168
rect 9272 208156 9278 208208
rect 3326 194488 3332 194540
rect 3384 194528 3390 194540
rect 9122 194528 9128 194540
rect 3384 194500 9128 194528
rect 3384 194488 3390 194500
rect 9122 194488 9128 194500
rect 9180 194488 9186 194540
rect 540238 182112 540244 182164
rect 540296 182152 540302 182164
rect 580166 182152 580172 182164
rect 540296 182124 580172 182152
rect 540296 182112 540302 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 3326 179596 3332 179648
rect 3384 179636 3390 179648
rect 9030 179636 9036 179648
rect 3384 179608 9036 179636
rect 3384 179596 3390 179608
rect 9030 179596 9036 179608
rect 9088 179596 9094 179648
rect 3050 165452 3056 165504
rect 3108 165492 3114 165504
rect 6178 165492 6184 165504
rect 3108 165464 6184 165492
rect 3108 165452 3114 165464
rect 6178 165452 6184 165464
rect 6236 165452 6242 165504
rect 539134 158652 539140 158704
rect 539192 158692 539198 158704
rect 580166 158692 580172 158704
rect 539192 158664 580172 158692
rect 539192 158652 539198 158664
rect 580166 158652 580172 158664
rect 580224 158652 580230 158704
rect 3326 122748 3332 122800
rect 3384 122788 3390 122800
rect 25498 122788 25504 122800
rect 3384 122760 25504 122788
rect 3384 122748 3390 122760
rect 25498 122748 25504 122760
rect 25556 122748 25562 122800
rect 539226 111732 539232 111784
rect 539284 111772 539290 111784
rect 580166 111772 580172 111784
rect 539284 111744 580172 111772
rect 539284 111732 539290 111744
rect 580166 111732 580172 111744
rect 580224 111732 580230 111784
rect 3326 93780 3332 93832
rect 3384 93820 3390 93832
rect 58618 93820 58624 93832
rect 3384 93792 58624 93820
rect 3384 93780 3390 93792
rect 58618 93780 58624 93792
rect 58676 93780 58682 93832
rect 538950 88272 538956 88324
rect 539008 88312 539014 88324
rect 580166 88312 580172 88324
rect 539008 88284 580172 88312
rect 539008 88272 539014 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 3142 79092 3148 79144
rect 3200 79132 3206 79144
rect 8938 79132 8944 79144
rect 3200 79104 8944 79132
rect 3200 79092 3206 79104
rect 8938 79092 8944 79104
rect 8996 79092 9002 79144
rect 539042 64812 539048 64864
rect 539100 64852 539106 64864
rect 579614 64852 579620 64864
rect 539100 64824 579620 64852
rect 539100 64812 539106 64824
rect 579614 64812 579620 64824
rect 579672 64812 579678 64864
rect 2774 64540 2780 64592
rect 2832 64580 2838 64592
rect 4798 64580 4804 64592
rect 2832 64552 4804 64580
rect 2832 64540 2838 64552
rect 4798 64540 4804 64552
rect 4856 64540 4862 64592
rect 60734 57944 60740 57996
rect 60792 57984 60798 57996
rect 61654 57984 61660 57996
rect 60792 57956 61660 57984
rect 60792 57944 60798 57956
rect 61654 57944 61660 57956
rect 61712 57944 61718 57996
rect 224129 57987 224187 57993
rect 224129 57953 224141 57987
rect 224175 57984 224187 57987
rect 224175 57956 224356 57984
rect 224175 57953 224187 57956
rect 224129 57947 224187 57953
rect 44082 57876 44088 57928
rect 44140 57916 44146 57928
rect 95234 57916 95240 57928
rect 44140 57888 95240 57916
rect 44140 57876 44146 57888
rect 95234 57876 95240 57888
rect 95292 57876 95298 57928
rect 108942 57876 108948 57928
rect 109000 57916 109006 57928
rect 109000 57888 112024 57916
rect 109000 57876 109006 57888
rect 41322 57808 41328 57860
rect 41380 57848 41386 57860
rect 93210 57848 93216 57860
rect 41380 57820 93216 57848
rect 41380 57808 41386 57820
rect 93210 57808 93216 57820
rect 93268 57808 93274 57860
rect 100662 57808 100668 57860
rect 100720 57848 100726 57860
rect 100720 57820 103192 57848
rect 100720 57808 100726 57820
rect 38470 57740 38476 57792
rect 38528 57780 38534 57792
rect 90358 57780 90364 57792
rect 38528 57752 90364 57780
rect 38528 57740 38534 57752
rect 90358 57740 90364 57752
rect 90416 57740 90422 57792
rect 96522 57740 96528 57792
rect 96580 57780 96586 57792
rect 103164 57780 103192 57820
rect 104158 57808 104164 57860
rect 104216 57848 104222 57860
rect 111886 57848 111892 57860
rect 104216 57820 111892 57848
rect 104216 57808 104222 57820
rect 111886 57808 111892 57820
rect 111944 57808 111950 57860
rect 111996 57848 112024 57888
rect 113082 57876 113088 57928
rect 113140 57916 113146 57928
rect 151998 57916 152004 57928
rect 113140 57888 152004 57916
rect 113140 57876 113146 57888
rect 151998 57876 152004 57888
rect 152056 57876 152062 57928
rect 152458 57876 152464 57928
rect 152516 57916 152522 57928
rect 156966 57916 156972 57928
rect 152516 57888 156972 57916
rect 152516 57876 152522 57888
rect 156966 57876 156972 57888
rect 157024 57876 157030 57928
rect 158622 57876 158628 57928
rect 158680 57916 158686 57928
rect 189258 57916 189264 57928
rect 158680 57888 189264 57916
rect 158680 57876 158686 57888
rect 189258 57876 189264 57888
rect 189316 57876 189322 57928
rect 190362 57876 190368 57928
rect 190420 57916 190426 57928
rect 215662 57916 215668 57928
rect 190420 57888 215668 57916
rect 190420 57876 190426 57888
rect 215662 57876 215668 57888
rect 215720 57876 215726 57928
rect 215757 57919 215815 57925
rect 215757 57885 215769 57919
rect 215803 57916 215815 57919
rect 224221 57919 224279 57925
rect 224221 57916 224233 57919
rect 215803 57888 224233 57916
rect 215803 57885 215815 57888
rect 215757 57879 215815 57885
rect 224221 57885 224233 57888
rect 224267 57885 224279 57919
rect 224328 57916 224356 57956
rect 242158 57916 242164 57928
rect 224328 57888 242164 57916
rect 224221 57879 224279 57885
rect 242158 57876 242164 57888
rect 242216 57876 242222 57928
rect 245562 57876 245568 57928
rect 245620 57916 245626 57928
rect 261754 57916 261760 57928
rect 245620 57888 261760 57916
rect 245620 57876 245626 57888
rect 261754 57876 261760 57888
rect 261812 57876 261818 57928
rect 263502 57876 263508 57928
rect 263560 57916 263566 57928
rect 275462 57916 275468 57928
rect 263560 57888 275468 57916
rect 263560 57876 263566 57888
rect 275462 57876 275468 57888
rect 275520 57876 275526 57928
rect 280062 57876 280068 57928
rect 280120 57916 280126 57928
rect 289170 57916 289176 57928
rect 280120 57888 289176 57916
rect 280120 57876 280126 57888
rect 289170 57876 289176 57888
rect 289228 57876 289234 57928
rect 460566 57876 460572 57928
rect 460624 57916 460630 57928
rect 485958 57916 485964 57928
rect 460624 57888 485964 57916
rect 460624 57876 460630 57888
rect 485958 57876 485964 57888
rect 486016 57876 486022 57928
rect 497826 57876 497832 57928
rect 497884 57916 497890 57928
rect 529198 57916 529204 57928
rect 497884 57888 529204 57916
rect 497884 57876 497890 57888
rect 529198 57876 529204 57888
rect 529256 57876 529262 57928
rect 149054 57848 149060 57860
rect 111996 57820 149060 57848
rect 149054 57808 149060 57820
rect 149112 57808 149118 57860
rect 150342 57808 150348 57860
rect 150400 57848 150406 57860
rect 182358 57848 182364 57860
rect 150400 57820 182364 57848
rect 150400 57808 150406 57820
rect 182358 57808 182364 57820
rect 182416 57808 182422 57860
rect 183462 57808 183468 57860
rect 183520 57848 183526 57860
rect 191193 57851 191251 57857
rect 191193 57848 191205 57851
rect 183520 57820 191205 57848
rect 183520 57808 183526 57820
rect 191193 57817 191205 57820
rect 191239 57817 191251 57851
rect 191193 57811 191251 57817
rect 191285 57851 191343 57857
rect 191285 57817 191297 57851
rect 191331 57848 191343 57851
rect 214742 57848 214748 57860
rect 191331 57820 214748 57848
rect 191331 57817 191343 57820
rect 191285 57811 191343 57817
rect 214742 57808 214748 57820
rect 214800 57808 214806 57860
rect 215202 57808 215208 57860
rect 215260 57848 215266 57860
rect 236270 57848 236276 57860
rect 215260 57820 236276 57848
rect 215260 57808 215266 57820
rect 236270 57808 236276 57820
rect 236328 57808 236334 57860
rect 240042 57808 240048 57860
rect 240100 57848 240106 57860
rect 256878 57848 256884 57860
rect 240100 57820 256884 57848
rect 240100 57808 240106 57820
rect 256878 57808 256884 57820
rect 256936 57808 256942 57860
rect 259362 57808 259368 57860
rect 259420 57848 259426 57860
rect 272518 57848 272524 57860
rect 259420 57820 272524 57848
rect 259420 57808 259426 57820
rect 272518 57808 272524 57820
rect 272576 57808 272582 57860
rect 274542 57808 274548 57860
rect 274600 57848 274606 57860
rect 285214 57848 285220 57860
rect 274600 57820 285220 57848
rect 274600 57808 274606 57820
rect 285214 57808 285220 57820
rect 285272 57808 285278 57860
rect 319438 57808 319444 57860
rect 319496 57848 319502 57860
rect 321462 57848 321468 57860
rect 319496 57820 321468 57848
rect 319496 57808 319502 57820
rect 321462 57808 321468 57820
rect 321520 57808 321526 57860
rect 480162 57808 480168 57860
rect 480220 57848 480226 57860
rect 489178 57848 489184 57860
rect 480220 57820 489184 57848
rect 480220 57808 480226 57820
rect 489178 57808 489184 57820
rect 489236 57808 489242 57860
rect 519354 57808 519360 57860
rect 519412 57848 519418 57860
rect 520182 57848 520188 57860
rect 519412 57820 520188 57848
rect 519412 57808 519418 57820
rect 520182 57808 520188 57820
rect 520240 57808 520246 57860
rect 520366 57808 520372 57860
rect 520424 57848 520430 57860
rect 521562 57848 521568 57860
rect 520424 57820 521568 57848
rect 520424 57808 520430 57820
rect 521562 57808 521568 57820
rect 521620 57808 521626 57860
rect 527174 57808 527180 57860
rect 527232 57848 527238 57860
rect 528462 57848 528468 57860
rect 527232 57820 528468 57848
rect 527232 57808 527238 57820
rect 528462 57808 528468 57820
rect 528520 57808 528526 57860
rect 532694 57848 532700 57860
rect 530044 57820 532700 57848
rect 142246 57780 142252 57792
rect 96580 57752 103100 57780
rect 103164 57752 142252 57780
rect 96580 57740 96586 57752
rect 38562 57672 38568 57724
rect 38620 57712 38626 57724
rect 91278 57712 91284 57724
rect 38620 57684 91284 57712
rect 38620 57672 38626 57684
rect 91278 57672 91284 57684
rect 91336 57672 91342 57724
rect 93762 57672 93768 57724
rect 93820 57712 93826 57724
rect 103072 57712 103100 57752
rect 142246 57740 142252 57752
rect 142304 57740 142310 57792
rect 142798 57740 142804 57792
rect 142856 57780 142862 57792
rect 151078 57780 151084 57792
rect 142856 57752 151084 57780
rect 142856 57740 142862 57752
rect 151078 57740 151084 57752
rect 151136 57740 151142 57792
rect 153838 57740 153844 57792
rect 153896 57780 153902 57792
rect 155954 57780 155960 57792
rect 153896 57752 155960 57780
rect 153896 57740 153902 57752
rect 155954 57740 155960 57752
rect 156012 57740 156018 57792
rect 156049 57783 156107 57789
rect 156049 57749 156061 57783
rect 156095 57780 156107 57783
rect 185302 57780 185308 57792
rect 156095 57752 185308 57780
rect 156095 57749 156107 57752
rect 156049 57743 156107 57749
rect 185302 57740 185308 57752
rect 185360 57740 185366 57792
rect 186222 57740 186228 57792
rect 186280 57780 186286 57792
rect 212718 57780 212724 57792
rect 186280 57752 212724 57780
rect 186280 57740 186286 57752
rect 212718 57740 212724 57752
rect 212776 57740 212782 57792
rect 212813 57783 212871 57789
rect 212813 57749 212825 57783
rect 212859 57780 212871 57783
rect 221550 57780 221556 57792
rect 212859 57752 221556 57780
rect 212859 57749 212871 57752
rect 212813 57743 212871 57749
rect 221550 57740 221556 57752
rect 221608 57740 221614 57792
rect 222102 57740 222108 57792
rect 222160 57780 222166 57792
rect 224129 57783 224187 57789
rect 224129 57780 224141 57783
rect 222160 57752 224141 57780
rect 222160 57740 222166 57752
rect 224129 57749 224141 57752
rect 224175 57749 224187 57783
rect 224129 57743 224187 57749
rect 224221 57783 224279 57789
rect 224221 57749 224233 57783
rect 224267 57780 224279 57783
rect 235258 57780 235264 57792
rect 224267 57752 235264 57780
rect 224267 57749 224279 57752
rect 224221 57743 224279 57749
rect 235258 57740 235264 57752
rect 235316 57740 235322 57792
rect 237282 57740 237288 57792
rect 237340 57780 237346 57792
rect 253934 57780 253940 57792
rect 237340 57752 253940 57780
rect 237340 57740 237346 57752
rect 253934 57740 253940 57752
rect 253992 57740 253998 57792
rect 257982 57740 257988 57792
rect 258040 57780 258046 57792
rect 271506 57780 271512 57792
rect 258040 57752 271512 57780
rect 258040 57740 258046 57752
rect 271506 57740 271512 57752
rect 271564 57740 271570 57792
rect 275922 57740 275928 57792
rect 275980 57780 275986 57792
rect 286226 57780 286232 57792
rect 275980 57752 286232 57780
rect 275980 57740 275986 57752
rect 286226 57740 286232 57752
rect 286284 57740 286290 57792
rect 326982 57740 326988 57792
rect 327040 57780 327046 57792
rect 328362 57780 328368 57792
rect 327040 57752 328368 57780
rect 327040 57740 327046 57752
rect 328362 57740 328368 57752
rect 328420 57740 328426 57792
rect 347958 57740 347964 57792
rect 348016 57780 348022 57792
rect 349062 57780 349068 57792
rect 348016 57752 349068 57780
rect 348016 57740 348022 57752
rect 349062 57740 349068 57752
rect 349120 57740 349126 57792
rect 371418 57740 371424 57792
rect 371476 57780 371482 57792
rect 374638 57780 374644 57792
rect 371476 57752 374644 57780
rect 371476 57740 371482 57752
rect 374638 57740 374644 57752
rect 374696 57740 374702 57792
rect 482094 57740 482100 57792
rect 482152 57780 482158 57792
rect 482922 57780 482928 57792
rect 482152 57752 482928 57780
rect 482152 57740 482158 57752
rect 482922 57740 482928 57752
rect 482980 57740 482986 57792
rect 483106 57740 483112 57792
rect 483164 57780 483170 57792
rect 484302 57780 484308 57792
rect 483164 57752 484308 57780
rect 483164 57740 483170 57752
rect 484302 57740 484308 57752
rect 484360 57740 484366 57792
rect 488994 57740 489000 57792
rect 489052 57780 489058 57792
rect 489822 57780 489828 57792
rect 489052 57752 489828 57780
rect 489052 57740 489058 57752
rect 489822 57740 489828 57752
rect 489880 57740 489886 57792
rect 498746 57740 498752 57792
rect 498804 57780 498810 57792
rect 530044 57780 530072 57820
rect 532694 57808 532700 57820
rect 532752 57808 532758 57860
rect 533062 57808 533068 57860
rect 533120 57848 533126 57860
rect 533120 57820 535684 57848
rect 533120 57808 533126 57820
rect 498804 57752 530072 57780
rect 498804 57740 498810 57752
rect 530118 57740 530124 57792
rect 530176 57780 530182 57792
rect 531222 57780 531228 57792
rect 530176 57752 531228 57780
rect 530176 57740 530182 57752
rect 531222 57740 531228 57752
rect 531280 57740 531286 57792
rect 534074 57740 534080 57792
rect 534132 57780 534138 57792
rect 535362 57780 535368 57792
rect 534132 57752 535368 57780
rect 534132 57740 534138 57752
rect 535362 57740 535368 57752
rect 535420 57740 535426 57792
rect 535656 57780 535684 57820
rect 537018 57808 537024 57860
rect 537076 57848 537082 57860
rect 538122 57848 538128 57860
rect 537076 57820 538128 57848
rect 537076 57808 537082 57820
rect 538122 57808 538128 57820
rect 538180 57808 538186 57860
rect 541618 57780 541624 57792
rect 535656 57752 541624 57780
rect 541618 57740 541624 57752
rect 541676 57740 541682 57792
rect 138290 57712 138296 57724
rect 93820 57684 96108 57712
rect 103072 57684 138296 57712
rect 93820 57672 93826 57684
rect 30190 57604 30196 57656
rect 30248 57644 30254 57656
rect 77941 57647 77999 57653
rect 77941 57644 77953 57647
rect 30248 57616 77953 57644
rect 30248 57604 30254 57616
rect 77941 57613 77953 57616
rect 77987 57613 77999 57647
rect 77941 57607 77999 57613
rect 78030 57604 78036 57656
rect 78088 57644 78094 57656
rect 81526 57644 81532 57656
rect 78088 57616 81532 57644
rect 78088 57604 78094 57616
rect 81526 57604 81532 57616
rect 81584 57604 81590 57656
rect 81621 57647 81679 57653
rect 81621 57613 81633 57647
rect 81667 57644 81679 57647
rect 83553 57647 83611 57653
rect 83553 57644 83565 57647
rect 81667 57616 83565 57644
rect 81667 57613 81679 57616
rect 81621 57607 81679 57613
rect 83553 57613 83565 57616
rect 83599 57613 83611 57647
rect 83553 57607 83611 57613
rect 85482 57604 85488 57656
rect 85540 57644 85546 57656
rect 94593 57647 94651 57653
rect 94593 57644 94605 57647
rect 85540 57616 94605 57644
rect 85540 57604 85546 57616
rect 94593 57613 94605 57616
rect 94639 57613 94651 57647
rect 96080 57644 96108 57684
rect 138290 57672 138296 57684
rect 138348 57672 138354 57724
rect 139118 57672 139124 57724
rect 139176 57712 139182 57724
rect 139176 57684 147352 57712
rect 139176 57672 139182 57684
rect 136358 57644 136364 57656
rect 96080 57616 136364 57644
rect 94593 57607 94651 57613
rect 136358 57604 136364 57616
rect 136416 57604 136422 57656
rect 140682 57604 140688 57656
rect 140740 57644 140746 57656
rect 147324 57644 147352 57684
rect 147582 57672 147588 57724
rect 147640 57712 147646 57724
rect 180426 57712 180432 57724
rect 147640 57684 180432 57712
rect 147640 57672 147646 57684
rect 180426 57672 180432 57684
rect 180484 57672 180490 57724
rect 182082 57672 182088 57724
rect 182140 57712 182146 57724
rect 191101 57715 191159 57721
rect 191101 57712 191113 57715
rect 182140 57684 191113 57712
rect 182140 57672 182146 57684
rect 191101 57681 191113 57684
rect 191147 57681 191159 57715
rect 191101 57675 191159 57681
rect 191193 57715 191251 57721
rect 191193 57681 191205 57715
rect 191239 57712 191251 57715
rect 209774 57712 209780 57724
rect 191239 57684 209780 57712
rect 191239 57681 191251 57684
rect 191193 57675 191251 57681
rect 209774 57672 209780 57684
rect 209832 57672 209838 57724
rect 213822 57672 213828 57724
rect 213880 57712 213886 57724
rect 215757 57715 215815 57721
rect 215757 57712 215769 57715
rect 213880 57684 215769 57712
rect 213880 57672 213886 57684
rect 215757 57681 215769 57684
rect 215803 57681 215815 57715
rect 215757 57675 215815 57681
rect 215849 57715 215907 57721
rect 215849 57681 215861 57715
rect 215895 57712 215907 57715
rect 232314 57712 232320 57724
rect 215895 57684 232320 57712
rect 215895 57681 215907 57684
rect 215849 57675 215907 57681
rect 232314 57672 232320 57684
rect 232372 57672 232378 57724
rect 233142 57672 233148 57724
rect 233200 57712 233206 57724
rect 250990 57712 250996 57724
rect 233200 57684 250996 57712
rect 233200 57672 233206 57684
rect 250990 57672 250996 57684
rect 251048 57672 251054 57724
rect 255222 57672 255228 57724
rect 255280 57712 255286 57724
rect 269574 57712 269580 57724
rect 255280 57684 269580 57712
rect 255280 57672 255286 57684
rect 269574 57672 269580 57684
rect 269632 57672 269638 57724
rect 271690 57672 271696 57724
rect 271748 57712 271754 57724
rect 282270 57712 282276 57724
rect 271748 57684 282276 57712
rect 271748 57672 271754 57684
rect 282270 57672 282276 57684
rect 282328 57672 282334 57724
rect 284202 57672 284208 57724
rect 284260 57712 284266 57724
rect 293034 57712 293040 57724
rect 284260 57684 293040 57712
rect 284260 57672 284266 57684
rect 293034 57672 293040 57684
rect 293092 57672 293098 57724
rect 296622 57672 296628 57724
rect 296680 57712 296686 57724
rect 302878 57712 302884 57724
rect 296680 57684 302884 57712
rect 296680 57672 296686 57684
rect 302878 57672 302884 57684
rect 302936 57672 302942 57724
rect 310422 57672 310428 57724
rect 310480 57712 310486 57724
rect 314654 57712 314660 57724
rect 310480 57684 314660 57712
rect 310480 57672 310486 57684
rect 314654 57672 314660 57684
rect 314712 57672 314718 57724
rect 321462 57672 321468 57724
rect 321520 57712 321526 57724
rect 323486 57712 323492 57724
rect 321520 57684 323492 57712
rect 321520 57672 321526 57684
rect 323486 57672 323492 57684
rect 323544 57672 323550 57724
rect 466454 57672 466460 57724
rect 466512 57712 466518 57724
rect 494238 57712 494244 57724
rect 466512 57684 494244 57712
rect 466512 57672 466518 57684
rect 494238 57672 494244 57684
rect 494296 57672 494302 57724
rect 496906 57712 496912 57724
rect 494348 57684 496912 57712
rect 173618 57644 173624 57656
rect 140740 57616 147260 57644
rect 147324 57616 173624 57644
rect 140740 57604 140746 57616
rect 31662 57536 31668 57588
rect 31720 57576 31726 57588
rect 85390 57576 85396 57588
rect 31720 57548 85396 57576
rect 31720 57536 31726 57548
rect 85390 57536 85396 57548
rect 85448 57536 85454 57588
rect 89622 57536 89628 57588
rect 89680 57576 89686 57588
rect 119985 57579 120043 57585
rect 119985 57576 119997 57579
rect 89680 57548 119997 57576
rect 89680 57536 89686 57548
rect 119985 57545 119997 57548
rect 120031 57545 120043 57579
rect 119985 57539 120043 57545
rect 120077 57579 120135 57585
rect 120077 57545 120089 57579
rect 120123 57576 120135 57579
rect 122466 57576 122472 57588
rect 120123 57548 122472 57576
rect 120123 57545 120135 57548
rect 120077 57539 120135 57545
rect 122466 57536 122472 57548
rect 122524 57536 122530 57588
rect 122561 57579 122619 57585
rect 122561 57545 122573 57579
rect 122607 57576 122619 57579
rect 130470 57576 130476 57588
rect 122607 57548 130476 57576
rect 122607 57545 122619 57548
rect 122561 57539 122619 57545
rect 130470 57536 130476 57548
rect 130528 57536 130534 57588
rect 130565 57579 130623 57585
rect 130565 57545 130577 57579
rect 130611 57576 130623 57579
rect 133414 57576 133420 57588
rect 130611 57548 133420 57576
rect 130611 57545 130623 57548
rect 130565 57539 130623 57545
rect 133414 57536 133420 57548
rect 133472 57536 133478 57588
rect 141973 57579 142031 57585
rect 141973 57545 141985 57579
rect 142019 57576 142031 57579
rect 147122 57576 147128 57588
rect 142019 57548 147128 57576
rect 142019 57545 142031 57548
rect 141973 57539 142031 57545
rect 147122 57536 147128 57548
rect 147180 57536 147186 57588
rect 23382 57468 23388 57520
rect 23440 57508 23446 57520
rect 78582 57508 78588 57520
rect 23440 57480 78588 57508
rect 23440 57468 23446 57480
rect 78582 57468 78588 57480
rect 78640 57468 78646 57520
rect 83458 57508 83464 57520
rect 79060 57480 83464 57508
rect 21910 57400 21916 57452
rect 21968 57440 21974 57452
rect 76558 57440 76564 57452
rect 21968 57412 76564 57440
rect 21968 57400 21974 57412
rect 76558 57400 76564 57412
rect 76616 57400 76622 57452
rect 77941 57443 77999 57449
rect 77941 57409 77953 57443
rect 77987 57440 77999 57443
rect 79060 57440 79088 57480
rect 83458 57468 83464 57480
rect 83516 57468 83522 57520
rect 83553 57511 83611 57517
rect 83553 57477 83565 57511
rect 83599 57508 83611 57511
rect 86402 57508 86408 57520
rect 83599 57480 86408 57508
rect 83599 57477 83611 57480
rect 83553 57471 83611 57477
rect 86402 57468 86408 57480
rect 86460 57468 86466 57520
rect 86862 57468 86868 57520
rect 86920 57508 86926 57520
rect 94593 57511 94651 57517
rect 86920 57480 94544 57508
rect 86920 57468 86926 57480
rect 77987 57412 79088 57440
rect 79137 57443 79195 57449
rect 77987 57409 77999 57412
rect 77941 57403 77999 57409
rect 79137 57409 79149 57443
rect 79183 57440 79195 57443
rect 81621 57443 81679 57449
rect 81621 57440 81633 57443
rect 79183 57412 81633 57440
rect 79183 57409 79195 57412
rect 79137 57403 79195 57409
rect 81621 57409 81633 57412
rect 81667 57409 81679 57443
rect 81621 57403 81679 57409
rect 82078 57400 82084 57452
rect 82136 57440 82142 57452
rect 92290 57440 92296 57452
rect 82136 57412 92296 57440
rect 82136 57400 82142 57412
rect 92290 57400 92296 57412
rect 92348 57400 92354 57452
rect 94516 57440 94544 57480
rect 94593 57477 94605 57511
rect 94639 57508 94651 57511
rect 129458 57508 129464 57520
rect 94639 57480 129464 57508
rect 94639 57477 94651 57480
rect 94593 57471 94651 57477
rect 129458 57468 129464 57480
rect 129516 57468 129522 57520
rect 129645 57511 129703 57517
rect 129645 57477 129657 57511
rect 129691 57508 129703 57511
rect 132402 57508 132408 57520
rect 129691 57480 132408 57508
rect 129691 57477 129703 57480
rect 129645 57471 129703 57477
rect 132402 57468 132408 57480
rect 132460 57468 132466 57520
rect 132497 57511 132555 57517
rect 132497 57477 132509 57511
rect 132543 57508 132555 57511
rect 145190 57508 145196 57520
rect 132543 57480 145196 57508
rect 132543 57477 132555 57480
rect 132497 57471 132555 57477
rect 145190 57468 145196 57480
rect 145248 57468 145254 57520
rect 122561 57443 122619 57449
rect 122561 57440 122573 57443
rect 94516 57412 122573 57440
rect 122561 57409 122573 57412
rect 122607 57409 122619 57443
rect 122561 57403 122619 57409
rect 124122 57400 124128 57452
rect 124180 57440 124186 57452
rect 132221 57443 132279 57449
rect 132221 57440 132233 57443
rect 124180 57412 132233 57440
rect 124180 57400 124186 57412
rect 132221 57409 132233 57412
rect 132267 57409 132279 57443
rect 132221 57403 132279 57409
rect 136542 57400 136548 57452
rect 136600 57440 136606 57452
rect 147232 57440 147260 57616
rect 173618 57604 173624 57616
rect 173676 57604 173682 57656
rect 176562 57604 176568 57656
rect 176620 57644 176626 57656
rect 203978 57644 203984 57656
rect 176620 57616 203984 57644
rect 176620 57604 176626 57616
rect 203978 57604 203984 57616
rect 204036 57604 204042 57656
rect 204162 57604 204168 57656
rect 204220 57644 204226 57656
rect 227438 57644 227444 57656
rect 204220 57616 227444 57644
rect 204220 57604 204226 57616
rect 227438 57604 227444 57616
rect 227496 57604 227502 57656
rect 229002 57604 229008 57656
rect 229060 57644 229066 57656
rect 247034 57644 247040 57656
rect 229060 57616 247040 57644
rect 229060 57604 229066 57616
rect 247034 57604 247040 57616
rect 247092 57604 247098 57656
rect 252462 57604 252468 57656
rect 252520 57644 252526 57656
rect 266630 57644 266636 57656
rect 252520 57616 266636 57644
rect 252520 57604 252526 57616
rect 266630 57604 266636 57616
rect 266688 57604 266694 57656
rect 267642 57604 267648 57656
rect 267700 57644 267706 57656
rect 279326 57644 279332 57656
rect 267700 57616 279332 57644
rect 267700 57604 267706 57616
rect 279326 57604 279332 57616
rect 279384 57604 279390 57656
rect 281442 57604 281448 57656
rect 281500 57644 281506 57656
rect 291102 57644 291108 57656
rect 281500 57616 291108 57644
rect 281500 57604 281506 57616
rect 291102 57604 291108 57616
rect 291160 57604 291166 57656
rect 311802 57604 311808 57656
rect 311860 57644 311866 57656
rect 315574 57644 315580 57656
rect 311860 57616 315580 57644
rect 311860 57604 311866 57616
rect 315574 57604 315580 57616
rect 315632 57604 315638 57656
rect 316678 57604 316684 57656
rect 316736 57644 316742 57656
rect 317598 57644 317604 57656
rect 316736 57616 317604 57644
rect 316736 57604 316742 57616
rect 317598 57604 317604 57616
rect 317656 57604 317662 57656
rect 322842 57604 322848 57656
rect 322900 57644 322906 57656
rect 325418 57644 325424 57656
rect 322900 57616 325424 57644
rect 322900 57604 322906 57616
rect 325418 57604 325424 57616
rect 325476 57604 325482 57656
rect 328362 57604 328368 57656
rect 328420 57644 328426 57656
rect 329282 57644 329288 57656
rect 328420 57616 329288 57644
rect 328420 57604 328426 57616
rect 329282 57604 329288 57616
rect 329340 57604 329346 57656
rect 344002 57604 344008 57656
rect 344060 57644 344066 57656
rect 344922 57644 344928 57656
rect 344060 57616 344928 57644
rect 344060 57604 344066 57616
rect 344922 57604 344928 57616
rect 344980 57604 344986 57656
rect 346946 57604 346952 57656
rect 347004 57644 347010 57656
rect 347958 57644 347964 57656
rect 347004 57616 347964 57644
rect 347004 57604 347010 57616
rect 347958 57604 347964 57616
rect 348016 57604 348022 57656
rect 350902 57604 350908 57656
rect 350960 57644 350966 57656
rect 351822 57644 351828 57656
rect 350960 57616 351828 57644
rect 350960 57604 350966 57616
rect 351822 57604 351828 57616
rect 351880 57604 351886 57656
rect 357710 57604 357716 57656
rect 357768 57644 357774 57656
rect 358630 57644 358636 57656
rect 357768 57616 358636 57644
rect 357768 57604 357774 57616
rect 358630 57604 358636 57616
rect 358688 57604 358694 57656
rect 360654 57604 360660 57656
rect 360712 57644 360718 57656
rect 362218 57644 362224 57656
rect 360712 57616 362224 57644
rect 360712 57604 360718 57616
rect 362218 57604 362224 57616
rect 362276 57604 362282 57656
rect 367554 57604 367560 57656
rect 367612 57644 367618 57656
rect 368382 57644 368388 57656
rect 367612 57616 368388 57644
rect 367612 57604 367618 57616
rect 368382 57604 368388 57616
rect 368440 57604 368446 57656
rect 368474 57604 368480 57656
rect 368532 57644 368538 57656
rect 369670 57644 369676 57656
rect 368532 57616 369676 57644
rect 368532 57604 368538 57616
rect 369670 57604 369676 57616
rect 369728 57604 369734 57656
rect 374362 57604 374368 57656
rect 374420 57644 374426 57656
rect 375282 57644 375288 57656
rect 374420 57616 375288 57644
rect 374420 57604 374426 57616
rect 375282 57604 375288 57616
rect 375340 57604 375346 57656
rect 375374 57604 375380 57656
rect 375432 57644 375438 57656
rect 376570 57644 376576 57656
rect 375432 57616 376576 57644
rect 375432 57604 375438 57616
rect 376570 57604 376576 57616
rect 376628 57604 376634 57656
rect 379238 57604 379244 57656
rect 379296 57644 379302 57656
rect 380158 57644 380164 57656
rect 379296 57616 380164 57644
rect 379296 57604 379302 57616
rect 380158 57604 380164 57616
rect 380216 57604 380222 57656
rect 381262 57604 381268 57656
rect 381320 57644 381326 57656
rect 382090 57644 382096 57656
rect 381320 57616 382096 57644
rect 381320 57604 381326 57616
rect 382090 57604 382096 57616
rect 382148 57604 382154 57656
rect 388070 57604 388076 57656
rect 388128 57644 388134 57656
rect 389082 57644 389088 57656
rect 388128 57616 389088 57644
rect 388128 57604 388134 57616
rect 389082 57604 389088 57616
rect 389140 57604 389146 57656
rect 391014 57604 391020 57656
rect 391072 57644 391078 57656
rect 391842 57644 391848 57656
rect 391072 57616 391848 57644
rect 391072 57604 391078 57616
rect 391842 57604 391848 57616
rect 391900 57604 391906 57656
rect 392026 57604 392032 57656
rect 392084 57644 392090 57656
rect 393222 57644 393228 57656
rect 392084 57616 393228 57644
rect 392084 57604 392090 57616
rect 393222 57604 393228 57616
rect 393280 57604 393286 57656
rect 394970 57604 394976 57656
rect 395028 57644 395034 57656
rect 395890 57644 395896 57656
rect 395028 57616 395896 57644
rect 395028 57604 395034 57616
rect 395890 57604 395896 57616
rect 395948 57604 395954 57656
rect 397914 57604 397920 57656
rect 397972 57644 397978 57656
rect 398742 57644 398748 57656
rect 397972 57616 398748 57644
rect 397972 57604 397978 57616
rect 398742 57604 398748 57616
rect 398800 57604 398806 57656
rect 398834 57604 398840 57656
rect 398892 57644 398898 57656
rect 400030 57644 400036 57656
rect 398892 57616 400036 57644
rect 398892 57604 398898 57616
rect 400030 57604 400036 57616
rect 400088 57604 400094 57656
rect 401778 57604 401784 57656
rect 401836 57644 401842 57656
rect 402790 57644 402796 57656
rect 401836 57616 402796 57644
rect 401836 57604 401842 57616
rect 402790 57604 402796 57616
rect 402848 57604 402854 57656
rect 404722 57604 404728 57656
rect 404780 57644 404786 57656
rect 405642 57644 405648 57656
rect 404780 57616 405648 57644
rect 404780 57604 404786 57616
rect 405642 57604 405648 57616
rect 405700 57604 405706 57656
rect 408678 57604 408684 57656
rect 408736 57644 408742 57656
rect 409690 57644 409696 57656
rect 408736 57616 409696 57644
rect 408736 57604 408742 57616
rect 409690 57604 409696 57616
rect 409748 57604 409754 57656
rect 411622 57604 411628 57656
rect 411680 57644 411686 57656
rect 412450 57644 412456 57656
rect 411680 57616 412456 57644
rect 411680 57604 411686 57616
rect 412450 57604 412456 57616
rect 412508 57604 412514 57656
rect 418430 57604 418436 57656
rect 418488 57644 418494 57656
rect 419442 57644 419448 57656
rect 418488 57616 419448 57644
rect 418488 57604 418494 57616
rect 419442 57604 419448 57616
rect 419500 57604 419506 57656
rect 421374 57604 421380 57656
rect 421432 57644 421438 57656
rect 422202 57644 422208 57656
rect 421432 57616 422208 57644
rect 421432 57604 421438 57616
rect 422202 57604 422208 57616
rect 422260 57604 422266 57656
rect 422386 57604 422392 57656
rect 422444 57644 422450 57656
rect 423490 57644 423496 57656
rect 422444 57616 423496 57644
rect 422444 57604 422450 57616
rect 423490 57604 423496 57616
rect 423548 57604 423554 57656
rect 425330 57604 425336 57656
rect 425388 57644 425394 57656
rect 426250 57644 426256 57656
rect 425388 57616 426256 57644
rect 425388 57604 425394 57616
rect 426250 57604 426256 57616
rect 426308 57604 426314 57656
rect 428274 57604 428280 57656
rect 428332 57644 428338 57656
rect 429102 57644 429108 57656
rect 428332 57616 429108 57644
rect 428332 57604 428338 57616
rect 429102 57604 429108 57616
rect 429160 57604 429166 57656
rect 432138 57604 432144 57656
rect 432196 57644 432202 57656
rect 433150 57644 433156 57656
rect 432196 57616 433156 57644
rect 432196 57604 432202 57616
rect 433150 57604 433156 57616
rect 433208 57604 433214 57656
rect 435082 57604 435088 57656
rect 435140 57644 435146 57656
rect 436002 57644 436008 57656
rect 435140 57616 436008 57644
rect 435140 57604 435146 57616
rect 436002 57604 436008 57616
rect 436060 57604 436066 57656
rect 439038 57604 439044 57656
rect 439096 57644 439102 57656
rect 440142 57644 440148 57656
rect 439096 57616 440148 57644
rect 439096 57604 439102 57616
rect 440142 57604 440148 57616
rect 440200 57604 440206 57656
rect 441982 57604 441988 57656
rect 442040 57644 442046 57656
rect 442902 57644 442908 57656
rect 442040 57616 442908 57644
rect 442040 57604 442046 57616
rect 442902 57604 442908 57616
rect 442960 57604 442966 57656
rect 448790 57604 448796 57656
rect 448848 57644 448854 57656
rect 449710 57644 449716 57656
rect 448848 57616 449716 57644
rect 448848 57604 448854 57616
rect 449710 57604 449716 57616
rect 449768 57604 449774 57656
rect 451734 57604 451740 57656
rect 451792 57644 451798 57656
rect 452562 57644 452568 57656
rect 451792 57616 452568 57644
rect 451792 57604 451798 57616
rect 452562 57604 452568 57616
rect 452620 57604 452626 57656
rect 452746 57604 452752 57656
rect 452804 57644 452810 57656
rect 453942 57644 453948 57656
rect 452804 57616 453948 57644
rect 452804 57604 452810 57616
rect 453942 57604 453948 57616
rect 454000 57604 454006 57656
rect 455690 57604 455696 57656
rect 455748 57644 455754 57656
rect 456702 57644 456708 57656
rect 455748 57616 456708 57644
rect 455748 57604 455754 57616
rect 456702 57604 456708 57616
rect 456760 57604 456766 57656
rect 458634 57604 458640 57656
rect 458692 57644 458698 57656
rect 459462 57644 459468 57656
rect 458692 57616 459468 57644
rect 458692 57604 458698 57616
rect 459462 57604 459468 57616
rect 459520 57604 459526 57656
rect 459554 57604 459560 57656
rect 459612 57644 459618 57656
rect 460842 57644 460848 57656
rect 459612 57616 460848 57644
rect 459612 57604 459618 57616
rect 460842 57604 460848 57616
rect 460900 57604 460906 57656
rect 462498 57604 462504 57656
rect 462556 57644 462562 57656
rect 463602 57644 463608 57656
rect 462556 57616 463608 57644
rect 462556 57604 462562 57616
rect 463602 57604 463608 57616
rect 463660 57604 463666 57656
rect 465442 57604 465448 57656
rect 465500 57644 465506 57656
rect 466362 57644 466368 57656
rect 465500 57616 466368 57644
rect 465500 57604 465506 57616
rect 466362 57604 466368 57616
rect 466420 57604 466426 57656
rect 469398 57604 469404 57656
rect 469456 57644 469462 57656
rect 494348 57644 494376 57684
rect 496906 57672 496912 57684
rect 496964 57672 496970 57724
rect 512454 57672 512460 57724
rect 512512 57712 512518 57724
rect 547138 57712 547144 57724
rect 512512 57684 547144 57712
rect 512512 57672 512518 57684
rect 547138 57672 547144 57684
rect 547196 57672 547202 57724
rect 469456 57616 494376 57644
rect 469456 57604 469462 57616
rect 496814 57604 496820 57656
rect 496872 57644 496878 57656
rect 498102 57644 498108 57656
rect 496872 57616 498108 57644
rect 496872 57604 496878 57616
rect 498102 57604 498108 57616
rect 498160 57604 498166 57656
rect 499758 57604 499764 57656
rect 499816 57644 499822 57656
rect 500862 57644 500868 57656
rect 499816 57616 500868 57644
rect 499816 57604 499822 57616
rect 500862 57604 500868 57616
rect 500920 57604 500926 57656
rect 502702 57604 502708 57656
rect 502760 57644 502766 57656
rect 503622 57644 503628 57656
rect 502760 57616 503628 57644
rect 502760 57604 502766 57616
rect 503622 57604 503628 57616
rect 503680 57604 503686 57656
rect 505646 57604 505652 57656
rect 505704 57644 505710 57656
rect 506382 57644 506388 57656
rect 505704 57616 506388 57644
rect 505704 57604 505710 57616
rect 506382 57604 506388 57616
rect 506440 57604 506446 57656
rect 513466 57604 513472 57656
rect 513524 57644 513530 57656
rect 514570 57644 514576 57656
rect 513524 57616 514576 57644
rect 513524 57604 513530 57616
rect 514570 57604 514576 57616
rect 514628 57604 514634 57656
rect 515398 57604 515404 57656
rect 515456 57644 515462 57656
rect 549898 57644 549904 57656
rect 515456 57616 549904 57644
rect 515456 57604 515462 57616
rect 549898 57604 549904 57616
rect 549956 57604 549962 57656
rect 151725 57579 151783 57585
rect 151725 57545 151737 57579
rect 151771 57576 151783 57579
rect 176470 57576 176476 57588
rect 151771 57548 176476 57576
rect 151771 57545 151783 57548
rect 151725 57539 151783 57545
rect 176470 57536 176476 57548
rect 176528 57536 176534 57588
rect 176657 57579 176715 57585
rect 176657 57545 176669 57579
rect 176703 57576 176715 57579
rect 183370 57576 183376 57588
rect 176703 57548 183376 57576
rect 176703 57545 176715 57548
rect 176657 57539 176715 57545
rect 183370 57536 183376 57548
rect 183428 57536 183434 57588
rect 184842 57536 184848 57588
rect 184900 57576 184906 57588
rect 191009 57579 191067 57585
rect 191009 57576 191021 57579
rect 184900 57548 191021 57576
rect 184900 57536 184906 57548
rect 191009 57545 191021 57548
rect 191055 57545 191067 57579
rect 191009 57539 191067 57545
rect 191101 57579 191159 57585
rect 191101 57545 191113 57579
rect 191147 57576 191159 57579
rect 208854 57576 208860 57588
rect 191147 57548 208860 57576
rect 191147 57545 191159 57548
rect 191101 57539 191159 57545
rect 208854 57536 208860 57548
rect 208912 57536 208918 57588
rect 211062 57536 211068 57588
rect 211120 57576 211126 57588
rect 233326 57576 233332 57588
rect 211120 57548 233332 57576
rect 211120 57536 211126 57548
rect 233326 57536 233332 57548
rect 233384 57536 233390 57588
rect 237190 57536 237196 57588
rect 237248 57576 237254 57588
rect 254854 57576 254860 57588
rect 237248 57548 254860 57576
rect 237248 57536 237254 57548
rect 254854 57536 254860 57548
rect 254912 57536 254918 57588
rect 256602 57536 256608 57588
rect 256660 57576 256666 57588
rect 270586 57576 270592 57588
rect 256660 57548 270592 57576
rect 256660 57536 256666 57548
rect 270586 57536 270592 57548
rect 270644 57536 270650 57588
rect 273162 57536 273168 57588
rect 273220 57576 273226 57588
rect 284294 57576 284300 57588
rect 273220 57548 284300 57576
rect 273220 57536 273226 57548
rect 284294 57536 284300 57548
rect 284352 57536 284358 57588
rect 286962 57536 286968 57588
rect 287020 57576 287026 57588
rect 295058 57576 295064 57588
rect 287020 57548 295064 57576
rect 287020 57536 287026 57548
rect 295058 57536 295064 57548
rect 295116 57536 295122 57588
rect 309042 57536 309048 57588
rect 309100 57576 309106 57588
rect 313642 57576 313648 57588
rect 309100 57548 313648 57576
rect 309100 57536 309106 57548
rect 313642 57536 313648 57548
rect 313700 57536 313706 57588
rect 317322 57536 317328 57588
rect 317380 57576 317386 57588
rect 320542 57576 320548 57588
rect 317380 57548 320548 57576
rect 317380 57536 317386 57548
rect 320542 57536 320548 57548
rect 320600 57536 320606 57588
rect 322750 57536 322756 57588
rect 322808 57576 322814 57588
rect 324406 57576 324412 57588
rect 322808 57548 324412 57576
rect 322808 57536 322814 57548
rect 324406 57536 324412 57548
rect 324464 57536 324470 57588
rect 349890 57536 349896 57588
rect 349948 57576 349954 57588
rect 352006 57576 352012 57588
rect 349948 57548 352012 57576
rect 349948 57536 349954 57548
rect 352006 57536 352012 57548
rect 352064 57536 352070 57588
rect 361666 57536 361672 57588
rect 361724 57576 361730 57588
rect 362770 57576 362776 57588
rect 361724 57548 362776 57576
rect 361724 57536 361730 57548
rect 362770 57536 362776 57548
rect 362828 57536 362834 57588
rect 364610 57536 364616 57588
rect 364668 57576 364674 57588
rect 369946 57576 369952 57588
rect 364668 57548 369952 57576
rect 364668 57536 364674 57548
rect 369946 57536 369952 57548
rect 370004 57536 370010 57588
rect 378318 57536 378324 57588
rect 378376 57576 378382 57588
rect 379422 57576 379428 57588
rect 378376 57548 379428 57576
rect 378376 57536 378382 57548
rect 379422 57536 379428 57548
rect 379480 57536 379486 57588
rect 429194 57536 429200 57588
rect 429252 57576 429258 57588
rect 430482 57576 430488 57588
rect 429252 57548 430488 57576
rect 429252 57536 429258 57548
rect 430482 57536 430488 57548
rect 430540 57536 430546 57588
rect 473354 57536 473360 57588
rect 473412 57576 473418 57588
rect 474550 57576 474556 57588
rect 473412 57548 474556 57576
rect 473412 57536 473418 57548
rect 474550 57536 474556 57548
rect 474608 57536 474614 57588
rect 475286 57536 475292 57588
rect 475344 57576 475350 57588
rect 503714 57576 503720 57588
rect 475344 57548 503720 57576
rect 475344 57536 475350 57548
rect 503714 57536 503720 57548
rect 503772 57536 503778 57588
rect 506658 57536 506664 57588
rect 506716 57576 506722 57588
rect 506716 57548 538904 57576
rect 506716 57536 506722 57548
rect 147677 57511 147735 57517
rect 147677 57477 147689 57511
rect 147723 57508 147735 57511
rect 177482 57508 177488 57520
rect 147723 57480 177488 57508
rect 147723 57477 147735 57480
rect 147677 57471 147735 57477
rect 177482 57468 177488 57480
rect 177540 57468 177546 57520
rect 185581 57511 185639 57517
rect 185581 57508 185593 57511
rect 177592 57480 185593 57508
rect 174538 57440 174544 57452
rect 136600 57412 142844 57440
rect 147232 57412 174544 57440
rect 136600 57400 136606 57412
rect 15102 57332 15108 57384
rect 15160 57372 15166 57384
rect 64877 57375 64935 57381
rect 64877 57372 64889 57375
rect 15160 57344 64889 57372
rect 15160 57332 15166 57344
rect 64877 57341 64889 57344
rect 64923 57341 64935 57375
rect 64877 57335 64935 57341
rect 64966 57332 64972 57384
rect 65024 57372 65030 57384
rect 65518 57372 65524 57384
rect 65024 57344 65524 57372
rect 65024 57332 65030 57344
rect 65518 57332 65524 57344
rect 65576 57332 65582 57384
rect 65613 57375 65671 57381
rect 65613 57341 65625 57375
rect 65659 57372 65671 57375
rect 70762 57372 70768 57384
rect 65659 57344 70768 57372
rect 65659 57341 65671 57344
rect 65613 57335 65671 57341
rect 70762 57332 70768 57344
rect 70820 57332 70826 57384
rect 71038 57332 71044 57384
rect 71096 57372 71102 57384
rect 79502 57372 79508 57384
rect 71096 57344 79508 57372
rect 71096 57332 71102 57344
rect 79502 57332 79508 57344
rect 79560 57332 79566 57384
rect 82541 57375 82599 57381
rect 82541 57372 82553 57375
rect 79612 57344 82553 57372
rect 12342 57264 12348 57316
rect 12400 57304 12406 57316
rect 68738 57304 68744 57316
rect 12400 57276 68744 57304
rect 12400 57264 12406 57276
rect 68738 57264 68744 57276
rect 68796 57264 68802 57316
rect 71130 57264 71136 57316
rect 71188 57304 71194 57316
rect 75638 57304 75644 57316
rect 71188 57276 75644 57304
rect 71188 57264 71194 57276
rect 75638 57264 75644 57276
rect 75696 57264 75702 57316
rect 75822 57264 75828 57316
rect 75880 57304 75886 57316
rect 79612 57304 79640 57344
rect 82541 57341 82553 57344
rect 82587 57341 82599 57375
rect 82541 57335 82599 57341
rect 82722 57332 82728 57384
rect 82780 57372 82786 57384
rect 119801 57375 119859 57381
rect 119801 57372 119813 57375
rect 82780 57344 119813 57372
rect 82780 57332 82786 57344
rect 119801 57341 119813 57344
rect 119847 57341 119859 57375
rect 124582 57372 124588 57384
rect 119801 57335 119859 57341
rect 119908 57344 124588 57372
rect 75880 57276 79640 57304
rect 75880 57264 75886 57276
rect 79962 57264 79968 57316
rect 80020 57304 80026 57316
rect 119908 57304 119936 57344
rect 124582 57332 124588 57344
rect 124640 57332 124646 57384
rect 126146 57372 126152 57384
rect 124692 57344 126152 57372
rect 80020 57276 119936 57304
rect 119985 57307 120043 57313
rect 80020 57264 80026 57276
rect 119985 57273 119997 57307
rect 120031 57304 120043 57307
rect 124493 57307 124551 57313
rect 124493 57304 124505 57307
rect 120031 57276 124505 57304
rect 120031 57273 120043 57276
rect 119985 57267 120043 57273
rect 124493 57273 124505 57276
rect 124539 57273 124551 57307
rect 124493 57267 124551 57273
rect 13630 57196 13636 57248
rect 13688 57236 13694 57248
rect 64877 57239 64935 57245
rect 64877 57236 64889 57239
rect 13688 57208 64889 57236
rect 13688 57196 13694 57208
rect 64877 57205 64889 57208
rect 64923 57205 64935 57239
rect 64877 57199 64935 57205
rect 64969 57239 65027 57245
rect 64969 57205 64981 57239
rect 65015 57236 65027 57239
rect 71682 57236 71688 57248
rect 65015 57208 71688 57236
rect 65015 57205 65027 57208
rect 64969 57199 65027 57205
rect 71682 57196 71688 57208
rect 71740 57196 71746 57248
rect 73798 57196 73804 57248
rect 73856 57236 73862 57248
rect 74626 57236 74632 57248
rect 73856 57208 74632 57236
rect 73856 57196 73862 57208
rect 74626 57196 74632 57208
rect 74684 57196 74690 57248
rect 75178 57196 75184 57248
rect 75236 57236 75242 57248
rect 82446 57236 82452 57248
rect 75236 57208 82452 57236
rect 75236 57196 75242 57208
rect 82446 57196 82452 57208
rect 82504 57196 82510 57248
rect 82541 57239 82599 57245
rect 82541 57205 82553 57239
rect 82587 57236 82599 57239
rect 115109 57239 115167 57245
rect 115109 57236 115121 57239
rect 82587 57208 115121 57236
rect 82587 57205 82599 57208
rect 82541 57199 82599 57205
rect 115109 57205 115121 57208
rect 115155 57205 115167 57239
rect 115109 57199 115167 57205
rect 115198 57196 115204 57248
rect 115256 57236 115262 57248
rect 118694 57236 118700 57248
rect 115256 57208 118700 57236
rect 115256 57196 115262 57208
rect 118694 57196 118700 57208
rect 118752 57196 118758 57248
rect 119801 57239 119859 57245
rect 119801 57205 119813 57239
rect 119847 57236 119859 57239
rect 124692 57236 124720 57344
rect 126146 57332 126152 57344
rect 126204 57332 126210 57384
rect 126238 57332 126244 57384
rect 126296 57372 126302 57384
rect 139302 57372 139308 57384
rect 126296 57344 139308 57372
rect 126296 57332 126302 57344
rect 139302 57332 139308 57344
rect 139360 57332 139366 57384
rect 142816 57372 142844 57412
rect 174538 57400 174544 57412
rect 174596 57400 174602 57452
rect 175182 57400 175188 57452
rect 175240 57440 175246 57452
rect 177592 57440 177620 57480
rect 185581 57477 185593 57480
rect 185627 57477 185639 57511
rect 185581 57471 185639 57477
rect 195885 57511 195943 57517
rect 195885 57477 195897 57511
rect 195931 57508 195943 57511
rect 211798 57508 211804 57520
rect 195931 57480 211804 57508
rect 195931 57477 195943 57480
rect 195885 57471 195943 57477
rect 211798 57468 211804 57480
rect 211856 57468 211862 57520
rect 211893 57511 211951 57517
rect 211893 57477 211905 57511
rect 211939 57508 211951 57511
rect 218606 57508 218612 57520
rect 211939 57480 218612 57508
rect 211939 57477 211951 57480
rect 211893 57471 211951 57477
rect 218606 57468 218612 57480
rect 218664 57468 218670 57520
rect 219250 57468 219256 57520
rect 219308 57508 219314 57520
rect 240226 57508 240232 57520
rect 219308 57480 240232 57508
rect 219308 57468 219314 57480
rect 240226 57468 240232 57480
rect 240284 57468 240290 57520
rect 241422 57468 241428 57520
rect 241480 57508 241486 57520
rect 257798 57508 257804 57520
rect 241480 57480 257804 57508
rect 241480 57468 241486 57480
rect 257798 57468 257804 57480
rect 257856 57468 257862 57520
rect 260742 57468 260748 57520
rect 260800 57508 260806 57520
rect 273530 57508 273536 57520
rect 260800 57480 273536 57508
rect 260800 57468 260806 57480
rect 273530 57468 273536 57480
rect 273588 57468 273594 57520
rect 277302 57468 277308 57520
rect 277360 57508 277366 57520
rect 287238 57508 287244 57520
rect 277360 57480 287244 57508
rect 277360 57468 277366 57480
rect 287238 57468 287244 57480
rect 287296 57468 287302 57520
rect 289722 57468 289728 57520
rect 289780 57508 289786 57520
rect 298002 57508 298008 57520
rect 289780 57480 298008 57508
rect 289780 57468 289786 57480
rect 298002 57468 298008 57480
rect 298060 57468 298066 57520
rect 299382 57468 299388 57520
rect 299440 57508 299446 57520
rect 305822 57508 305828 57520
rect 299440 57480 305828 57508
rect 299440 57468 299446 57480
rect 305822 57468 305828 57480
rect 305880 57468 305886 57520
rect 306282 57468 306288 57520
rect 306340 57508 306346 57520
rect 311710 57508 311716 57520
rect 306340 57480 311716 57508
rect 306340 57468 306346 57480
rect 311710 57468 311716 57480
rect 311768 57468 311774 57520
rect 320082 57468 320088 57520
rect 320140 57508 320146 57520
rect 322474 57508 322480 57520
rect 320140 57480 322480 57508
rect 320140 57468 320146 57480
rect 322474 57468 322480 57480
rect 322532 57468 322538 57520
rect 478230 57468 478236 57520
rect 478288 57508 478294 57520
rect 507946 57508 507952 57520
rect 478288 57480 507952 57508
rect 478288 57468 478294 57480
rect 507946 57468 507952 57480
rect 508004 57468 508010 57520
rect 509510 57468 509516 57520
rect 509568 57508 509574 57520
rect 538769 57511 538827 57517
rect 538769 57508 538781 57511
rect 509568 57480 538781 57508
rect 509568 57468 509574 57480
rect 538769 57477 538781 57480
rect 538815 57477 538827 57511
rect 538876 57508 538904 57548
rect 538950 57536 538956 57588
rect 539008 57576 539014 57588
rect 544378 57576 544384 57588
rect 539008 57548 544384 57576
rect 539008 57536 539014 57548
rect 544378 57536 544384 57548
rect 544436 57536 544442 57588
rect 542354 57508 542360 57520
rect 538876 57480 542360 57508
rect 538769 57471 538827 57477
rect 542354 57468 542360 57480
rect 542412 57468 542418 57520
rect 175240 57412 177620 57440
rect 175240 57400 175246 57412
rect 177942 57400 177948 57452
rect 178000 57440 178006 57452
rect 205910 57440 205916 57452
rect 178000 57412 205916 57440
rect 178000 57400 178006 57412
rect 205910 57400 205916 57412
rect 205968 57400 205974 57452
rect 206738 57400 206744 57452
rect 206796 57440 206802 57452
rect 229370 57440 229376 57452
rect 206796 57412 229376 57440
rect 206796 57400 206802 57412
rect 229370 57400 229376 57412
rect 229428 57400 229434 57452
rect 230474 57400 230480 57452
rect 230532 57440 230538 57452
rect 248966 57440 248972 57452
rect 230532 57412 248972 57440
rect 230532 57400 230538 57412
rect 248966 57400 248972 57412
rect 249024 57400 249030 57452
rect 251082 57400 251088 57452
rect 251140 57440 251146 57452
rect 265618 57440 265624 57452
rect 251140 57412 265624 57440
rect 251140 57400 251146 57412
rect 265618 57400 265624 57412
rect 265676 57400 265682 57452
rect 266262 57400 266268 57452
rect 266320 57440 266326 57452
rect 278406 57440 278412 57452
rect 266320 57412 278412 57440
rect 266320 57400 266326 57412
rect 278406 57400 278412 57412
rect 278464 57400 278470 57452
rect 282822 57400 282828 57452
rect 282880 57440 282886 57452
rect 292114 57440 292120 57452
rect 282880 57412 292120 57440
rect 282880 57400 282886 57412
rect 292114 57400 292120 57412
rect 292172 57400 292178 57452
rect 292482 57400 292488 57452
rect 292540 57440 292546 57452
rect 299934 57440 299940 57452
rect 292540 57412 299940 57440
rect 292540 57400 292546 57412
rect 299934 57400 299940 57412
rect 299992 57400 299998 57452
rect 472342 57400 472348 57452
rect 472400 57440 472406 57452
rect 501046 57440 501052 57452
rect 472400 57412 501052 57440
rect 472400 57400 472406 57412
rect 501046 57400 501052 57412
rect 501104 57400 501110 57452
rect 507578 57400 507584 57452
rect 507636 57440 507642 57452
rect 543734 57440 543740 57452
rect 507636 57412 543740 57440
rect 507636 57400 507642 57412
rect 543734 57400 543740 57412
rect 543792 57400 543798 57452
rect 171594 57372 171600 57384
rect 142816 57344 171600 57372
rect 171594 57332 171600 57344
rect 171652 57332 171658 57384
rect 173069 57375 173127 57381
rect 173069 57341 173081 57375
rect 173115 57372 173127 57375
rect 176657 57375 176715 57381
rect 176657 57372 176669 57375
rect 173115 57344 176669 57372
rect 173115 57341 173127 57344
rect 173069 57335 173127 57341
rect 176657 57341 176669 57344
rect 176703 57341 176715 57375
rect 176657 57335 176715 57341
rect 179322 57332 179328 57384
rect 179380 57372 179386 57384
rect 185489 57375 185547 57381
rect 185489 57372 185501 57375
rect 179380 57344 185501 57372
rect 179380 57332 179386 57344
rect 185489 57341 185501 57344
rect 185535 57341 185547 57375
rect 185489 57335 185547 57341
rect 185581 57375 185639 57381
rect 185581 57341 185593 57375
rect 185627 57372 185639 57375
rect 202966 57372 202972 57384
rect 185627 57344 202972 57372
rect 185627 57341 185639 57344
rect 185581 57335 185639 57341
rect 202966 57332 202972 57344
rect 203024 57332 203030 57384
rect 205542 57332 205548 57384
rect 205600 57372 205606 57384
rect 228450 57372 228456 57384
rect 205600 57344 228456 57372
rect 205600 57332 205606 57344
rect 228450 57332 228456 57344
rect 228508 57332 228514 57384
rect 230382 57372 230388 57384
rect 228560 57344 230388 57372
rect 124769 57307 124827 57313
rect 124769 57273 124781 57307
rect 124815 57304 124827 57307
rect 129645 57307 129703 57313
rect 129645 57304 129657 57307
rect 124815 57276 129657 57304
rect 124815 57273 124827 57276
rect 124769 57267 124827 57273
rect 129645 57273 129657 57276
rect 129691 57273 129703 57307
rect 161842 57304 161848 57316
rect 129645 57267 129703 57273
rect 129752 57276 161848 57304
rect 119847 57208 124720 57236
rect 119847 57205 119859 57208
rect 119801 57199 119859 57205
rect 125502 57196 125508 57248
rect 125560 57236 125566 57248
rect 129752 57236 129780 57276
rect 161842 57264 161848 57276
rect 161900 57264 161906 57316
rect 168374 57264 168380 57316
rect 168432 57304 168438 57316
rect 169294 57304 169300 57316
rect 168432 57276 169300 57304
rect 168432 57264 168438 57276
rect 169294 57264 169300 57276
rect 169352 57264 169358 57316
rect 169389 57307 169447 57313
rect 169389 57273 169401 57307
rect 169435 57304 169447 57307
rect 194134 57304 194140 57316
rect 169435 57276 194140 57304
rect 169435 57273 169447 57276
rect 169389 57267 169447 57273
rect 194134 57264 194140 57276
rect 194192 57264 194198 57316
rect 200022 57264 200028 57316
rect 200080 57304 200086 57316
rect 223574 57304 223580 57316
rect 200080 57276 223580 57304
rect 200080 57264 200086 57276
rect 223574 57264 223580 57276
rect 223632 57264 223638 57316
rect 224221 57307 224279 57313
rect 224221 57273 224233 57307
rect 224267 57304 224279 57307
rect 228560 57304 228588 57344
rect 230382 57332 230388 57344
rect 230440 57332 230446 57384
rect 231762 57332 231768 57384
rect 231820 57372 231826 57384
rect 249978 57372 249984 57384
rect 231820 57344 249984 57372
rect 231820 57332 231826 57344
rect 249978 57332 249984 57344
rect 250036 57332 250042 57384
rect 253750 57332 253756 57384
rect 253808 57372 253814 57384
rect 268562 57372 268568 57384
rect 253808 57344 268568 57372
rect 253808 57332 253814 57344
rect 268562 57332 268568 57344
rect 268620 57332 268626 57384
rect 271782 57332 271788 57384
rect 271840 57372 271846 57384
rect 283282 57372 283288 57384
rect 271840 57344 283288 57372
rect 271840 57332 271846 57344
rect 283282 57332 283288 57344
rect 283340 57332 283346 57384
rect 285582 57332 285588 57384
rect 285640 57372 285646 57384
rect 294046 57372 294052 57384
rect 285640 57344 294052 57372
rect 285640 57332 285646 57344
rect 294046 57332 294052 57344
rect 294104 57332 294110 57384
rect 295242 57332 295248 57384
rect 295300 57372 295306 57384
rect 301866 57372 301872 57384
rect 295300 57344 301872 57372
rect 295300 57332 295306 57344
rect 301866 57332 301872 57344
rect 301924 57332 301930 57384
rect 304902 57332 304908 57384
rect 304960 57372 304966 57384
rect 309686 57372 309692 57384
rect 304960 57344 309692 57372
rect 304960 57332 304966 57344
rect 309686 57332 309692 57344
rect 309744 57332 309750 57384
rect 384206 57332 384212 57384
rect 384264 57372 384270 57384
rect 384942 57372 384948 57384
rect 384264 57344 384948 57372
rect 384264 57332 384270 57344
rect 384942 57332 384948 57344
rect 385000 57332 385006 57384
rect 414566 57332 414572 57384
rect 414624 57372 414630 57384
rect 415302 57372 415308 57384
rect 414624 57344 415308 57372
rect 414624 57332 414630 57344
rect 415302 57332 415308 57344
rect 415360 57332 415366 57384
rect 444926 57332 444932 57384
rect 444984 57372 444990 57384
rect 445662 57372 445668 57384
rect 444984 57344 445668 57372
rect 444984 57332 444990 57344
rect 445662 57332 445668 57344
rect 445720 57332 445726 57384
rect 457622 57332 457628 57384
rect 457680 57372 457686 57384
rect 483106 57372 483112 57384
rect 457680 57344 483112 57372
rect 457680 57332 457686 57344
rect 483106 57332 483112 57344
rect 483164 57332 483170 57384
rect 484118 57332 484124 57384
rect 484176 57372 484182 57384
rect 514754 57372 514760 57384
rect 484176 57344 514760 57372
rect 484176 57332 484182 57344
rect 514754 57332 514760 57344
rect 514812 57332 514818 57384
rect 516410 57332 516416 57384
rect 516468 57372 516474 57384
rect 554866 57372 554872 57384
rect 516468 57344 554872 57372
rect 516468 57332 516474 57344
rect 554866 57332 554872 57344
rect 554924 57332 554930 57384
rect 224267 57276 228588 57304
rect 224267 57273 224279 57276
rect 224221 57267 224279 57273
rect 228910 57264 228916 57316
rect 228968 57304 228974 57316
rect 248046 57304 248052 57316
rect 228968 57276 248052 57304
rect 228968 57264 228974 57276
rect 248046 57264 248052 57276
rect 248104 57264 248110 57316
rect 248322 57264 248328 57316
rect 248380 57304 248386 57316
rect 263686 57304 263692 57316
rect 248380 57276 263692 57304
rect 248380 57264 248386 57276
rect 263686 57264 263692 57276
rect 263744 57264 263750 57316
rect 264882 57264 264888 57316
rect 264940 57304 264946 57316
rect 277394 57304 277400 57316
rect 264940 57276 277400 57304
rect 264940 57264 264946 57276
rect 277394 57264 277400 57276
rect 277452 57264 277458 57316
rect 278682 57264 278688 57316
rect 278740 57304 278746 57316
rect 288158 57304 288164 57316
rect 278740 57276 288164 57304
rect 278740 57264 278746 57276
rect 288158 57264 288164 57276
rect 288216 57264 288222 57316
rect 288250 57264 288256 57316
rect 288308 57304 288314 57316
rect 296990 57304 296996 57316
rect 288308 57276 296996 57304
rect 288308 57264 288314 57276
rect 296990 57264 296996 57276
rect 297048 57264 297054 57316
rect 298002 57264 298008 57316
rect 298060 57304 298066 57316
rect 304810 57304 304816 57316
rect 298060 57276 304816 57304
rect 298060 57264 298066 57276
rect 304810 57264 304816 57276
rect 304868 57264 304874 57316
rect 306190 57264 306196 57316
rect 306248 57304 306254 57316
rect 310698 57304 310704 57316
rect 306248 57276 310704 57304
rect 306248 57264 306254 57276
rect 310698 57264 310704 57276
rect 310756 57264 310762 57316
rect 463510 57264 463516 57316
rect 463568 57304 463574 57316
rect 490098 57304 490104 57316
rect 463568 57276 490104 57304
rect 463568 57264 463574 57276
rect 490098 57264 490104 57276
rect 490156 57264 490162 57316
rect 492858 57264 492864 57316
rect 492916 57304 492922 57316
rect 525794 57304 525800 57316
rect 492916 57276 525800 57304
rect 492916 57264 492922 57276
rect 525794 57264 525800 57276
rect 525852 57264 525858 57316
rect 528186 57264 528192 57316
rect 528244 57304 528250 57316
rect 566458 57304 566464 57316
rect 528244 57276 566464 57304
rect 528244 57264 528250 57276
rect 566458 57264 566464 57276
rect 566516 57264 566522 57316
rect 125560 57208 129780 57236
rect 132221 57239 132279 57245
rect 125560 57196 125566 57208
rect 132221 57205 132233 57239
rect 132267 57236 132279 57239
rect 160830 57236 160836 57248
rect 132267 57208 160836 57236
rect 132267 57205 132279 57208
rect 132221 57199 132279 57205
rect 160830 57196 160836 57208
rect 160888 57196 160894 57248
rect 168190 57196 168196 57248
rect 168248 57236 168254 57248
rect 198090 57236 198096 57248
rect 168248 57208 198096 57236
rect 168248 57196 168254 57208
rect 198090 57196 198096 57208
rect 198148 57196 198154 57248
rect 198642 57196 198648 57248
rect 198700 57236 198706 57248
rect 222562 57236 222568 57248
rect 198700 57208 222568 57236
rect 198700 57196 198706 57208
rect 222562 57196 222568 57208
rect 222620 57196 222626 57248
rect 223482 57196 223488 57248
rect 223540 57236 223546 57248
rect 243078 57236 243084 57248
rect 223540 57208 243084 57236
rect 223540 57196 223546 57208
rect 243078 57196 243084 57208
rect 243136 57196 243142 57248
rect 244182 57196 244188 57248
rect 244240 57236 244246 57248
rect 259730 57236 259736 57248
rect 244240 57208 259736 57236
rect 244240 57196 244246 57208
rect 259730 57196 259736 57208
rect 259788 57196 259794 57248
rect 263410 57196 263416 57248
rect 263468 57236 263474 57248
rect 276382 57236 276388 57248
rect 263468 57208 276388 57236
rect 263468 57196 263474 57208
rect 276382 57196 276388 57208
rect 276440 57196 276446 57248
rect 279970 57196 279976 57248
rect 280028 57236 280034 57248
rect 290182 57236 290188 57248
rect 280028 57208 290188 57236
rect 280028 57196 280034 57208
rect 290182 57196 290188 57208
rect 290240 57196 290246 57248
rect 293862 57196 293868 57248
rect 293920 57236 293926 57248
rect 300946 57236 300952 57248
rect 293920 57208 300952 57236
rect 293920 57196 293926 57208
rect 300946 57196 300952 57208
rect 301004 57196 301010 57248
rect 315942 57196 315948 57248
rect 316000 57236 316006 57248
rect 319530 57236 319536 57248
rect 316000 57208 319536 57236
rect 316000 57196 316006 57208
rect 319530 57196 319536 57208
rect 319588 57196 319594 57248
rect 354766 57196 354772 57248
rect 354824 57236 354830 57248
rect 355870 57236 355876 57248
rect 354824 57208 355876 57236
rect 354824 57196 354830 57208
rect 355870 57196 355876 57208
rect 355928 57196 355934 57248
rect 385126 57196 385132 57248
rect 385184 57236 385190 57248
rect 386322 57236 386328 57248
rect 385184 57208 386328 57236
rect 385184 57196 385190 57208
rect 386322 57196 386328 57208
rect 386380 57196 386386 57248
rect 415486 57196 415492 57248
rect 415544 57236 415550 57248
rect 416682 57236 416688 57248
rect 415544 57208 416688 57236
rect 415544 57196 415550 57208
rect 416682 57196 416688 57208
rect 416740 57196 416746 57248
rect 437106 57196 437112 57248
rect 437164 57236 437170 57248
rect 458266 57236 458272 57248
rect 437164 57208 458272 57236
rect 437164 57196 437170 57208
rect 458266 57196 458272 57208
rect 458324 57196 458330 57248
rect 479150 57196 479156 57248
rect 479208 57236 479214 57248
rect 480162 57236 480168 57248
rect 479208 57208 480168 57236
rect 479208 57196 479214 57208
rect 480162 57196 480168 57208
rect 480220 57196 480226 57248
rect 481174 57196 481180 57248
rect 481232 57236 481238 57248
rect 512086 57236 512092 57248
rect 481232 57208 512092 57236
rect 481232 57196 481238 57208
rect 512086 57196 512092 57208
rect 512144 57196 512150 57248
rect 525242 57196 525248 57248
rect 525300 57236 525306 57248
rect 564434 57236 564440 57248
rect 525300 57208 564440 57236
rect 525300 57196 525306 57208
rect 564434 57196 564440 57208
rect 564492 57196 564498 57248
rect 37182 57128 37188 57180
rect 37240 57168 37246 57180
rect 89346 57168 89352 57180
rect 37240 57140 89352 57168
rect 37240 57128 37246 57140
rect 89346 57128 89352 57140
rect 89404 57128 89410 57180
rect 91649 57171 91707 57177
rect 91649 57137 91661 57171
rect 91695 57168 91707 57171
rect 97166 57168 97172 57180
rect 91695 57140 97172 57168
rect 91695 57137 91707 57140
rect 91649 57131 91707 57137
rect 97166 57128 97172 57140
rect 97224 57128 97230 57180
rect 102870 57128 102876 57180
rect 102928 57168 102934 57180
rect 105998 57168 106004 57180
rect 102928 57140 106004 57168
rect 102928 57128 102934 57140
rect 105998 57128 106004 57140
rect 106056 57128 106062 57180
rect 107562 57128 107568 57180
rect 107620 57168 107626 57180
rect 141973 57171 142031 57177
rect 141973 57168 141985 57171
rect 107620 57140 141985 57168
rect 107620 57128 107626 57140
rect 141973 57137 141985 57140
rect 142019 57137 142031 57171
rect 141973 57131 142031 57137
rect 142062 57128 142068 57180
rect 142120 57168 142126 57180
rect 151725 57171 151783 57177
rect 151725 57168 151737 57171
rect 142120 57140 151737 57168
rect 142120 57128 142126 57140
rect 151725 57137 151737 57140
rect 151771 57137 151783 57171
rect 151725 57131 151783 57137
rect 153102 57128 153108 57180
rect 153160 57168 153166 57180
rect 156049 57171 156107 57177
rect 156049 57168 156061 57171
rect 153160 57140 156061 57168
rect 153160 57128 153166 57140
rect 156049 57137 156061 57140
rect 156095 57137 156107 57171
rect 156049 57131 156107 57137
rect 157242 57128 157248 57180
rect 157300 57168 157306 57180
rect 188246 57168 188252 57180
rect 157300 57140 188252 57168
rect 157300 57128 157306 57140
rect 188246 57128 188252 57140
rect 188304 57128 188310 57180
rect 188982 57128 188988 57180
rect 189040 57168 189046 57180
rect 191285 57171 191343 57177
rect 191285 57168 191297 57171
rect 189040 57140 191297 57168
rect 189040 57128 189046 57140
rect 191285 57137 191297 57140
rect 191331 57137 191343 57171
rect 191285 57131 191343 57137
rect 195977 57171 196035 57177
rect 195977 57137 195989 57171
rect 196023 57168 196035 57171
rect 220630 57168 220636 57180
rect 196023 57140 220636 57168
rect 196023 57137 196035 57140
rect 195977 57131 196035 57137
rect 220630 57128 220636 57140
rect 220688 57128 220694 57180
rect 220722 57128 220728 57180
rect 220780 57168 220786 57180
rect 241146 57168 241152 57180
rect 220780 57140 241152 57168
rect 220780 57128 220786 57140
rect 241146 57128 241152 57140
rect 241204 57128 241210 57180
rect 246942 57128 246948 57180
rect 247000 57168 247006 57180
rect 262674 57168 262680 57180
rect 247000 57140 262680 57168
rect 247000 57128 247006 57140
rect 262674 57128 262680 57140
rect 262732 57128 262738 57180
rect 269022 57128 269028 57180
rect 269080 57168 269086 57180
rect 280338 57168 280344 57180
rect 269080 57140 280344 57168
rect 269080 57128 269086 57140
rect 280338 57128 280344 57140
rect 280396 57128 280402 57180
rect 494882 57128 494888 57180
rect 494940 57168 494946 57180
rect 526438 57168 526444 57180
rect 494940 57140 526444 57168
rect 494940 57128 494946 57140
rect 526438 57128 526444 57140
rect 526496 57128 526502 57180
rect 529106 57128 529112 57180
rect 529164 57168 529170 57180
rect 537478 57168 537484 57180
rect 529164 57140 537484 57168
rect 529164 57128 529170 57140
rect 537478 57128 537484 57140
rect 537536 57128 537542 57180
rect 538769 57171 538827 57177
rect 538769 57137 538781 57171
rect 538815 57168 538827 57171
rect 545758 57168 545764 57180
rect 538815 57140 545764 57168
rect 538815 57137 538827 57140
rect 538769 57131 538827 57137
rect 545758 57128 545764 57140
rect 545816 57128 545822 57180
rect 45462 57060 45468 57112
rect 45520 57100 45526 57112
rect 96154 57100 96160 57112
rect 45520 57072 96160 57100
rect 45520 57060 45526 57072
rect 96154 57060 96160 57072
rect 96212 57060 96218 57112
rect 102045 57103 102103 57109
rect 102045 57069 102057 57103
rect 102091 57100 102103 57103
rect 112806 57100 112812 57112
rect 102091 57072 112812 57100
rect 102091 57069 102103 57072
rect 102045 57063 102103 57069
rect 112806 57060 112812 57072
rect 112864 57060 112870 57112
rect 117222 57060 117228 57112
rect 117280 57100 117286 57112
rect 154942 57100 154948 57112
rect 117280 57072 154948 57100
rect 117280 57060 117286 57072
rect 154942 57060 154948 57072
rect 155000 57060 155006 57112
rect 156598 57060 156604 57112
rect 156656 57100 156662 57112
rect 159818 57100 159824 57112
rect 156656 57072 159824 57100
rect 156656 57060 156662 57072
rect 159818 57060 159824 57072
rect 159876 57060 159882 57112
rect 160002 57060 160008 57112
rect 160060 57100 160066 57112
rect 191190 57100 191196 57112
rect 160060 57072 191196 57100
rect 160060 57060 160066 57072
rect 191190 57060 191196 57072
rect 191248 57060 191254 57112
rect 193122 57060 193128 57112
rect 193180 57100 193186 57112
rect 217686 57100 217692 57112
rect 193180 57072 217692 57100
rect 193180 57060 193186 57072
rect 217686 57060 217692 57072
rect 217744 57060 217750 57112
rect 219342 57060 219348 57112
rect 219400 57100 219406 57112
rect 239214 57100 239220 57112
rect 219400 57072 239220 57100
rect 219400 57060 219406 57072
rect 239214 57060 239220 57072
rect 239272 57060 239278 57112
rect 242802 57060 242808 57112
rect 242860 57100 242866 57112
rect 258810 57100 258816 57112
rect 242860 57072 258816 57100
rect 242860 57060 242866 57072
rect 258810 57060 258816 57072
rect 258868 57060 258874 57112
rect 262122 57060 262128 57112
rect 262180 57100 262186 57112
rect 274450 57100 274456 57112
rect 262180 57072 274456 57100
rect 262180 57060 262186 57072
rect 274450 57060 274456 57072
rect 274508 57060 274514 57112
rect 297910 57060 297916 57112
rect 297968 57100 297974 57112
rect 303890 57100 303896 57112
rect 297968 57072 303896 57100
rect 297968 57060 297974 57072
rect 303890 57060 303896 57072
rect 303948 57060 303954 57112
rect 353846 57060 353852 57112
rect 353904 57100 353910 57112
rect 356146 57100 356152 57112
rect 353904 57072 356152 57100
rect 353904 57060 353910 57072
rect 356146 57060 356152 57072
rect 356204 57060 356210 57112
rect 405734 57060 405740 57112
rect 405792 57100 405798 57112
rect 406930 57100 406936 57112
rect 405792 57072 406936 57100
rect 405792 57060 405798 57072
rect 406930 57060 406936 57072
rect 406988 57060 406994 57112
rect 436094 57060 436100 57112
rect 436152 57100 436158 57112
rect 437382 57100 437388 57112
rect 436152 57072 437388 57100
rect 436152 57060 436158 57072
rect 437382 57060 437388 57072
rect 437440 57060 437446 57112
rect 445846 57060 445852 57112
rect 445904 57100 445910 57112
rect 446950 57100 446956 57112
rect 445904 57072 446956 57100
rect 445904 57060 445910 57072
rect 446950 57060 446956 57072
rect 447008 57060 447014 57112
rect 490006 57060 490012 57112
rect 490064 57100 490070 57112
rect 521654 57100 521660 57112
rect 490064 57072 521660 57100
rect 490064 57060 490070 57072
rect 521654 57060 521660 57072
rect 521712 57060 521718 57112
rect 526162 57060 526168 57112
rect 526220 57100 526226 57112
rect 533338 57100 533344 57112
rect 526220 57072 533344 57100
rect 526220 57060 526226 57072
rect 533338 57060 533344 57072
rect 533396 57060 533402 57112
rect 50982 56992 50988 57044
rect 51040 57032 51046 57044
rect 101122 57032 101128 57044
rect 51040 57004 101128 57032
rect 51040 56992 51046 57004
rect 101122 56992 101128 57004
rect 101180 56992 101186 57044
rect 105538 56992 105544 57044
rect 105596 57032 105602 57044
rect 117774 57032 117780 57044
rect 105596 57004 117780 57032
rect 105596 56992 105602 57004
rect 117774 56992 117780 57004
rect 117832 56992 117838 57044
rect 117958 56992 117964 57044
rect 118016 57032 118022 57044
rect 119893 57035 119951 57041
rect 119893 57032 119905 57035
rect 118016 57004 119905 57032
rect 118016 56992 118022 57004
rect 119893 57001 119905 57004
rect 119939 57001 119951 57035
rect 119893 56995 119951 57001
rect 119982 56992 119988 57044
rect 120040 57032 120046 57044
rect 157886 57032 157892 57044
rect 120040 57004 157892 57032
rect 120040 56992 120046 57004
rect 157886 56992 157892 57004
rect 157944 56992 157950 57044
rect 159910 56992 159916 57044
rect 159968 57032 159974 57044
rect 190270 57032 190276 57044
rect 159968 57004 190276 57032
rect 159968 56992 159974 57004
rect 190270 56992 190276 57004
rect 190328 56992 190334 57044
rect 191009 57035 191067 57041
rect 191009 57001 191021 57035
rect 191055 57032 191067 57035
rect 195885 57035 195943 57041
rect 195885 57032 195897 57035
rect 191055 57004 195897 57032
rect 191055 57001 191067 57004
rect 191009 56995 191067 57001
rect 195885 57001 195897 57004
rect 195931 57001 195943 57035
rect 195885 56995 195943 57001
rect 197262 56992 197268 57044
rect 197320 57032 197326 57044
rect 212813 57035 212871 57041
rect 212813 57032 212825 57035
rect 197320 57004 212825 57032
rect 197320 56992 197326 57004
rect 212813 57001 212825 57004
rect 212859 57001 212871 57035
rect 212813 56995 212871 57001
rect 217962 56992 217968 57044
rect 218020 57032 218026 57044
rect 238202 57032 238208 57044
rect 218020 57004 238208 57032
rect 218020 56992 218026 57004
rect 238202 56992 238208 57004
rect 238260 56992 238266 57044
rect 238662 56992 238668 57044
rect 238720 57032 238726 57044
rect 255866 57032 255872 57044
rect 238720 57004 255872 57032
rect 238720 56992 238726 57004
rect 255866 56992 255872 57004
rect 255924 56992 255930 57044
rect 270402 56992 270408 57044
rect 270460 57032 270466 57044
rect 281350 57032 281356 57044
rect 270460 57004 281356 57032
rect 270460 56992 270466 57004
rect 281350 56992 281356 57004
rect 281408 56992 281414 57044
rect 495802 56992 495808 57044
rect 495860 57032 495866 57044
rect 528738 57032 528744 57044
rect 495860 57004 528744 57032
rect 495860 56992 495866 57004
rect 528738 56992 528744 57004
rect 528796 56992 528802 57044
rect 46842 56924 46848 56976
rect 46900 56964 46906 56976
rect 91649 56967 91707 56973
rect 91649 56964 91661 56967
rect 46900 56936 91661 56964
rect 46900 56924 46906 56936
rect 91649 56933 91661 56936
rect 91695 56933 91707 56967
rect 91649 56927 91707 56933
rect 91738 56924 91744 56976
rect 91796 56964 91802 56976
rect 98178 56964 98184 56976
rect 91796 56936 98184 56964
rect 91796 56924 91802 56936
rect 98178 56924 98184 56936
rect 98236 56924 98242 56976
rect 99377 56967 99435 56973
rect 99377 56933 99389 56967
rect 99423 56964 99435 56967
rect 102597 56967 102655 56973
rect 102597 56964 102609 56967
rect 99423 56936 102609 56964
rect 99423 56933 99435 56936
rect 99377 56927 99435 56933
rect 102597 56933 102609 56936
rect 102643 56933 102655 56967
rect 102597 56927 102655 56933
rect 102689 56967 102747 56973
rect 102689 56933 102701 56967
rect 102735 56964 102747 56967
rect 108574 56964 108580 56976
rect 102735 56936 108580 56964
rect 102735 56933 102747 56936
rect 102689 56927 102747 56933
rect 108574 56924 108580 56936
rect 108632 56924 108638 56976
rect 111058 56924 111064 56976
rect 111116 56964 111122 56976
rect 115017 56967 115075 56973
rect 115017 56964 115029 56967
rect 111116 56936 115029 56964
rect 111116 56924 111122 56936
rect 115017 56933 115029 56936
rect 115063 56933 115075 56967
rect 115017 56927 115075 56933
rect 115109 56967 115167 56973
rect 115109 56933 115121 56967
rect 115155 56964 115167 56967
rect 121270 56964 121276 56976
rect 115155 56936 121276 56964
rect 115155 56933 115167 56936
rect 115109 56927 115167 56933
rect 121270 56924 121276 56936
rect 121328 56924 121334 56976
rect 121362 56924 121368 56976
rect 121420 56964 121426 56976
rect 158898 56964 158904 56976
rect 121420 56936 158904 56964
rect 121420 56924 121426 56936
rect 158898 56924 158904 56936
rect 158956 56924 158962 56976
rect 165522 56924 165528 56976
rect 165580 56964 165586 56976
rect 195146 56964 195152 56976
rect 165580 56936 195152 56964
rect 165580 56924 165586 56936
rect 195146 56924 195152 56936
rect 195204 56924 195210 56976
rect 202690 56924 202696 56976
rect 202748 56964 202754 56976
rect 225506 56964 225512 56976
rect 202748 56936 225512 56964
rect 202748 56924 202754 56936
rect 225506 56924 225512 56936
rect 225564 56924 225570 56976
rect 227622 56924 227628 56976
rect 227680 56964 227686 56976
rect 246022 56964 246028 56976
rect 227680 56936 246028 56964
rect 227680 56924 227686 56936
rect 246022 56924 246028 56936
rect 246080 56924 246086 56976
rect 249702 56924 249708 56976
rect 249760 56964 249766 56976
rect 264698 56964 264704 56976
rect 249760 56936 264704 56964
rect 249760 56924 249766 56936
rect 264698 56924 264704 56936
rect 264756 56924 264762 56976
rect 288342 56924 288348 56976
rect 288400 56964 288406 56976
rect 295978 56964 295984 56976
rect 288400 56936 295984 56964
rect 288400 56924 288406 56936
rect 295978 56924 295984 56936
rect 296036 56924 296042 56976
rect 345014 56924 345020 56976
rect 345072 56964 345078 56976
rect 346302 56964 346308 56976
rect 345072 56936 346308 56964
rect 345072 56924 345078 56936
rect 346302 56924 346308 56936
rect 346360 56924 346366 56976
rect 476206 56924 476212 56976
rect 476264 56964 476270 56976
rect 477402 56964 477408 56976
rect 476264 56936 477408 56964
rect 476264 56924 476270 56936
rect 477402 56924 477408 56936
rect 477460 56924 477466 56976
rect 486050 56924 486056 56976
rect 486108 56964 486114 56976
rect 491938 56964 491944 56976
rect 486108 56936 491944 56964
rect 486108 56924 486114 56936
rect 491938 56924 491944 56936
rect 491996 56924 492002 56976
rect 534994 56924 535000 56976
rect 535052 56964 535058 56976
rect 538950 56964 538956 56976
rect 535052 56936 538956 56964
rect 535052 56924 535058 56936
rect 538950 56924 538956 56936
rect 539008 56924 539014 56976
rect 61378 56856 61384 56908
rect 61436 56896 61442 56908
rect 62850 56896 62856 56908
rect 61436 56868 62856 56896
rect 61436 56856 61442 56868
rect 62850 56856 62856 56868
rect 62908 56856 62914 56908
rect 62945 56899 63003 56905
rect 62945 56865 62957 56899
rect 62991 56896 63003 56899
rect 107010 56896 107016 56908
rect 62991 56868 107016 56896
rect 62991 56865 63003 56868
rect 62945 56859 63003 56865
rect 107010 56856 107016 56868
rect 107068 56856 107074 56908
rect 114462 56856 114468 56908
rect 114520 56896 114526 56908
rect 153010 56896 153016 56908
rect 114520 56868 153016 56896
rect 114520 56856 114526 56868
rect 153010 56856 153016 56868
rect 153068 56856 153074 56908
rect 164142 56856 164148 56908
rect 164200 56896 164206 56908
rect 169389 56899 169447 56905
rect 169389 56896 169401 56899
rect 164200 56868 169401 56896
rect 164200 56856 164206 56868
rect 169389 56865 169401 56868
rect 169435 56865 169447 56899
rect 169389 56859 169447 56865
rect 172422 56856 172428 56908
rect 172480 56896 172486 56908
rect 201034 56896 201040 56908
rect 172480 56868 201040 56896
rect 172480 56856 172486 56868
rect 201034 56856 201040 56868
rect 201092 56856 201098 56908
rect 201402 56856 201408 56908
rect 201460 56896 201466 56908
rect 224494 56896 224500 56908
rect 201460 56868 224500 56896
rect 201460 56856 201466 56868
rect 224494 56856 224500 56868
rect 224552 56856 224558 56908
rect 224862 56856 224868 56908
rect 224920 56896 224926 56908
rect 244090 56896 244096 56908
rect 224920 56868 244096 56896
rect 224920 56856 224926 56868
rect 244090 56856 244096 56868
rect 244148 56856 244154 56908
rect 245470 56856 245476 56908
rect 245528 56896 245534 56908
rect 260374 56896 260380 56908
rect 245528 56868 260380 56896
rect 245528 56856 245534 56868
rect 260374 56856 260380 56868
rect 260432 56856 260438 56908
rect 307662 56856 307668 56908
rect 307720 56896 307726 56908
rect 312630 56896 312636 56908
rect 307720 56868 312636 56896
rect 307720 56856 307726 56868
rect 312630 56856 312636 56868
rect 312688 56856 312694 56908
rect 53742 56788 53748 56840
rect 53800 56828 53806 56840
rect 103054 56828 103060 56840
rect 53800 56800 103060 56828
rect 53800 56788 53806 56800
rect 103054 56788 103060 56800
rect 103112 56788 103118 56840
rect 112438 56788 112444 56840
rect 112496 56828 112502 56840
rect 128817 56831 128875 56837
rect 128817 56828 128829 56831
rect 112496 56800 128829 56828
rect 112496 56788 112502 56800
rect 128817 56797 128829 56800
rect 128863 56797 128875 56831
rect 128817 56791 128875 56797
rect 135898 56788 135904 56840
rect 135956 56828 135962 56840
rect 135956 56800 142752 56828
rect 135956 56788 135962 56800
rect 57882 56720 57888 56772
rect 57940 56760 57946 56772
rect 62945 56763 63003 56769
rect 62945 56760 62957 56763
rect 57940 56732 62957 56760
rect 57940 56720 57946 56732
rect 62945 56729 62957 56732
rect 62991 56729 63003 56763
rect 62945 56723 63003 56729
rect 64782 56720 64788 56772
rect 64840 56760 64846 56772
rect 102045 56763 102103 56769
rect 102045 56760 102057 56763
rect 64840 56732 102057 56760
rect 64840 56720 64846 56732
rect 102045 56729 102057 56732
rect 102091 56729 102103 56763
rect 102045 56723 102103 56729
rect 102597 56763 102655 56769
rect 102597 56729 102609 56763
rect 102643 56760 102655 56763
rect 102643 56732 104204 56760
rect 102643 56729 102655 56732
rect 102597 56723 102655 56729
rect 61470 56652 61476 56704
rect 61528 56692 61534 56704
rect 66806 56692 66812 56704
rect 61528 56664 66812 56692
rect 61528 56652 61534 56664
rect 66806 56652 66812 56664
rect 66864 56652 66870 56704
rect 67542 56652 67548 56704
rect 67600 56692 67606 56704
rect 69569 56695 69627 56701
rect 69569 56692 69581 56695
rect 67600 56664 69581 56692
rect 67600 56652 67606 56664
rect 69569 56661 69581 56664
rect 69615 56661 69627 56695
rect 102689 56695 102747 56701
rect 102689 56692 102701 56695
rect 69569 56655 69627 56661
rect 69676 56664 102701 56692
rect 60642 56584 60648 56636
rect 60700 56624 60706 56636
rect 69676 56624 69704 56664
rect 102689 56661 102701 56664
rect 102735 56661 102747 56695
rect 102689 56655 102747 56661
rect 102778 56652 102784 56704
rect 102836 56692 102842 56704
rect 104066 56692 104072 56704
rect 102836 56664 104072 56692
rect 102836 56652 102842 56664
rect 104066 56652 104072 56664
rect 104124 56652 104130 56704
rect 104176 56692 104204 56732
rect 108298 56720 108304 56772
rect 108356 56760 108362 56772
rect 109862 56760 109868 56772
rect 108356 56732 109868 56760
rect 108356 56720 108362 56732
rect 109862 56720 109868 56732
rect 109920 56720 109926 56772
rect 119338 56720 119344 56772
rect 119396 56760 119402 56772
rect 141234 56760 141240 56772
rect 119396 56732 141240 56760
rect 119396 56720 119402 56732
rect 141234 56720 141240 56732
rect 141292 56720 141298 56772
rect 114830 56692 114836 56704
rect 104176 56664 114836 56692
rect 114830 56652 114836 56664
rect 114888 56652 114894 56704
rect 115017 56695 115075 56701
rect 115017 56661 115029 56695
rect 115063 56692 115075 56695
rect 120718 56692 120724 56704
rect 115063 56664 120724 56692
rect 115063 56661 115075 56664
rect 115017 56655 115075 56661
rect 120718 56652 120724 56664
rect 120776 56652 120782 56704
rect 122098 56652 122104 56704
rect 122156 56692 122162 56704
rect 142617 56695 142675 56701
rect 142617 56692 142629 56695
rect 122156 56664 142629 56692
rect 122156 56652 122162 56664
rect 142617 56661 142629 56664
rect 142663 56661 142675 56695
rect 142617 56655 142675 56661
rect 60700 56596 69704 56624
rect 69753 56627 69811 56633
rect 60700 56584 60706 56596
rect 69753 56593 69765 56627
rect 69799 56624 69811 56627
rect 99377 56627 99435 56633
rect 99377 56624 99389 56627
rect 69799 56596 99389 56624
rect 69799 56593 69811 56596
rect 69753 56587 69811 56593
rect 99377 56593 99389 56596
rect 99423 56593 99435 56627
rect 99377 56587 99435 56593
rect 109678 56584 109684 56636
rect 109736 56624 109742 56636
rect 115750 56624 115756 56636
rect 109736 56596 115756 56624
rect 109736 56584 109742 56596
rect 115750 56584 115756 56596
rect 115808 56584 115814 56636
rect 122190 56584 122196 56636
rect 122248 56624 122254 56636
rect 128817 56627 128875 56633
rect 122248 56596 128768 56624
rect 122248 56584 122254 56596
rect 77938 56516 77944 56568
rect 77996 56556 78002 56568
rect 79137 56559 79195 56565
rect 79137 56556 79149 56559
rect 77996 56528 79149 56556
rect 77996 56516 78002 56528
rect 79137 56525 79149 56528
rect 79183 56525 79195 56559
rect 128740 56556 128768 56596
rect 128817 56593 128829 56627
rect 128863 56624 128875 56627
rect 135346 56624 135352 56636
rect 128863 56596 135352 56624
rect 128863 56593 128875 56596
rect 128817 56587 128875 56593
rect 135346 56584 135352 56596
rect 135404 56584 135410 56636
rect 142724 56624 142752 56800
rect 143442 56788 143448 56840
rect 143500 56828 143506 56840
rect 147677 56831 147735 56837
rect 147677 56828 147689 56831
rect 143500 56800 147689 56828
rect 143500 56788 143506 56800
rect 147677 56797 147689 56800
rect 147723 56797 147735 56831
rect 147677 56791 147735 56797
rect 168282 56788 168288 56840
rect 168340 56828 168346 56840
rect 197078 56828 197084 56840
rect 168340 56800 197084 56828
rect 168340 56788 168346 56800
rect 197078 56788 197084 56800
rect 197136 56788 197142 56840
rect 209682 56788 209688 56840
rect 209740 56828 209746 56840
rect 231394 56828 231400 56840
rect 209740 56800 231400 56828
rect 209740 56788 209746 56800
rect 231394 56788 231400 56800
rect 231452 56788 231458 56840
rect 234522 56788 234528 56840
rect 234580 56828 234586 56840
rect 251910 56828 251916 56840
rect 234580 56800 251916 56828
rect 234580 56788 234586 56800
rect 251910 56788 251916 56800
rect 251968 56788 251974 56840
rect 253842 56788 253848 56840
rect 253900 56828 253906 56840
rect 267366 56828 267372 56840
rect 253900 56800 267372 56828
rect 253900 56788 253906 56800
rect 267366 56788 267372 56800
rect 267424 56788 267430 56840
rect 536006 56788 536012 56840
rect 536064 56828 536070 56840
rect 536742 56828 536748 56840
rect 536064 56800 536748 56828
rect 536064 56788 536070 56800
rect 536742 56788 536748 56800
rect 536800 56788 536806 56840
rect 171042 56720 171048 56772
rect 171100 56760 171106 56772
rect 199654 56760 199660 56772
rect 171100 56732 199660 56760
rect 171100 56720 171106 56732
rect 199654 56720 199660 56732
rect 199712 56720 199718 56772
rect 211893 56763 211951 56769
rect 211893 56760 211905 56763
rect 208228 56732 211905 56760
rect 142801 56695 142859 56701
rect 142801 56661 142813 56695
rect 142847 56692 142859 56695
rect 144178 56692 144184 56704
rect 142847 56664 144184 56692
rect 142847 56661 142859 56664
rect 142801 56655 142859 56661
rect 144178 56652 144184 56664
rect 144236 56652 144242 56704
rect 148134 56692 148140 56704
rect 144288 56664 148140 56692
rect 144288 56624 144316 56664
rect 148134 56652 148140 56664
rect 148192 56652 148198 56704
rect 169018 56652 169024 56704
rect 169076 56692 169082 56704
rect 171137 56695 171195 56701
rect 171137 56692 171149 56695
rect 169076 56664 171149 56692
rect 169076 56652 169082 56664
rect 171137 56661 171149 56664
rect 171183 56661 171195 56695
rect 171137 56655 171195 56661
rect 185489 56695 185547 56701
rect 185489 56661 185501 56695
rect 185535 56692 185547 56695
rect 206922 56692 206928 56704
rect 185535 56664 206928 56692
rect 185535 56661 185547 56664
rect 185489 56655 185547 56661
rect 206922 56652 206928 56664
rect 206980 56652 206986 56704
rect 142724 56596 144316 56624
rect 145558 56584 145564 56636
rect 145616 56624 145622 56636
rect 154022 56624 154028 56636
rect 145616 56596 154028 56624
rect 145616 56584 145622 56596
rect 154022 56584 154028 56596
rect 154080 56584 154086 56636
rect 160738 56584 160744 56636
rect 160796 56624 160802 56636
rect 162762 56624 162768 56636
rect 160796 56596 162768 56624
rect 160796 56584 160802 56596
rect 162762 56584 162768 56596
rect 162820 56584 162826 56636
rect 164878 56584 164884 56636
rect 164936 56624 164942 56636
rect 173069 56627 173127 56633
rect 173069 56624 173081 56627
rect 164936 56596 173081 56624
rect 164936 56584 164942 56596
rect 173069 56593 173081 56596
rect 173115 56593 173127 56627
rect 173069 56587 173127 56593
rect 173158 56584 173164 56636
rect 173216 56624 173222 56636
rect 192202 56624 192208 56636
rect 173216 56596 192208 56624
rect 173216 56584 173222 56596
rect 192202 56584 192208 56596
rect 192260 56584 192266 56636
rect 194502 56584 194508 56636
rect 194560 56624 194566 56636
rect 208228 56624 208256 56732
rect 211893 56729 211905 56732
rect 211939 56729 211951 56763
rect 211893 56723 211951 56729
rect 212442 56720 212448 56772
rect 212500 56760 212506 56772
rect 234338 56760 234344 56772
rect 212500 56732 234344 56760
rect 212500 56720 212506 56732
rect 234338 56720 234344 56732
rect 234396 56720 234402 56772
rect 235902 56720 235908 56772
rect 235960 56760 235966 56772
rect 252922 56760 252928 56772
rect 235960 56732 252928 56760
rect 235960 56720 235966 56732
rect 252922 56720 252928 56732
rect 252980 56720 252986 56772
rect 302142 56720 302148 56772
rect 302200 56760 302206 56772
rect 307754 56760 307760 56772
rect 302200 56732 307760 56760
rect 302200 56720 302206 56732
rect 307754 56720 307760 56732
rect 307812 56720 307818 56772
rect 313182 56720 313188 56772
rect 313240 56760 313246 56772
rect 316586 56760 316592 56772
rect 313240 56732 316592 56760
rect 313240 56720 313246 56732
rect 316586 56720 316592 56732
rect 316644 56720 316650 56772
rect 208302 56652 208308 56704
rect 208360 56692 208366 56704
rect 224221 56695 224279 56701
rect 224221 56692 224233 56695
rect 208360 56664 224233 56692
rect 208360 56652 208366 56664
rect 224221 56661 224233 56664
rect 224267 56661 224279 56695
rect 224221 56655 224279 56661
rect 226242 56652 226248 56704
rect 226300 56692 226306 56704
rect 245102 56692 245108 56704
rect 226300 56664 245108 56692
rect 226300 56652 226306 56664
rect 245102 56652 245108 56664
rect 245160 56652 245166 56704
rect 303522 56652 303528 56704
rect 303580 56692 303586 56704
rect 308766 56692 308772 56704
rect 303580 56664 308772 56692
rect 303580 56652 303586 56664
rect 308766 56652 308772 56664
rect 308824 56652 308830 56704
rect 315298 56652 315304 56704
rect 315356 56692 315362 56704
rect 318518 56692 318524 56704
rect 315356 56664 318524 56692
rect 315356 56652 315362 56664
rect 318518 56652 318524 56664
rect 318576 56652 318582 56704
rect 324222 56652 324228 56704
rect 324280 56692 324286 56704
rect 326338 56692 326344 56704
rect 324280 56664 326344 56692
rect 324280 56652 324286 56664
rect 326338 56652 326344 56664
rect 326396 56652 326402 56704
rect 342990 56652 342996 56704
rect 343048 56692 343054 56704
rect 343726 56692 343732 56704
rect 343048 56664 343732 56692
rect 343048 56652 343054 56664
rect 343726 56652 343732 56664
rect 343784 56652 343790 56704
rect 504082 56652 504088 56704
rect 504140 56692 504146 56704
rect 509878 56692 509884 56704
rect 504140 56664 509884 56692
rect 504140 56652 504146 56664
rect 509878 56652 509884 56664
rect 509936 56652 509942 56704
rect 523310 56652 523316 56704
rect 523368 56692 523374 56704
rect 524322 56692 524328 56704
rect 523368 56664 524328 56692
rect 523368 56652 523374 56664
rect 524322 56652 524328 56664
rect 524380 56652 524386 56704
rect 194560 56596 208256 56624
rect 194560 56584 194566 56596
rect 210970 56584 210976 56636
rect 211028 56624 211034 56636
rect 215849 56627 215907 56633
rect 215849 56624 215861 56627
rect 211028 56596 215861 56624
rect 211028 56584 211034 56596
rect 215849 56593 215861 56596
rect 215895 56593 215907 56627
rect 215849 56587 215907 56593
rect 216582 56584 216588 56636
rect 216640 56624 216646 56636
rect 237006 56624 237012 56636
rect 216640 56596 237012 56624
rect 216640 56584 216646 56596
rect 237006 56584 237012 56596
rect 237064 56584 237070 56636
rect 291102 56584 291108 56636
rect 291160 56624 291166 56636
rect 298922 56624 298928 56636
rect 291160 56596 298928 56624
rect 291160 56584 291166 56596
rect 298922 56584 298928 56596
rect 298980 56584 298986 56636
rect 304258 56584 304264 56636
rect 304316 56624 304322 56636
rect 306834 56624 306840 56636
rect 304316 56596 306840 56624
rect 304316 56584 304322 56596
rect 306834 56584 306840 56596
rect 306892 56584 306898 56636
rect 327350 56624 327356 56636
rect 326356 56596 327356 56624
rect 326356 56568 326384 56596
rect 327350 56584 327356 56596
rect 327408 56584 327414 56636
rect 336734 56584 336740 56636
rect 336792 56624 336798 56636
rect 337194 56624 337200 56636
rect 336792 56596 337200 56624
rect 336792 56584 336798 56596
rect 337194 56584 337200 56596
rect 337252 56584 337258 56636
rect 338114 56584 338120 56636
rect 338172 56624 338178 56636
rect 338206 56624 338212 56636
rect 338172 56596 338212 56624
rect 338172 56584 338178 56596
rect 338206 56584 338212 56596
rect 338264 56584 338270 56636
rect 537938 56584 537944 56636
rect 537996 56624 538002 56636
rect 540238 56624 540244 56636
rect 537996 56596 540244 56624
rect 537996 56584 538002 56596
rect 540238 56584 540244 56596
rect 540296 56584 540302 56636
rect 130565 56559 130623 56565
rect 130565 56556 130577 56559
rect 128740 56528 130577 56556
rect 79137 56519 79195 56525
rect 130565 56525 130577 56528
rect 130611 56525 130623 56559
rect 130565 56519 130623 56525
rect 171137 56559 171195 56565
rect 171137 56525 171149 56559
rect 171183 56556 171195 56559
rect 186314 56556 186320 56568
rect 171183 56528 186320 56556
rect 171183 56525 171195 56528
rect 171137 56519 171195 56525
rect 186314 56516 186320 56528
rect 186372 56516 186378 56568
rect 326338 56516 326344 56568
rect 326396 56516 326402 56568
rect 336734 56448 336740 56500
rect 336792 56488 336798 56500
rect 336792 56460 336837 56488
rect 336792 56448 336798 56460
rect 165614 55836 165620 55888
rect 165672 55876 165678 55888
rect 166350 55876 166356 55888
rect 165672 55848 166356 55876
rect 165672 55836 165678 55848
rect 166350 55836 166356 55848
rect 166408 55836 166414 55888
rect 334161 55607 334219 55613
rect 334161 55573 334173 55607
rect 334207 55604 334219 55607
rect 334342 55604 334348 55616
rect 334207 55576 334348 55604
rect 334207 55573 334219 55576
rect 334161 55567 334219 55573
rect 334342 55564 334348 55576
rect 334400 55564 334406 55616
rect 100849 52343 100907 52349
rect 100849 52309 100861 52343
rect 100895 52340 100907 52343
rect 101214 52340 101220 52352
rect 100895 52312 101220 52340
rect 100895 52309 100907 52312
rect 100849 52303 100907 52309
rect 101214 52300 101220 52312
rect 101272 52300 101278 52352
rect 121549 51595 121607 51601
rect 121549 51561 121561 51595
rect 121595 51592 121607 51595
rect 121730 51592 121736 51604
rect 121595 51564 121736 51592
rect 121595 51561 121607 51564
rect 121549 51555 121607 51561
rect 121730 51552 121736 51564
rect 121788 51552 121794 51604
rect 98546 48328 98552 48340
rect 98507 48300 98552 48328
rect 98546 48288 98552 48300
rect 98604 48288 98610 48340
rect 100846 48328 100852 48340
rect 100807 48300 100852 48328
rect 100846 48288 100852 48300
rect 100904 48288 100910 48340
rect 121546 48328 121552 48340
rect 121507 48300 121552 48328
rect 121546 48288 121552 48300
rect 121604 48288 121610 48340
rect 128998 48288 129004 48340
rect 129056 48328 129062 48340
rect 132497 48331 132555 48337
rect 132497 48328 132509 48331
rect 129056 48300 132509 48328
rect 129056 48288 129062 48300
rect 132497 48297 132509 48300
rect 132543 48297 132555 48331
rect 132497 48291 132555 48297
rect 145190 48288 145196 48340
rect 145248 48328 145254 48340
rect 145282 48328 145288 48340
rect 145248 48300 145288 48328
rect 145248 48288 145254 48300
rect 145282 48288 145288 48300
rect 145340 48288 145346 48340
rect 195882 48288 195888 48340
rect 195940 48328 195946 48340
rect 195977 48331 196035 48337
rect 195977 48328 195989 48331
rect 195940 48300 195989 48328
rect 195940 48288 195946 48300
rect 195977 48297 195989 48300
rect 196023 48297 196035 48331
rect 195977 48291 196035 48297
rect 212626 48288 212632 48340
rect 212684 48328 212690 48340
rect 213454 48328 213460 48340
rect 212684 48300 213460 48328
rect 212684 48288 212690 48300
rect 213454 48288 213460 48300
rect 213512 48288 213518 48340
rect 334158 48328 334164 48340
rect 334119 48300 334164 48328
rect 334158 48288 334164 48300
rect 334216 48288 334222 48340
rect 98638 48220 98644 48272
rect 98696 48260 98702 48272
rect 100110 48260 100116 48272
rect 98696 48232 100116 48260
rect 98696 48220 98702 48232
rect 100110 48220 100116 48232
rect 100168 48220 100174 48272
rect 98546 46968 98552 46980
rect 98507 46940 98552 46968
rect 98546 46928 98552 46940
rect 98604 46928 98610 46980
rect 336734 46928 336740 46980
rect 336792 46968 336798 46980
rect 336792 46940 336837 46968
rect 336792 46928 336798 46940
rect 338114 46900 338120 46912
rect 338075 46872 338120 46900
rect 338114 46860 338120 46872
rect 338172 46860 338178 46912
rect 121454 41352 121460 41404
rect 121512 41392 121518 41404
rect 121638 41392 121644 41404
rect 121512 41364 121644 41392
rect 121512 41352 121518 41364
rect 121638 41352 121644 41364
rect 121696 41352 121702 41404
rect 212534 41352 212540 41404
rect 212592 41392 212598 41404
rect 212718 41392 212724 41404
rect 212592 41364 212724 41392
rect 212592 41352 212598 41364
rect 212718 41352 212724 41364
rect 212776 41352 212782 41404
rect 145006 38632 145012 38684
rect 145064 38672 145070 38684
rect 145098 38672 145104 38684
rect 145064 38644 145104 38672
rect 145064 38632 145070 38644
rect 145098 38632 145104 38644
rect 145156 38632 145162 38684
rect 101030 38604 101036 38616
rect 100991 38576 101036 38604
rect 101030 38564 101036 38576
rect 101088 38564 101094 38616
rect 192021 38607 192079 38613
rect 192021 38573 192033 38607
rect 192067 38604 192079 38607
rect 192110 38604 192116 38616
rect 192067 38576 192116 38604
rect 192067 38573 192079 38576
rect 192021 38567 192079 38573
rect 192110 38564 192116 38576
rect 192168 38564 192174 38616
rect 195882 38604 195888 38616
rect 195843 38576 195888 38604
rect 195882 38564 195888 38576
rect 195940 38564 195946 38616
rect 98270 37952 98276 38004
rect 98328 37992 98334 38004
rect 98454 37992 98460 38004
rect 98328 37964 98460 37992
rect 98328 37952 98334 37964
rect 98454 37952 98460 37964
rect 98512 37952 98518 38004
rect 338114 37312 338120 37324
rect 338075 37284 338120 37312
rect 338114 37272 338120 37284
rect 338172 37272 338178 37324
rect 128633 37247 128691 37253
rect 128633 37213 128645 37247
rect 128679 37244 128691 37247
rect 128814 37244 128820 37256
rect 128679 37216 128820 37244
rect 128679 37213 128691 37216
rect 128633 37207 128691 37213
rect 128814 37204 128820 37216
rect 128872 37204 128878 37256
rect 336734 37204 336740 37256
rect 336792 37244 336798 37256
rect 336792 37216 336837 37244
rect 336792 37204 336798 37216
rect 145006 35748 145012 35760
rect 144967 35720 145012 35748
rect 145006 35708 145012 35720
rect 145064 35708 145070 35760
rect 121638 31764 121644 31816
rect 121696 31764 121702 31816
rect 333974 31764 333980 31816
rect 334032 31764 334038 31816
rect 101033 31671 101091 31677
rect 101033 31637 101045 31671
rect 101079 31668 101091 31671
rect 101214 31668 101220 31680
rect 101079 31640 101220 31668
rect 101079 31637 101091 31640
rect 101033 31631 101091 31637
rect 101214 31628 101220 31640
rect 101272 31628 101278 31680
rect 121656 31668 121684 31764
rect 121730 31668 121736 31680
rect 121656 31640 121736 31668
rect 121730 31628 121736 31640
rect 121788 31628 121794 31680
rect 333992 31668 334020 31764
rect 334066 31668 334072 31680
rect 333992 31640 334072 31668
rect 334066 31628 334072 31640
rect 334124 31628 334130 31680
rect 145009 29019 145067 29025
rect 145009 28985 145021 29019
rect 145055 29016 145067 29019
rect 145190 29016 145196 29028
rect 145055 28988 145196 29016
rect 145055 28985 145067 28988
rect 145009 28979 145067 28985
rect 145190 28976 145196 28988
rect 145248 28976 145254 29028
rect 192018 29016 192024 29028
rect 191979 28988 192024 29016
rect 192018 28976 192024 28988
rect 192076 28976 192082 29028
rect 195882 29016 195888 29028
rect 195843 28988 195888 29016
rect 195882 28976 195888 28988
rect 195940 28976 195946 29028
rect 97994 28908 98000 28960
rect 98052 28948 98058 28960
rect 98454 28948 98460 28960
rect 98052 28920 98460 28948
rect 98052 28908 98058 28920
rect 98454 28908 98460 28920
rect 98512 28908 98518 28960
rect 100754 28908 100760 28960
rect 100812 28948 100818 28960
rect 101214 28948 101220 28960
rect 100812 28920 101220 28948
rect 100812 28908 100818 28920
rect 101214 28908 101220 28920
rect 101272 28908 101278 28960
rect 128630 27724 128636 27736
rect 128591 27696 128636 27724
rect 128630 27684 128636 27696
rect 128688 27684 128694 27736
rect 336734 27616 336740 27668
rect 336792 27656 336798 27668
rect 336792 27628 336837 27656
rect 336792 27616 336798 27628
rect 121641 27591 121699 27597
rect 121641 27557 121653 27591
rect 121687 27588 121699 27591
rect 121730 27588 121736 27600
rect 121687 27560 121736 27588
rect 121687 27557 121699 27560
rect 121641 27551 121699 27557
rect 121730 27548 121736 27560
rect 121788 27548 121794 27600
rect 128630 27548 128636 27600
rect 128688 27588 128694 27600
rect 128909 27591 128967 27597
rect 128909 27588 128921 27591
rect 128688 27560 128921 27588
rect 128688 27548 128694 27560
rect 128909 27557 128921 27560
rect 128955 27557 128967 27591
rect 212534 27588 212540 27600
rect 212495 27560 212540 27588
rect 128909 27551 128967 27557
rect 212534 27548 212540 27560
rect 212592 27548 212598 27600
rect 338114 27588 338120 27600
rect 338075 27560 338120 27588
rect 338114 27548 338120 27560
rect 338172 27548 338178 27600
rect 2866 22040 2872 22092
rect 2924 22080 2930 22092
rect 538030 22080 538036 22092
rect 2924 22052 538036 22080
rect 2924 22040 2930 22052
rect 538030 22040 538036 22052
rect 538088 22040 538094 22092
rect 195882 19456 195888 19508
rect 195940 19456 195946 19508
rect 195900 19372 195928 19456
rect 145006 19320 145012 19372
rect 145064 19360 145070 19372
rect 145098 19360 145104 19372
rect 145064 19332 145104 19360
rect 145064 19320 145070 19332
rect 145098 19320 145104 19332
rect 145156 19320 145162 19372
rect 195882 19320 195888 19372
rect 195940 19320 195946 19372
rect 192202 19292 192208 19304
rect 192163 19264 192208 19292
rect 192202 19252 192208 19264
rect 192260 19252 192266 19304
rect 128906 19224 128912 19236
rect 128867 19196 128912 19224
rect 128906 19184 128912 19196
rect 128964 19184 128970 19236
rect 121638 18000 121644 18012
rect 121599 17972 121644 18000
rect 121638 17960 121644 17972
rect 121696 17960 121702 18012
rect 212537 18003 212595 18009
rect 212537 17969 212549 18003
rect 212583 18000 212595 18003
rect 212626 18000 212632 18012
rect 212583 17972 212632 18000
rect 212583 17969 212595 17972
rect 212537 17963 212595 17969
rect 212626 17960 212632 17972
rect 212684 17960 212690 18012
rect 333974 17932 333980 17944
rect 333935 17904 333980 17932
rect 333974 17892 333980 17904
rect 334032 17892 334038 17944
rect 336734 17892 336740 17944
rect 336792 17932 336798 17944
rect 336792 17904 336837 17932
rect 336792 17892 336798 17904
rect 538858 17892 538864 17944
rect 538916 17932 538922 17944
rect 579798 17932 579804 17944
rect 538916 17904 579804 17932
rect 538916 17892 538922 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 203702 13132 203708 13184
rect 203760 13172 203766 13184
rect 204162 13172 204168 13184
rect 203760 13144 204168 13172
rect 203760 13132 203766 13144
rect 204162 13132 204168 13144
rect 204220 13132 204226 13184
rect 121638 12492 121644 12504
rect 121564 12464 121644 12492
rect 121564 12436 121592 12464
rect 121638 12452 121644 12464
rect 121696 12452 121702 12504
rect 128906 12452 128912 12504
rect 128964 12452 128970 12504
rect 121546 12384 121552 12436
rect 121604 12384 121610 12436
rect 128924 12368 128952 12452
rect 128906 12316 128912 12368
rect 128964 12316 128970 12368
rect 192205 9707 192263 9713
rect 192205 9673 192217 9707
rect 192251 9704 192263 9707
rect 192294 9704 192300 9716
rect 192251 9676 192300 9704
rect 192251 9673 192263 9676
rect 192205 9667 192263 9673
rect 192294 9664 192300 9676
rect 192352 9664 192358 9716
rect 338117 9707 338175 9713
rect 338117 9673 338129 9707
rect 338163 9704 338175 9707
rect 338298 9704 338304 9716
rect 338163 9676 338304 9704
rect 338163 9673 338175 9676
rect 338117 9667 338175 9673
rect 338298 9664 338304 9676
rect 338356 9664 338362 9716
rect 195609 9639 195667 9645
rect 195609 9605 195621 9639
rect 195655 9636 195667 9639
rect 195882 9636 195888 9648
rect 195655 9608 195888 9636
rect 195655 9605 195667 9608
rect 195609 9599 195667 9605
rect 195882 9596 195888 9608
rect 195940 9596 195946 9648
rect 212442 9636 212448 9648
rect 212403 9608 212448 9636
rect 212442 9596 212448 9608
rect 212500 9596 212506 9648
rect 336737 9571 336795 9577
rect 336737 9537 336749 9571
rect 336783 9568 336795 9571
rect 337102 9568 337108 9580
rect 336783 9540 337108 9568
rect 336783 9537 336795 9540
rect 336737 9531 336795 9537
rect 337102 9528 337108 9540
rect 337160 9528 337166 9580
rect 333977 8347 334035 8353
rect 333977 8313 333989 8347
rect 334023 8344 334035 8347
rect 334066 8344 334072 8356
rect 334023 8316 334072 8344
rect 334023 8313 334035 8316
rect 333977 8307 334035 8313
rect 334066 8304 334072 8316
rect 334124 8304 334130 8356
rect 106277 6375 106335 6381
rect 106277 6341 106289 6375
rect 106323 6372 106335 6375
rect 111058 6372 111064 6384
rect 106323 6344 111064 6372
rect 106323 6341 106335 6344
rect 106277 6335 106335 6341
rect 111058 6332 111064 6344
rect 111116 6332 111122 6384
rect 94498 6196 94504 6248
rect 94556 6236 94562 6248
rect 136634 6236 136640 6248
rect 94556 6208 136640 6236
rect 94556 6196 94562 6208
rect 136634 6196 136640 6208
rect 136692 6196 136698 6248
rect 87322 6128 87328 6180
rect 87380 6168 87386 6180
rect 131206 6168 131212 6180
rect 87380 6140 131212 6168
rect 87380 6128 87386 6140
rect 131206 6128 131212 6140
rect 131264 6128 131270 6180
rect 51626 5448 51632 5500
rect 51684 5488 51690 5500
rect 100938 5488 100944 5500
rect 51684 5460 100944 5488
rect 51684 5448 51690 5460
rect 100938 5448 100944 5460
rect 100996 5448 101002 5500
rect 105170 5448 105176 5500
rect 105228 5488 105234 5500
rect 145098 5488 145104 5500
rect 105228 5460 145104 5488
rect 105228 5448 105234 5460
rect 145098 5448 145104 5460
rect 145156 5448 145162 5500
rect 521378 5448 521384 5500
rect 521436 5488 521442 5500
rect 521562 5488 521568 5500
rect 521436 5460 521568 5488
rect 521436 5448 521442 5460
rect 521562 5448 521568 5460
rect 521620 5448 521626 5500
rect 58802 5380 58808 5432
rect 58860 5420 58866 5432
rect 107746 5420 107752 5432
rect 58860 5392 107752 5420
rect 58860 5380 58866 5392
rect 107746 5380 107752 5392
rect 107804 5380 107810 5432
rect 48130 5312 48136 5364
rect 48188 5352 48194 5364
rect 98178 5352 98184 5364
rect 48188 5324 98184 5352
rect 48188 5312 48194 5324
rect 98178 5312 98184 5324
rect 98236 5312 98242 5364
rect 101582 5312 101588 5364
rect 101640 5352 101646 5364
rect 142338 5352 142344 5364
rect 101640 5324 142344 5352
rect 101640 5312 101646 5324
rect 142338 5312 142344 5324
rect 142396 5312 142402 5364
rect 30282 5244 30288 5296
rect 30340 5284 30346 5296
rect 84286 5284 84292 5296
rect 30340 5256 84292 5284
rect 30340 5244 30346 5256
rect 84286 5244 84292 5256
rect 84344 5244 84350 5296
rect 90910 5244 90916 5296
rect 90968 5284 90974 5296
rect 133874 5284 133880 5296
rect 90968 5256 133880 5284
rect 90968 5244 90974 5256
rect 133874 5244 133880 5256
rect 133932 5244 133938 5296
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 69014 5216 69020 5228
rect 12492 5188 69020 5216
rect 12492 5176 12498 5188
rect 69014 5176 69020 5188
rect 69072 5176 69078 5228
rect 76650 5176 76656 5228
rect 76708 5216 76714 5228
rect 121546 5216 121552 5228
rect 76708 5188 121552 5216
rect 76708 5176 76714 5188
rect 121546 5176 121552 5188
rect 121604 5176 121610 5228
rect 155126 5176 155132 5228
rect 155184 5216 155190 5228
rect 186406 5216 186412 5228
rect 155184 5188 186412 5216
rect 155184 5176 155190 5188
rect 186406 5176 186412 5188
rect 186464 5176 186470 5228
rect 502242 5176 502248 5228
rect 502300 5216 502306 5228
rect 536926 5216 536932 5228
rect 502300 5188 536932 5216
rect 502300 5176 502306 5188
rect 536926 5176 536932 5188
rect 536984 5176 536990 5228
rect 22002 5108 22008 5160
rect 22060 5148 22066 5160
rect 77386 5148 77392 5160
rect 22060 5120 77392 5148
rect 22060 5108 22066 5120
rect 77386 5108 77392 5120
rect 77444 5108 77450 5160
rect 80238 5108 80244 5160
rect 80296 5148 80302 5160
rect 125594 5148 125600 5160
rect 80296 5120 125600 5148
rect 80296 5108 80302 5120
rect 125594 5108 125600 5120
rect 125652 5108 125658 5160
rect 148042 5108 148048 5160
rect 148100 5148 148106 5160
rect 180794 5148 180800 5160
rect 148100 5120 180800 5148
rect 148100 5108 148106 5120
rect 180794 5108 180800 5120
rect 180852 5108 180858 5160
rect 505002 5108 505008 5160
rect 505060 5148 505066 5160
rect 540514 5148 540520 5160
rect 505060 5120 540520 5148
rect 505060 5108 505066 5120
rect 540514 5108 540520 5120
rect 540572 5108 540578 5160
rect 17218 5040 17224 5092
rect 17276 5080 17282 5092
rect 73154 5080 73160 5092
rect 17276 5052 73160 5080
rect 17276 5040 17282 5052
rect 73154 5040 73160 5052
rect 73212 5040 73218 5092
rect 83826 5040 83832 5092
rect 83884 5080 83890 5092
rect 128446 5080 128452 5092
rect 83884 5052 128452 5080
rect 83884 5040 83890 5052
rect 128446 5040 128452 5052
rect 128504 5040 128510 5092
rect 134886 5040 134892 5092
rect 134944 5080 134950 5092
rect 169754 5080 169760 5092
rect 134944 5052 169760 5080
rect 134944 5040 134950 5052
rect 169754 5040 169760 5052
rect 169812 5040 169818 5092
rect 510522 5040 510528 5092
rect 510580 5080 510586 5092
rect 547690 5080 547696 5092
rect 510580 5052 547696 5080
rect 510580 5040 510586 5052
rect 547690 5040 547696 5052
rect 547748 5040 547754 5092
rect 2866 4972 2872 5024
rect 2924 5012 2930 5024
rect 60734 5012 60740 5024
rect 2924 4984 60740 5012
rect 2924 4972 2930 4984
rect 60734 4972 60740 4984
rect 60792 4972 60798 5024
rect 69474 4972 69480 5024
rect 69532 5012 69538 5024
rect 115934 5012 115940 5024
rect 69532 4984 115940 5012
rect 69532 4972 69538 4984
rect 115934 4972 115940 4984
rect 115992 4972 115998 5024
rect 131390 4972 131396 5024
rect 131448 5012 131454 5024
rect 166994 5012 167000 5024
rect 131448 4984 167000 5012
rect 131448 4972 131454 4984
rect 166994 4972 167000 4984
rect 167052 4972 167058 5024
rect 514570 4972 514576 5024
rect 514628 5012 514634 5024
rect 551186 5012 551192 5024
rect 514628 4984 551192 5012
rect 514628 4972 514634 4984
rect 551186 4972 551192 4984
rect 551244 4972 551250 5024
rect 7650 4904 7656 4956
rect 7708 4944 7714 4956
rect 64966 4944 64972 4956
rect 7708 4916 64972 4944
rect 7708 4904 7714 4916
rect 64966 4904 64972 4916
rect 65024 4904 65030 4956
rect 73062 4904 73068 4956
rect 73120 4944 73126 4956
rect 118786 4944 118792 4956
rect 73120 4916 118792 4944
rect 73120 4904 73126 4916
rect 118786 4904 118792 4916
rect 118844 4904 118850 4956
rect 132586 4904 132592 4956
rect 132644 4944 132650 4956
rect 168466 4944 168472 4956
rect 132644 4916 168472 4944
rect 132644 4904 132650 4916
rect 168466 4904 168472 4916
rect 168524 4904 168530 4956
rect 520182 4904 520188 4956
rect 520240 4944 520246 4956
rect 558362 4944 558368 4956
rect 520240 4916 558368 4944
rect 520240 4904 520246 4916
rect 558362 4904 558368 4916
rect 558420 4904 558426 4956
rect 566 4836 572 4888
rect 624 4876 630 4888
rect 59354 4876 59360 4888
rect 624 4848 59360 4876
rect 624 4836 630 4848
rect 59354 4836 59360 4848
rect 59412 4836 59418 4888
rect 65978 4836 65984 4888
rect 66036 4876 66042 4888
rect 113174 4876 113180 4888
rect 66036 4848 113180 4876
rect 66036 4836 66042 4848
rect 113174 4836 113180 4848
rect 113232 4836 113238 4888
rect 127802 4836 127808 4888
rect 127860 4876 127866 4888
rect 164234 4876 164240 4888
rect 127860 4848 164240 4876
rect 127860 4836 127866 4848
rect 164234 4836 164240 4848
rect 164292 4836 164298 4888
rect 522942 4836 522948 4888
rect 523000 4876 523006 4888
rect 561950 4876 561956 4888
rect 523000 4848 561956 4876
rect 523000 4836 523006 4848
rect 561950 4836 561956 4848
rect 562008 4836 562014 4888
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 60826 4808 60832 4820
rect 1728 4780 60832 4808
rect 1728 4768 1734 4780
rect 60826 4768 60832 4780
rect 60884 4768 60890 4820
rect 62390 4768 62396 4820
rect 62448 4808 62454 4820
rect 110414 4808 110420 4820
rect 62448 4780 110420 4808
rect 62448 4768 62454 4780
rect 110414 4768 110420 4780
rect 110472 4768 110478 4820
rect 128998 4768 129004 4820
rect 129056 4808 129062 4820
rect 165706 4808 165712 4820
rect 129056 4780 165712 4808
rect 129056 4768 129062 4780
rect 165706 4768 165712 4780
rect 165764 4768 165770 4820
rect 487062 4768 487068 4820
rect 487120 4808 487126 4820
rect 519078 4808 519084 4820
rect 487120 4780 519084 4808
rect 487120 4768 487126 4780
rect 519078 4768 519084 4780
rect 519136 4768 519142 4820
rect 531130 4768 531136 4820
rect 531188 4808 531194 4820
rect 572622 4808 572628 4820
rect 531188 4780 572628 4808
rect 531188 4768 531194 4780
rect 572622 4768 572628 4780
rect 572680 4768 572686 4820
rect 55214 4700 55220 4752
rect 55272 4740 55278 4752
rect 104986 4740 104992 4752
rect 55272 4712 104992 4740
rect 55272 4700 55278 4712
rect 104986 4700 104992 4712
rect 105044 4700 105050 4752
rect 98086 4632 98092 4684
rect 98144 4672 98150 4684
rect 139394 4672 139400 4684
rect 98144 4644 139400 4672
rect 98144 4632 98150 4644
rect 139394 4632 139400 4644
rect 139452 4632 139458 4684
rect 55217 4267 55275 4273
rect 55217 4233 55229 4267
rect 55263 4264 55275 4267
rect 64785 4267 64843 4273
rect 64785 4264 64797 4267
rect 55263 4236 64797 4264
rect 55263 4233 55275 4236
rect 55217 4227 55275 4233
rect 64785 4233 64797 4236
rect 64831 4233 64843 4267
rect 64785 4227 64843 4233
rect 356146 4224 356152 4276
rect 356204 4264 356210 4276
rect 357342 4264 357348 4276
rect 356204 4236 357348 4264
rect 356204 4224 356210 4236
rect 357342 4224 357348 4236
rect 357400 4224 357406 4276
rect 59909 4199 59967 4205
rect 59909 4165 59921 4199
rect 59955 4196 59967 4199
rect 61378 4196 61384 4208
rect 59955 4168 61384 4196
rect 59955 4165 59967 4168
rect 59909 4159 59967 4165
rect 61378 4156 61384 4168
rect 61436 4156 61442 4208
rect 96617 4199 96675 4205
rect 96617 4196 96629 4199
rect 74460 4168 75316 4196
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 21910 4128 21916 4140
rect 20772 4100 21916 4128
rect 20772 4088 20778 4100
rect 21910 4088 21916 4100
rect 21968 4088 21974 4140
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4128 22063 4131
rect 71130 4128 71136 4140
rect 22051 4100 71136 4128
rect 22051 4097 22063 4100
rect 22005 4091 22063 4097
rect 71130 4088 71136 4100
rect 71188 4088 71194 4140
rect 74258 4088 74264 4140
rect 74316 4128 74322 4140
rect 74460 4128 74488 4168
rect 75288 4137 75316 4168
rect 93228 4168 93900 4196
rect 74316 4100 74488 4128
rect 75273 4131 75331 4137
rect 74316 4088 74322 4100
rect 75273 4097 75285 4131
rect 75319 4097 75331 4131
rect 75273 4091 75331 4097
rect 84105 4131 84163 4137
rect 84105 4097 84117 4131
rect 84151 4128 84163 4131
rect 93228 4128 93256 4168
rect 84151 4100 93256 4128
rect 84151 4097 84163 4100
rect 84105 4091 84163 4097
rect 93302 4088 93308 4140
rect 93360 4128 93366 4140
rect 93762 4128 93768 4140
rect 93360 4100 93768 4128
rect 93360 4088 93366 4100
rect 93762 4088 93768 4100
rect 93820 4088 93826 4140
rect 93872 4128 93900 4168
rect 95620 4168 96629 4196
rect 95620 4128 95648 4168
rect 96617 4165 96629 4168
rect 96663 4165 96675 4199
rect 96617 4159 96675 4165
rect 145576 4168 146340 4196
rect 93872 4100 95648 4128
rect 95694 4088 95700 4140
rect 95752 4128 95758 4140
rect 96522 4128 96528 4140
rect 95752 4100 96528 4128
rect 95752 4088 95758 4100
rect 96522 4088 96528 4100
rect 96580 4088 96586 4140
rect 96709 4131 96767 4137
rect 96709 4097 96721 4131
rect 96755 4128 96767 4131
rect 106277 4131 106335 4137
rect 106277 4128 106289 4131
rect 96755 4100 106289 4128
rect 96755 4097 96767 4100
rect 96709 4091 96767 4097
rect 106277 4097 106289 4100
rect 106323 4097 106335 4131
rect 106277 4091 106335 4097
rect 112346 4088 112352 4140
rect 112404 4128 112410 4140
rect 113082 4128 113088 4140
rect 112404 4100 113088 4128
rect 112404 4088 112410 4100
rect 113082 4088 113088 4100
rect 113140 4088 113146 4140
rect 113542 4088 113548 4140
rect 113600 4128 113606 4140
rect 114462 4128 114468 4140
rect 113600 4100 114468 4128
rect 113600 4088 113606 4100
rect 114462 4088 114468 4100
rect 114520 4088 114526 4140
rect 119430 4088 119436 4140
rect 119488 4128 119494 4140
rect 119982 4128 119988 4140
rect 119488 4100 119988 4128
rect 119488 4088 119494 4100
rect 119982 4088 119988 4100
rect 120040 4088 120046 4140
rect 120626 4088 120632 4140
rect 120684 4128 120690 4140
rect 121362 4128 121368 4140
rect 120684 4100 121368 4128
rect 120684 4088 120690 4100
rect 121362 4088 121368 4100
rect 121420 4088 121426 4140
rect 123018 4088 123024 4140
rect 123076 4128 123082 4140
rect 124122 4128 124128 4140
rect 123076 4100 124128 4128
rect 123076 4088 123082 4100
rect 124122 4088 124128 4100
rect 124180 4088 124186 4140
rect 136082 4088 136088 4140
rect 136140 4128 136146 4140
rect 136542 4128 136548 4140
rect 136140 4100 136548 4128
rect 136140 4088 136146 4100
rect 136542 4088 136548 4100
rect 136600 4088 136606 4140
rect 138474 4088 138480 4140
rect 138532 4128 138538 4140
rect 139302 4128 139308 4140
rect 138532 4100 139308 4128
rect 138532 4088 138538 4100
rect 139302 4088 139308 4100
rect 139360 4088 139366 4140
rect 140866 4088 140872 4140
rect 140924 4128 140930 4140
rect 145576 4128 145604 4168
rect 140924 4100 145604 4128
rect 140924 4088 140930 4100
rect 145650 4088 145656 4140
rect 145708 4128 145714 4140
rect 146202 4128 146208 4140
rect 145708 4100 146208 4128
rect 145708 4088 145714 4100
rect 146202 4088 146208 4100
rect 146260 4088 146266 4140
rect 146312 4128 146340 4168
rect 453942 4156 453948 4208
rect 454000 4196 454006 4208
rect 456245 4199 456303 4205
rect 456245 4196 456257 4199
rect 454000 4168 456257 4196
rect 454000 4156 454006 4168
rect 456245 4165 456257 4168
rect 456291 4165 456303 4199
rect 456245 4159 456303 4165
rect 175366 4128 175372 4140
rect 146312 4100 175372 4128
rect 175366 4088 175372 4100
rect 175424 4088 175430 4140
rect 193214 4088 193220 4140
rect 193272 4128 193278 4140
rect 194502 4128 194508 4140
rect 193272 4100 194508 4128
rect 193272 4088 193278 4100
rect 194502 4088 194508 4100
rect 194560 4088 194566 4140
rect 196802 4088 196808 4140
rect 196860 4128 196866 4140
rect 197262 4128 197268 4140
rect 196860 4100 197268 4128
rect 196860 4088 196866 4100
rect 197262 4088 197268 4100
rect 197320 4088 197326 4140
rect 199194 4088 199200 4140
rect 199252 4128 199258 4140
rect 200022 4128 200028 4140
rect 199252 4100 200028 4128
rect 199252 4088 199258 4100
rect 200022 4088 200028 4100
rect 200080 4088 200086 4140
rect 201494 4088 201500 4140
rect 201552 4128 201558 4140
rect 202690 4128 202696 4140
rect 201552 4100 202696 4128
rect 201552 4088 201558 4100
rect 202690 4088 202696 4100
rect 202748 4088 202754 4140
rect 205082 4088 205088 4140
rect 205140 4128 205146 4140
rect 205542 4128 205548 4140
rect 205140 4100 205548 4128
rect 205140 4088 205146 4100
rect 205542 4088 205548 4100
rect 205600 4088 205606 4140
rect 207474 4088 207480 4140
rect 207532 4128 207538 4140
rect 208302 4128 208308 4140
rect 207532 4100 208308 4128
rect 207532 4088 207538 4100
rect 208302 4088 208308 4100
rect 208360 4088 208366 4140
rect 208670 4088 208676 4140
rect 208728 4128 208734 4140
rect 209682 4128 209688 4140
rect 208728 4100 209688 4128
rect 208728 4088 208734 4100
rect 209682 4088 209688 4100
rect 209740 4088 209746 4140
rect 214650 4088 214656 4140
rect 214708 4128 214714 4140
rect 215202 4128 215208 4140
rect 214708 4100 215208 4128
rect 214708 4088 214714 4100
rect 215202 4088 215208 4100
rect 215260 4088 215266 4140
rect 332410 4088 332416 4140
rect 332468 4128 332474 4140
rect 332686 4128 332692 4140
rect 332468 4100 332692 4128
rect 332468 4088 332474 4100
rect 332686 4088 332692 4100
rect 332744 4088 332750 4140
rect 335354 4088 335360 4140
rect 335412 4128 335418 4140
rect 335906 4128 335912 4140
rect 335412 4100 335912 4128
rect 335412 4088 335418 4100
rect 335906 4088 335912 4100
rect 335964 4088 335970 4140
rect 339494 4088 339500 4140
rect 339552 4128 339558 4140
rect 340690 4128 340696 4140
rect 339552 4100 340696 4128
rect 339552 4088 339558 4100
rect 340690 4088 340696 4100
rect 340748 4088 340754 4140
rect 344922 4088 344928 4140
rect 344980 4128 344986 4140
rect 345474 4128 345480 4140
rect 344980 4100 345480 4128
rect 344980 4088 344986 4100
rect 345474 4088 345480 4100
rect 345532 4088 345538 4140
rect 353202 4088 353208 4140
rect 353260 4128 353266 4140
rect 356146 4128 356152 4140
rect 353260 4100 356152 4128
rect 353260 4088 353266 4100
rect 356146 4088 356152 4100
rect 356204 4088 356210 4140
rect 357434 4088 357440 4140
rect 357492 4128 357498 4140
rect 360930 4128 360936 4140
rect 357492 4100 360936 4128
rect 357492 4088 357498 4100
rect 360930 4088 360936 4100
rect 360988 4088 360994 4140
rect 362218 4088 362224 4140
rect 362276 4128 362282 4140
rect 365714 4128 365720 4140
rect 362276 4100 365720 4128
rect 362276 4088 362282 4100
rect 365714 4088 365720 4100
rect 365772 4088 365778 4140
rect 379422 4088 379428 4140
rect 379480 4128 379486 4140
rect 387058 4128 387064 4140
rect 379480 4100 387064 4128
rect 379480 4088 379486 4100
rect 387058 4088 387064 4100
rect 387116 4088 387122 4140
rect 397362 4088 397368 4140
rect 397420 4128 397426 4140
rect 409598 4128 409604 4140
rect 397420 4100 409604 4128
rect 397420 4088 397426 4100
rect 409598 4088 409604 4100
rect 409656 4088 409662 4140
rect 409690 4088 409696 4140
rect 409748 4128 409754 4140
rect 423950 4128 423956 4140
rect 409748 4100 423956 4128
rect 409748 4088 409754 4100
rect 423950 4088 423956 4100
rect 424008 4088 424014 4140
rect 430390 4088 430396 4140
rect 430448 4128 430454 4140
rect 431221 4131 431279 4137
rect 431221 4128 431233 4131
rect 430448 4100 431233 4128
rect 430448 4088 430454 4100
rect 431221 4097 431233 4100
rect 431267 4097 431279 4131
rect 431221 4091 431279 4097
rect 431862 4088 431868 4140
rect 431920 4128 431926 4140
rect 451274 4128 451280 4140
rect 431920 4100 451280 4128
rect 431920 4088 431926 4100
rect 451274 4088 451280 4100
rect 451332 4088 451338 4140
rect 452562 4088 452568 4140
rect 452620 4128 452626 4140
rect 476298 4128 476304 4140
rect 452620 4100 476304 4128
rect 452620 4088 452626 4100
rect 476298 4088 476304 4100
rect 476356 4088 476362 4140
rect 484302 4088 484308 4140
rect 484360 4128 484366 4140
rect 514386 4128 514392 4140
rect 484360 4100 514392 4128
rect 484360 4088 484366 4100
rect 514386 4088 514392 4100
rect 514444 4088 514450 4140
rect 514662 4088 514668 4140
rect 514720 4128 514726 4140
rect 552382 4128 552388 4140
rect 514720 4100 552388 4128
rect 514720 4088 514726 4100
rect 552382 4088 552388 4100
rect 552440 4088 552446 4140
rect 566458 4088 566464 4140
rect 566516 4128 566522 4140
rect 569034 4128 569040 4140
rect 566516 4100 569040 4128
rect 566516 4088 566522 4100
rect 569034 4088 569040 4100
rect 569092 4088 569098 4140
rect 35897 4063 35955 4069
rect 35897 4029 35909 4063
rect 35943 4060 35955 4063
rect 45465 4063 45523 4069
rect 45465 4060 45477 4063
rect 35943 4032 45477 4060
rect 35943 4029 35955 4032
rect 35897 4023 35955 4029
rect 45465 4029 45477 4032
rect 45511 4029 45523 4063
rect 45465 4023 45523 4029
rect 45649 4063 45707 4069
rect 45649 4029 45661 4063
rect 45695 4060 45707 4063
rect 88981 4063 89039 4069
rect 88981 4060 88993 4063
rect 45695 4032 88993 4060
rect 45695 4029 45707 4032
rect 45649 4023 45707 4029
rect 88981 4029 88993 4032
rect 89027 4029 89039 4063
rect 88981 4023 89039 4029
rect 111150 4020 111156 4072
rect 111208 4060 111214 4072
rect 142798 4060 142804 4072
rect 111208 4032 142804 4060
rect 111208 4020 111214 4032
rect 142798 4020 142804 4032
rect 142856 4020 142862 4072
rect 144454 4020 144460 4072
rect 144512 4060 144518 4072
rect 178034 4060 178040 4072
rect 144512 4032 178040 4060
rect 144512 4020 144518 4032
rect 178034 4020 178040 4032
rect 178092 4020 178098 4072
rect 190822 4020 190828 4072
rect 190880 4060 190886 4072
rect 200761 4063 200819 4069
rect 200761 4060 200773 4063
rect 190880 4032 200773 4060
rect 190880 4020 190886 4032
rect 200761 4029 200773 4032
rect 200807 4029 200819 4063
rect 200761 4023 200819 4029
rect 362770 4020 362776 4072
rect 362828 4060 362834 4072
rect 366910 4060 366916 4072
rect 362828 4032 366916 4060
rect 362828 4020 362834 4032
rect 366910 4020 366916 4032
rect 366968 4020 366974 4072
rect 384942 4020 384948 4072
rect 385000 4060 385006 4072
rect 394234 4060 394240 4072
rect 385000 4032 394240 4060
rect 385000 4020 385006 4032
rect 394234 4020 394240 4032
rect 394292 4020 394298 4072
rect 395890 4020 395896 4072
rect 395948 4060 395954 4072
rect 407298 4060 407304 4072
rect 395948 4032 407304 4060
rect 395948 4020 395954 4032
rect 407298 4020 407304 4032
rect 407356 4020 407362 4072
rect 412450 4020 412456 4072
rect 412508 4060 412514 4072
rect 427538 4060 427544 4072
rect 412508 4032 427544 4060
rect 412508 4020 412514 4032
rect 427538 4020 427544 4032
rect 427596 4020 427602 4072
rect 430482 4020 430488 4072
rect 430540 4060 430546 4072
rect 448974 4060 448980 4072
rect 430540 4032 448980 4060
rect 430540 4020 430546 4032
rect 448974 4020 448980 4032
rect 449032 4020 449038 4072
rect 449710 4020 449716 4072
rect 449768 4060 449774 4072
rect 472710 4060 472716 4072
rect 449768 4032 472716 4060
rect 449768 4020 449774 4032
rect 472710 4020 472716 4032
rect 472768 4020 472774 4072
rect 474550 4020 474556 4072
rect 474608 4060 474614 4072
rect 502426 4060 502432 4072
rect 474608 4032 502432 4060
rect 474608 4020 474614 4032
rect 502426 4020 502432 4032
rect 502484 4020 502490 4072
rect 503622 4020 503628 4072
rect 503680 4060 503686 4072
rect 503680 4032 531176 4060
rect 503680 4020 503686 4032
rect 8846 3952 8852 4004
rect 8904 3992 8910 4004
rect 61470 3992 61476 4004
rect 8904 3964 61476 3992
rect 8904 3952 8910 3964
rect 61470 3952 61476 3964
rect 61528 3952 61534 4004
rect 63586 3952 63592 4004
rect 63644 3992 63650 4004
rect 104158 3992 104164 4004
rect 63644 3964 104164 3992
rect 63644 3952 63650 3964
rect 104158 3952 104164 3964
rect 104216 3952 104222 4004
rect 121822 3952 121828 4004
rect 121880 3992 121886 4004
rect 156598 3992 156604 4004
rect 121880 3964 156604 3992
rect 121880 3952 121886 3964
rect 156598 3952 156604 3964
rect 156656 3952 156662 4004
rect 156693 3995 156751 4001
rect 156693 3961 156705 3995
rect 156739 3992 156751 3995
rect 160738 3992 160744 4004
rect 156739 3964 160744 3992
rect 156739 3961 156751 3964
rect 156693 3955 156751 3961
rect 160738 3952 160744 3964
rect 160796 3952 160802 4004
rect 161106 3952 161112 4004
rect 161164 3992 161170 4004
rect 161477 3995 161535 4001
rect 161477 3992 161489 3995
rect 161164 3964 161489 3992
rect 161164 3952 161170 3964
rect 161477 3961 161489 3964
rect 161523 3961 161535 3995
rect 161477 3955 161535 3961
rect 183738 3952 183744 4004
rect 183796 3992 183802 4004
rect 209866 3992 209872 4004
rect 183796 3964 209872 3992
rect 183796 3952 183802 3964
rect 209866 3952 209872 3964
rect 209924 3952 209930 4004
rect 313366 3952 313372 4004
rect 313424 3992 313430 4004
rect 316678 3992 316684 4004
rect 313424 3964 316684 3992
rect 313424 3952 313430 3964
rect 316678 3952 316684 3964
rect 316736 3952 316742 4004
rect 386322 3952 386328 4004
rect 386380 3992 386386 4004
rect 395430 3992 395436 4004
rect 386380 3964 395436 3992
rect 386380 3952 386386 3964
rect 395430 3952 395436 3964
rect 395488 3952 395494 4004
rect 400030 3952 400036 4004
rect 400088 3992 400094 4004
rect 412082 3992 412088 4004
rect 400088 3964 412088 3992
rect 400088 3952 400094 3964
rect 412082 3952 412088 3964
rect 412140 3952 412146 4004
rect 412542 3952 412548 4004
rect 412600 3992 412606 4004
rect 428734 3992 428740 4004
rect 412600 3964 428740 3992
rect 412600 3952 412606 3964
rect 428734 3952 428740 3964
rect 428792 3952 428798 4004
rect 429102 3952 429108 4004
rect 429160 3992 429166 4004
rect 447778 3992 447784 4004
rect 429160 3964 447784 3992
rect 429160 3952 429166 3964
rect 447778 3952 447784 3964
rect 447836 3952 447842 4004
rect 449802 3952 449808 4004
rect 449860 3992 449866 4004
rect 473906 3992 473912 4004
rect 449860 3964 473912 3992
rect 449860 3952 449866 3964
rect 473906 3952 473912 3964
rect 473964 3952 473970 4004
rect 477310 3952 477316 4004
rect 477368 3992 477374 4004
rect 507210 3992 507216 4004
rect 477368 3964 507216 3992
rect 477368 3952 477374 3964
rect 507210 3952 507216 3964
rect 507268 3952 507274 4004
rect 526438 3952 526444 4004
rect 526496 3992 526502 4004
rect 528646 3992 528652 4004
rect 526496 3964 528652 3992
rect 526496 3952 526502 3964
rect 528646 3952 528652 3964
rect 528704 3952 528710 4004
rect 531148 3992 531176 4032
rect 531222 4020 531228 4072
rect 531280 4060 531286 4072
rect 533433 4063 533491 4069
rect 533433 4060 533445 4063
rect 531280 4032 533445 4060
rect 531280 4020 531286 4032
rect 533433 4029 533445 4032
rect 533479 4029 533491 4063
rect 533433 4023 533491 4029
rect 538950 4020 538956 4072
rect 539008 4060 539014 4072
rect 577406 4060 577412 4072
rect 539008 4032 577412 4060
rect 539008 4020 539014 4032
rect 577406 4020 577412 4032
rect 577464 4020 577470 4072
rect 532881 3995 532939 4001
rect 532881 3992 532893 3995
rect 531148 3964 532893 3992
rect 532881 3961 532893 3964
rect 532927 3961 532939 3995
rect 532881 3955 532939 3961
rect 532973 3995 533031 4001
rect 532973 3961 532985 3995
rect 533019 3992 533031 3995
rect 563146 3992 563152 4004
rect 533019 3964 563152 3992
rect 533019 3961 533031 3964
rect 532973 3955 533031 3961
rect 563146 3952 563152 3964
rect 563204 3952 563210 4004
rect 16022 3884 16028 3936
rect 16080 3924 16086 3936
rect 26145 3927 26203 3933
rect 26145 3924 26157 3927
rect 16080 3896 26157 3924
rect 16080 3884 16086 3896
rect 26145 3893 26157 3896
rect 26191 3893 26203 3927
rect 26145 3887 26203 3893
rect 33870 3884 33876 3936
rect 33928 3924 33934 3936
rect 86954 3924 86960 3936
rect 33928 3896 86960 3924
rect 33928 3884 33934 3896
rect 86954 3884 86960 3896
rect 87012 3884 87018 3936
rect 92106 3884 92112 3936
rect 92164 3924 92170 3936
rect 112438 3924 112444 3936
rect 92164 3896 112444 3924
rect 92164 3884 92170 3896
rect 112438 3884 112444 3896
rect 112496 3884 112502 3936
rect 118234 3884 118240 3936
rect 118292 3924 118298 3936
rect 148689 3927 148747 3933
rect 148689 3924 148701 3927
rect 118292 3896 148701 3924
rect 118292 3884 118298 3896
rect 148689 3893 148701 3896
rect 148735 3893 148747 3927
rect 148689 3887 148747 3893
rect 149238 3884 149244 3936
rect 149296 3924 149302 3936
rect 150342 3924 150348 3936
rect 149296 3896 150348 3924
rect 149296 3884 149302 3896
rect 150342 3884 150348 3896
rect 150400 3884 150406 3936
rect 153930 3884 153936 3936
rect 153988 3924 153994 3936
rect 169018 3924 169024 3936
rect 153988 3896 169024 3924
rect 153988 3884 153994 3896
rect 169018 3884 169024 3896
rect 169076 3884 169082 3936
rect 169113 3927 169171 3933
rect 169113 3893 169125 3927
rect 169159 3924 169171 3927
rect 173158 3924 173164 3936
rect 169159 3896 173164 3924
rect 169159 3893 169171 3896
rect 169113 3887 169171 3893
rect 173158 3884 173164 3896
rect 173216 3884 173222 3936
rect 191101 3927 191159 3933
rect 191101 3893 191113 3927
rect 191147 3924 191159 3927
rect 198826 3924 198832 3936
rect 191147 3896 198832 3924
rect 191147 3893 191159 3896
rect 191101 3887 191159 3893
rect 198826 3884 198832 3896
rect 198884 3884 198890 3936
rect 200761 3927 200819 3933
rect 200761 3893 200773 3927
rect 200807 3924 200819 3927
rect 216674 3924 216680 3936
rect 200807 3896 216680 3924
rect 200807 3893 200819 3896
rect 200761 3887 200819 3893
rect 216674 3884 216680 3896
rect 216732 3884 216738 3936
rect 382182 3884 382188 3936
rect 382240 3924 382246 3936
rect 391750 3924 391756 3936
rect 382240 3896 391756 3924
rect 382240 3884 382246 3896
rect 391750 3884 391756 3896
rect 391808 3884 391814 3936
rect 393130 3884 393136 3936
rect 393188 3924 393194 3936
rect 404906 3924 404912 3936
rect 393188 3896 404912 3924
rect 393188 3884 393194 3896
rect 404906 3884 404912 3896
rect 404964 3884 404970 3936
rect 407022 3884 407028 3936
rect 407080 3924 407086 3936
rect 421558 3924 421564 3936
rect 407080 3896 421564 3924
rect 407080 3884 407086 3896
rect 421558 3884 421564 3896
rect 421616 3884 421622 3936
rect 423490 3884 423496 3936
rect 423548 3924 423554 3936
rect 440602 3924 440608 3936
rect 423548 3896 440608 3924
rect 423548 3884 423554 3896
rect 440602 3884 440608 3896
rect 440660 3884 440666 3936
rect 441522 3884 441528 3936
rect 441580 3924 441586 3936
rect 456061 3927 456119 3933
rect 441580 3896 456012 3924
rect 441580 3884 441586 3896
rect 19518 3816 19524 3868
rect 19576 3856 19582 3868
rect 22005 3859 22063 3865
rect 22005 3856 22017 3859
rect 19576 3828 22017 3856
rect 19576 3816 19582 3828
rect 22005 3825 22017 3828
rect 22051 3825 22063 3859
rect 22005 3819 22063 3825
rect 34974 3816 34980 3868
rect 35032 3856 35038 3868
rect 88334 3856 88340 3868
rect 35032 3828 88340 3856
rect 35032 3816 35038 3828
rect 88334 3816 88340 3828
rect 88392 3816 88398 3868
rect 88981 3859 89039 3865
rect 88981 3825 88993 3859
rect 89027 3856 89039 3859
rect 93854 3856 93860 3868
rect 89027 3828 93860 3856
rect 89027 3825 89039 3828
rect 88981 3819 89039 3825
rect 93854 3816 93860 3828
rect 93912 3816 93918 3868
rect 96890 3816 96896 3868
rect 96948 3856 96954 3868
rect 126238 3856 126244 3868
rect 96948 3828 126244 3856
rect 96948 3816 96954 3828
rect 126238 3816 126244 3828
rect 126296 3816 126302 3868
rect 130194 3816 130200 3868
rect 130252 3856 130258 3868
rect 165614 3856 165620 3868
rect 130252 3828 165620 3856
rect 130252 3816 130258 3828
rect 165614 3816 165620 3828
rect 165672 3816 165678 3868
rect 180150 3816 180156 3868
rect 180208 3856 180214 3868
rect 207014 3856 207020 3868
rect 180208 3828 207020 3856
rect 180208 3816 180214 3828
rect 207014 3816 207020 3828
rect 207072 3816 207078 3868
rect 360102 3816 360108 3868
rect 360160 3856 360166 3868
rect 364518 3856 364524 3868
rect 360160 3828 364524 3856
rect 360160 3816 360166 3828
rect 364518 3816 364524 3828
rect 364576 3816 364582 3868
rect 369762 3816 369768 3868
rect 369820 3856 369826 3868
rect 376386 3856 376392 3868
rect 369820 3828 376392 3856
rect 369820 3816 369826 3828
rect 376386 3816 376392 3828
rect 376444 3816 376450 3868
rect 383562 3816 383568 3868
rect 383620 3856 383626 3868
rect 393038 3856 393044 3868
rect 383620 3828 393044 3856
rect 383620 3816 383626 3828
rect 393038 3816 393044 3828
rect 393096 3816 393102 3868
rect 393222 3816 393228 3868
rect 393280 3856 393286 3868
rect 403710 3856 403716 3868
rect 393280 3828 403716 3856
rect 393280 3816 393286 3828
rect 403710 3816 403716 3828
rect 403768 3816 403774 3868
rect 404262 3816 404268 3868
rect 404320 3856 404326 3868
rect 417970 3856 417976 3868
rect 404320 3828 417976 3856
rect 404320 3816 404326 3828
rect 417970 3816 417976 3828
rect 418028 3816 418034 3868
rect 418062 3816 418068 3868
rect 418120 3856 418126 3868
rect 434530 3856 434536 3868
rect 418120 3828 434536 3856
rect 418120 3816 418126 3828
rect 434530 3816 434536 3828
rect 434588 3816 434594 3868
rect 434622 3816 434628 3868
rect 434680 3856 434686 3868
rect 454862 3856 454868 3868
rect 434680 3828 454868 3856
rect 434680 3816 434686 3828
rect 454862 3816 454868 3828
rect 454920 3816 454926 3868
rect 455984 3856 456012 3896
rect 456061 3893 456073 3927
rect 456107 3924 456119 3927
rect 462038 3924 462044 3936
rect 456107 3896 462044 3924
rect 456107 3893 456119 3896
rect 456061 3887 456119 3893
rect 462038 3884 462044 3896
rect 462096 3884 462102 3936
rect 464982 3884 464988 3936
rect 465040 3924 465046 3936
rect 491754 3924 491760 3936
rect 465040 3896 491760 3924
rect 465040 3884 465046 3896
rect 491754 3884 491760 3896
rect 491812 3884 491818 3936
rect 492582 3884 492588 3936
rect 492640 3924 492646 3936
rect 525058 3924 525064 3936
rect 492640 3896 525064 3924
rect 492640 3884 492646 3896
rect 525058 3884 525064 3896
rect 525116 3884 525122 3936
rect 528462 3884 528468 3936
rect 528520 3924 528526 3936
rect 567838 3924 567844 3936
rect 528520 3896 567844 3924
rect 528520 3884 528526 3896
rect 567838 3884 567844 3896
rect 567896 3884 567902 3936
rect 456153 3859 456211 3865
rect 456153 3856 456165 3859
rect 455984 3828 456165 3856
rect 456153 3825 456165 3828
rect 456199 3825 456211 3859
rect 456153 3819 456211 3825
rect 456702 3816 456708 3868
rect 456760 3856 456766 3868
rect 462133 3859 462191 3865
rect 462133 3856 462145 3859
rect 456760 3828 462145 3856
rect 456760 3816 456766 3828
rect 462133 3825 462145 3828
rect 462179 3825 462191 3859
rect 462133 3819 462191 3825
rect 462222 3816 462228 3868
rect 462280 3856 462286 3868
rect 488166 3856 488172 3868
rect 462280 3828 488172 3856
rect 462280 3816 462286 3828
rect 488166 3816 488172 3828
rect 488224 3816 488230 3868
rect 489822 3816 489828 3868
rect 489880 3856 489886 3868
rect 521470 3856 521476 3868
rect 489880 3828 521476 3856
rect 489880 3816 489886 3828
rect 521470 3816 521476 3828
rect 521528 3816 521534 3868
rect 524322 3816 524328 3868
rect 524380 3856 524386 3868
rect 532973 3859 533031 3865
rect 532973 3856 532985 3859
rect 524380 3828 532985 3856
rect 524380 3816 524386 3828
rect 532973 3825 532985 3828
rect 533019 3825 533031 3859
rect 532973 3819 533031 3825
rect 533341 3859 533399 3865
rect 533341 3825 533353 3859
rect 533387 3856 533399 3859
rect 564342 3856 564348 3868
rect 533387 3828 564348 3856
rect 533387 3825 533399 3828
rect 533341 3819 533399 3825
rect 564342 3816 564348 3828
rect 564400 3816 564406 3868
rect 25498 3748 25504 3800
rect 25556 3788 25562 3800
rect 80054 3788 80060 3800
rect 25556 3760 80060 3788
rect 25556 3748 25562 3760
rect 80054 3748 80060 3760
rect 80112 3748 80118 3800
rect 84105 3791 84163 3797
rect 84105 3788 84117 3791
rect 80164 3760 84117 3788
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 10100 3692 16528 3720
rect 10100 3680 10106 3692
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 12342 3584 12348 3596
rect 11296 3556 12348 3584
rect 11296 3544 11302 3556
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 16500 3584 16528 3692
rect 18322 3680 18328 3732
rect 18380 3720 18386 3732
rect 35897 3723 35955 3729
rect 35897 3720 35909 3723
rect 18380 3692 35909 3720
rect 18380 3680 18386 3692
rect 35897 3689 35909 3692
rect 35943 3689 35955 3723
rect 35897 3683 35955 3689
rect 45465 3723 45523 3729
rect 45465 3689 45477 3723
rect 45511 3720 45523 3723
rect 55217 3723 55275 3729
rect 55217 3720 55229 3723
rect 45511 3692 55229 3720
rect 45511 3689 45523 3692
rect 45465 3683 45523 3689
rect 55217 3689 55229 3692
rect 55263 3689 55275 3723
rect 55217 3683 55275 3689
rect 64785 3723 64843 3729
rect 64785 3689 64797 3723
rect 64831 3720 64843 3723
rect 64877 3723 64935 3729
rect 64877 3720 64889 3723
rect 64831 3692 64889 3720
rect 64831 3689 64843 3692
rect 64785 3683 64843 3689
rect 64877 3689 64889 3692
rect 64923 3689 64935 3723
rect 64877 3683 64935 3689
rect 69661 3723 69719 3729
rect 69661 3689 69673 3723
rect 69707 3720 69719 3723
rect 75178 3720 75184 3732
rect 69707 3692 75184 3720
rect 69707 3689 69719 3692
rect 69661 3683 69719 3689
rect 75178 3680 75184 3692
rect 75236 3680 75242 3732
rect 75273 3723 75331 3729
rect 75273 3689 75285 3723
rect 75319 3720 75331 3723
rect 80164 3720 80192 3760
rect 84105 3757 84117 3760
rect 84151 3757 84163 3791
rect 84105 3751 84163 3757
rect 89714 3748 89720 3800
rect 89772 3788 89778 3800
rect 122190 3788 122196 3800
rect 89772 3760 122196 3788
rect 89772 3748 89778 3760
rect 122190 3748 122196 3760
rect 122248 3748 122254 3800
rect 133782 3748 133788 3800
rect 133840 3788 133846 3800
rect 168374 3788 168380 3800
rect 133840 3760 168380 3788
rect 133840 3748 133846 3760
rect 168374 3748 168380 3760
rect 168432 3748 168438 3800
rect 172974 3748 172980 3800
rect 173032 3788 173038 3800
rect 201678 3788 201684 3800
rect 173032 3760 201684 3788
rect 173032 3748 173038 3760
rect 201678 3748 201684 3760
rect 201736 3748 201742 3800
rect 371142 3748 371148 3800
rect 371200 3788 371206 3800
rect 377582 3788 377588 3800
rect 371200 3760 377588 3788
rect 371200 3748 371206 3760
rect 377582 3748 377588 3760
rect 377640 3748 377646 3800
rect 380802 3748 380808 3800
rect 380860 3788 380866 3800
rect 389450 3788 389456 3800
rect 380860 3760 389456 3788
rect 380860 3748 380866 3760
rect 389450 3748 389456 3760
rect 389508 3748 389514 3800
rect 390462 3748 390468 3800
rect 390520 3788 390526 3800
rect 401318 3788 401324 3800
rect 390520 3760 401324 3788
rect 390520 3748 390526 3760
rect 401318 3748 401324 3760
rect 401376 3748 401382 3800
rect 401502 3748 401508 3800
rect 401560 3788 401566 3800
rect 414474 3788 414480 3800
rect 401560 3760 414480 3788
rect 401560 3748 401566 3760
rect 414474 3748 414480 3760
rect 414532 3748 414538 3800
rect 415302 3748 415308 3800
rect 415360 3788 415366 3800
rect 431126 3788 431132 3800
rect 415360 3760 431132 3788
rect 415360 3748 415366 3760
rect 431126 3748 431132 3760
rect 431184 3748 431190 3800
rect 431221 3791 431279 3797
rect 431221 3757 431233 3791
rect 431267 3788 431279 3791
rect 433153 3791 433211 3797
rect 433153 3788 433165 3791
rect 431267 3760 433165 3788
rect 431267 3757 431279 3760
rect 431221 3751 431279 3757
rect 433153 3757 433165 3760
rect 433199 3757 433211 3791
rect 433153 3751 433211 3757
rect 433242 3748 433248 3800
rect 433300 3788 433306 3800
rect 433300 3760 442304 3788
rect 433300 3748 433306 3760
rect 75319 3692 80192 3720
rect 75319 3689 75331 3692
rect 75273 3683 75331 3689
rect 82630 3680 82636 3732
rect 82688 3720 82694 3732
rect 115290 3720 115296 3732
rect 82688 3692 115296 3720
rect 82688 3680 82694 3692
rect 115290 3680 115296 3692
rect 115348 3680 115354 3732
rect 115934 3680 115940 3732
rect 115992 3720 115998 3732
rect 117222 3720 117228 3732
rect 115992 3692 117228 3720
rect 115992 3680 115998 3692
rect 117222 3680 117228 3692
rect 117280 3680 117286 3732
rect 124214 3680 124220 3732
rect 124272 3720 124278 3732
rect 125502 3720 125508 3732
rect 124272 3692 125508 3720
rect 124272 3680 124278 3692
rect 125502 3680 125508 3692
rect 125560 3680 125566 3732
rect 137278 3680 137284 3732
rect 137336 3720 137342 3732
rect 166261 3723 166319 3729
rect 166261 3720 166273 3723
rect 137336 3692 166273 3720
rect 137336 3680 137342 3692
rect 166261 3689 166273 3692
rect 166307 3689 166319 3723
rect 166261 3683 166319 3689
rect 176470 3680 176476 3732
rect 176528 3720 176534 3732
rect 204254 3720 204260 3732
rect 176528 3692 204260 3720
rect 176528 3680 176534 3692
rect 204254 3680 204260 3692
rect 204312 3680 204318 3732
rect 364242 3680 364248 3732
rect 364300 3720 364306 3732
rect 369210 3720 369216 3732
rect 364300 3692 369216 3720
rect 364300 3680 364306 3692
rect 369210 3680 369216 3692
rect 369268 3680 369274 3732
rect 389082 3680 389088 3732
rect 389140 3720 389146 3732
rect 399018 3720 399024 3732
rect 389140 3692 399024 3720
rect 389140 3680 389146 3692
rect 399018 3680 399024 3692
rect 399076 3680 399082 3732
rect 400122 3680 400128 3732
rect 400180 3720 400186 3732
rect 413278 3720 413284 3732
rect 400180 3692 413284 3720
rect 400180 3680 400186 3692
rect 413278 3680 413284 3692
rect 413336 3680 413342 3732
rect 413922 3680 413928 3732
rect 413980 3720 413986 3732
rect 429930 3720 429936 3732
rect 413980 3692 429936 3720
rect 413980 3680 413986 3692
rect 429930 3680 429936 3692
rect 429988 3680 429994 3732
rect 442276 3720 442304 3760
rect 445662 3748 445668 3800
rect 445720 3788 445726 3800
rect 453761 3791 453819 3797
rect 453761 3788 453773 3791
rect 445720 3760 453773 3788
rect 445720 3748 445726 3760
rect 453761 3757 453773 3760
rect 453807 3757 453819 3791
rect 453761 3751 453819 3757
rect 453850 3748 453856 3800
rect 453908 3788 453914 3800
rect 471793 3791 471851 3797
rect 471793 3788 471805 3791
rect 453908 3760 471805 3788
rect 453908 3748 453914 3760
rect 471793 3757 471805 3760
rect 471839 3757 471851 3791
rect 471793 3751 471851 3757
rect 471882 3748 471888 3800
rect 471940 3788 471946 3800
rect 476117 3791 476175 3797
rect 476117 3788 476129 3791
rect 471940 3760 476129 3788
rect 471940 3748 471946 3760
rect 476117 3757 476129 3760
rect 476163 3757 476175 3791
rect 476117 3751 476175 3757
rect 485682 3748 485688 3800
rect 485740 3788 485746 3800
rect 516778 3788 516784 3800
rect 485740 3760 516784 3788
rect 485740 3748 485746 3760
rect 516778 3748 516784 3760
rect 516836 3748 516842 3800
rect 521562 3748 521568 3800
rect 521620 3788 521626 3800
rect 560754 3788 560760 3800
rect 521620 3760 560760 3788
rect 521620 3748 521626 3760
rect 560754 3748 560760 3760
rect 560812 3748 560818 3800
rect 446677 3723 446735 3729
rect 446677 3720 446689 3723
rect 442276 3692 446689 3720
rect 446677 3689 446689 3692
rect 446723 3689 446735 3723
rect 446677 3683 446735 3689
rect 447042 3680 447048 3732
rect 447100 3720 447106 3732
rect 456245 3723 456303 3729
rect 447100 3692 456196 3720
rect 447100 3680 447106 3692
rect 26145 3655 26203 3661
rect 26145 3621 26157 3655
rect 26191 3652 26203 3655
rect 35989 3655 36047 3661
rect 35989 3652 36001 3655
rect 26191 3624 36001 3652
rect 26191 3621 26203 3624
rect 26145 3615 26203 3621
rect 35989 3621 36001 3624
rect 36035 3621 36047 3655
rect 35989 3615 36047 3621
rect 45373 3655 45431 3661
rect 45373 3621 45385 3655
rect 45419 3652 45431 3655
rect 55306 3652 55312 3664
rect 45419 3624 55312 3652
rect 45419 3621 45431 3624
rect 45373 3615 45431 3621
rect 55306 3612 55312 3624
rect 55364 3612 55370 3664
rect 64690 3612 64696 3664
rect 64748 3652 64754 3664
rect 68373 3655 68431 3661
rect 64748 3624 68324 3652
rect 64748 3612 64754 3624
rect 67818 3584 67824 3596
rect 16500 3556 67824 3584
rect 67818 3544 67824 3556
rect 67876 3544 67882 3596
rect 68296 3584 68324 3624
rect 68373 3621 68385 3655
rect 68419 3652 68431 3655
rect 108298 3652 108304 3664
rect 68419 3624 108304 3652
rect 68419 3621 68431 3624
rect 68373 3615 68431 3621
rect 108298 3612 108304 3624
rect 108356 3612 108362 3664
rect 109954 3612 109960 3664
rect 110012 3652 110018 3664
rect 149146 3652 149152 3664
rect 110012 3624 149152 3652
rect 110012 3612 110018 3624
rect 149146 3612 149152 3624
rect 149204 3612 149210 3664
rect 151538 3612 151544 3664
rect 151596 3652 151602 3664
rect 183554 3652 183560 3664
rect 151596 3624 183560 3652
rect 151596 3612 151602 3624
rect 183554 3612 183560 3624
rect 183612 3612 183618 3664
rect 187234 3612 187240 3664
rect 187292 3652 187298 3664
rect 212718 3652 212724 3664
rect 187292 3624 212724 3652
rect 187292 3612 187298 3624
rect 212718 3612 212724 3624
rect 212776 3612 212782 3664
rect 362862 3612 362868 3664
rect 362920 3652 362926 3664
rect 368014 3652 368020 3664
rect 362920 3624 368020 3652
rect 362920 3612 362926 3624
rect 368014 3612 368020 3624
rect 368072 3612 368078 3664
rect 387702 3612 387708 3664
rect 387760 3652 387766 3664
rect 397822 3652 397828 3664
rect 387760 3624 397828 3652
rect 387760 3612 387766 3624
rect 397822 3612 397828 3624
rect 397880 3612 397886 3664
rect 402790 3612 402796 3664
rect 402848 3652 402854 3664
rect 415670 3652 415676 3664
rect 402848 3624 415676 3652
rect 402848 3612 402854 3624
rect 415670 3612 415676 3624
rect 415728 3612 415734 3664
rect 416590 3612 416596 3664
rect 416648 3652 416654 3664
rect 433518 3652 433524 3664
rect 416648 3624 433524 3652
rect 416648 3612 416654 3624
rect 433518 3612 433524 3624
rect 433576 3612 433582 3664
rect 438762 3612 438768 3664
rect 438820 3652 438826 3664
rect 456058 3652 456064 3664
rect 438820 3624 456064 3652
rect 438820 3612 438826 3624
rect 456058 3612 456064 3624
rect 456116 3612 456122 3664
rect 71774 3584 71780 3596
rect 68296 3556 71780 3584
rect 71774 3544 71780 3556
rect 71832 3544 71838 3596
rect 71869 3587 71927 3593
rect 71869 3553 71881 3587
rect 71915 3584 71927 3587
rect 73798 3584 73804 3596
rect 71915 3556 73804 3584
rect 71915 3553 71927 3556
rect 71869 3547 71927 3553
rect 73798 3544 73804 3556
rect 73856 3544 73862 3596
rect 77294 3544 77300 3596
rect 77352 3584 77358 3596
rect 77938 3584 77944 3596
rect 77352 3556 77944 3584
rect 77352 3544 77358 3556
rect 77938 3544 77944 3556
rect 77996 3544 78002 3596
rect 79042 3544 79048 3596
rect 79100 3584 79106 3596
rect 79962 3584 79968 3596
rect 79100 3556 79968 3584
rect 79100 3544 79106 3556
rect 79962 3544 79968 3556
rect 80020 3544 80026 3596
rect 81434 3544 81440 3596
rect 81492 3584 81498 3596
rect 82722 3584 82728 3596
rect 81492 3556 82728 3584
rect 81492 3544 81498 3556
rect 82722 3544 82728 3556
rect 82780 3544 82786 3596
rect 82817 3587 82875 3593
rect 82817 3553 82829 3587
rect 82863 3584 82875 3587
rect 117958 3584 117964 3596
rect 82863 3556 117964 3584
rect 82863 3553 82875 3556
rect 82817 3547 82875 3553
rect 117958 3544 117964 3556
rect 118016 3544 118022 3596
rect 125410 3544 125416 3596
rect 125468 3584 125474 3596
rect 156693 3587 156751 3593
rect 156693 3584 156705 3587
rect 125468 3556 156705 3584
rect 125468 3544 125474 3556
rect 156693 3553 156705 3556
rect 156739 3553 156751 3587
rect 156693 3547 156751 3553
rect 158714 3544 158720 3596
rect 158772 3584 158778 3596
rect 159910 3584 159916 3596
rect 158772 3556 159916 3584
rect 158772 3544 158778 3556
rect 159910 3544 159916 3556
rect 159968 3544 159974 3596
rect 161477 3587 161535 3593
rect 161477 3553 161489 3587
rect 161523 3584 161535 3587
rect 169113 3587 169171 3593
rect 169113 3584 169125 3587
rect 161523 3556 169125 3584
rect 161523 3553 161535 3556
rect 161477 3547 161535 3553
rect 169113 3553 169125 3556
rect 169159 3553 169171 3587
rect 169113 3547 169171 3553
rect 169386 3544 169392 3596
rect 169444 3584 169450 3596
rect 191101 3587 191159 3593
rect 191101 3584 191113 3587
rect 169444 3556 191113 3584
rect 169444 3544 169450 3556
rect 191101 3553 191113 3556
rect 191147 3553 191159 3587
rect 196066 3584 196072 3596
rect 191101 3547 191159 3553
rect 191208 3556 196072 3584
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 59909 3519 59967 3525
rect 59909 3516 59921 3519
rect 4120 3488 59921 3516
rect 4120 3476 4126 3488
rect 59909 3485 59921 3488
rect 59955 3485 59967 3519
rect 59909 3479 59967 3485
rect 59998 3476 60004 3528
rect 60056 3516 60062 3528
rect 60642 3516 60648 3528
rect 60056 3488 60648 3516
rect 60056 3476 60062 3488
rect 60642 3476 60648 3488
rect 60700 3476 60706 3528
rect 61194 3476 61200 3528
rect 61252 3516 61258 3528
rect 68189 3519 68247 3525
rect 68189 3516 68201 3519
rect 61252 3488 68201 3516
rect 61252 3476 61258 3488
rect 68189 3485 68201 3488
rect 68235 3485 68247 3519
rect 68189 3479 68247 3485
rect 68278 3476 68284 3528
rect 68336 3516 68342 3528
rect 104161 3519 104219 3525
rect 104161 3516 104173 3519
rect 68336 3488 104173 3516
rect 68336 3476 68342 3488
rect 104161 3485 104173 3488
rect 104207 3485 104219 3519
rect 104161 3479 104219 3485
rect 126606 3476 126612 3528
rect 126664 3516 126670 3528
rect 162946 3516 162952 3528
rect 126664 3488 162952 3516
rect 126664 3476 126670 3488
rect 162946 3476 162952 3488
rect 163004 3476 163010 3528
rect 163498 3476 163504 3528
rect 163556 3516 163562 3528
rect 164142 3516 164148 3528
rect 163556 3488 164148 3516
rect 163556 3476 163562 3488
rect 164142 3476 164148 3488
rect 164200 3476 164206 3528
rect 164694 3476 164700 3528
rect 164752 3516 164758 3528
rect 165522 3516 165528 3528
rect 164752 3488 165528 3516
rect 164752 3476 164758 3488
rect 165522 3476 165528 3488
rect 165580 3476 165586 3528
rect 165890 3476 165896 3528
rect 165948 3516 165954 3528
rect 191208 3516 191236 3556
rect 196066 3544 196072 3556
rect 196124 3544 196130 3596
rect 218146 3544 218152 3596
rect 218204 3584 218210 3596
rect 219342 3584 219348 3596
rect 218204 3556 219348 3584
rect 218204 3544 218210 3556
rect 219342 3544 219348 3556
rect 219400 3544 219406 3596
rect 252646 3544 252652 3596
rect 252704 3584 252710 3596
rect 253842 3584 253848 3596
rect 252704 3556 253848 3584
rect 252704 3544 252710 3556
rect 253842 3544 253848 3556
rect 253900 3544 253906 3596
rect 270494 3544 270500 3596
rect 270552 3584 270558 3596
rect 271690 3584 271696 3596
rect 270552 3556 271696 3584
rect 270552 3544 270558 3556
rect 271690 3544 271696 3556
rect 271748 3544 271754 3596
rect 278866 3544 278872 3596
rect 278924 3584 278930 3596
rect 280062 3584 280068 3596
rect 278924 3556 280068 3584
rect 278924 3544 278930 3556
rect 280062 3544 280068 3556
rect 280120 3544 280126 3596
rect 287146 3544 287152 3596
rect 287204 3584 287210 3596
rect 288342 3584 288348 3596
rect 287204 3556 288348 3584
rect 287204 3544 287210 3556
rect 288342 3544 288348 3556
rect 288400 3544 288406 3596
rect 296714 3544 296720 3596
rect 296772 3584 296778 3596
rect 297910 3584 297916 3596
rect 296772 3556 297916 3584
rect 296772 3544 296778 3556
rect 297910 3544 297916 3556
rect 297968 3544 297974 3596
rect 304994 3544 305000 3596
rect 305052 3584 305058 3596
rect 306190 3584 306196 3596
rect 305052 3556 306196 3584
rect 305052 3544 305058 3556
rect 306190 3544 306196 3556
rect 306248 3544 306254 3596
rect 348970 3544 348976 3596
rect 349028 3584 349034 3596
rect 351362 3584 351368 3596
rect 349028 3556 351368 3584
rect 349028 3544 349034 3556
rect 351362 3544 351368 3556
rect 351420 3544 351426 3596
rect 351730 3544 351736 3596
rect 351788 3584 351794 3596
rect 354950 3584 354956 3596
rect 351788 3556 354956 3584
rect 351788 3544 351794 3556
rect 354950 3544 354956 3556
rect 355008 3544 355014 3596
rect 358722 3544 358728 3596
rect 358780 3584 358786 3596
rect 363322 3584 363328 3596
rect 358780 3556 363328 3584
rect 358780 3544 358786 3556
rect 363322 3544 363328 3556
rect 363380 3544 363386 3596
rect 373902 3544 373908 3596
rect 373960 3584 373966 3596
rect 381170 3584 381176 3596
rect 373960 3556 381176 3584
rect 373960 3544 373966 3556
rect 381170 3544 381176 3556
rect 381228 3544 381234 3596
rect 382090 3544 382096 3596
rect 382148 3584 382154 3596
rect 390646 3584 390652 3596
rect 382148 3556 390652 3584
rect 382148 3544 382154 3556
rect 390646 3544 390652 3556
rect 390704 3544 390710 3596
rect 395982 3544 395988 3596
rect 396040 3584 396046 3596
rect 408494 3584 408500 3596
rect 396040 3556 408500 3584
rect 396040 3544 396046 3556
rect 408494 3544 408500 3556
rect 408552 3544 408558 3596
rect 409782 3544 409788 3596
rect 409840 3584 409846 3596
rect 425146 3584 425152 3596
rect 409840 3556 425152 3584
rect 409840 3544 409846 3556
rect 425146 3544 425152 3556
rect 425204 3544 425210 3596
rect 426342 3544 426348 3596
rect 426400 3584 426406 3596
rect 445386 3584 445392 3596
rect 426400 3556 445392 3584
rect 426400 3544 426406 3556
rect 445386 3544 445392 3556
rect 445444 3544 445450 3596
rect 445481 3587 445539 3593
rect 445481 3553 445493 3587
rect 445527 3584 445539 3587
rect 450170 3584 450176 3596
rect 445527 3556 450176 3584
rect 445527 3553 445539 3556
rect 445481 3547 445539 3553
rect 450170 3544 450176 3556
rect 450228 3544 450234 3596
rect 451182 3544 451188 3596
rect 451240 3584 451246 3596
rect 455969 3587 456027 3593
rect 455969 3584 455981 3587
rect 451240 3556 455981 3584
rect 451240 3544 451246 3556
rect 455969 3553 455981 3556
rect 456015 3553 456027 3587
rect 456168 3584 456196 3692
rect 456245 3689 456257 3723
rect 456291 3720 456303 3723
rect 457349 3723 457407 3729
rect 457349 3720 457361 3723
rect 456291 3692 457361 3720
rect 456291 3689 456303 3692
rect 456245 3683 456303 3689
rect 457349 3689 457361 3692
rect 457395 3689 457407 3723
rect 457349 3683 457407 3689
rect 459462 3680 459468 3732
rect 459520 3720 459526 3732
rect 484578 3720 484584 3732
rect 459520 3692 484584 3720
rect 459520 3680 459526 3692
rect 484578 3680 484584 3692
rect 484636 3680 484642 3732
rect 488442 3680 488448 3732
rect 488500 3720 488506 3732
rect 520274 3720 520280 3732
rect 488500 3692 520280 3720
rect 488500 3680 488506 3692
rect 520274 3680 520280 3692
rect 520332 3680 520338 3732
rect 524230 3680 524236 3732
rect 524288 3720 524294 3732
rect 533341 3723 533399 3729
rect 533341 3720 533353 3723
rect 524288 3692 533353 3720
rect 524288 3680 524294 3692
rect 533341 3689 533353 3692
rect 533387 3689 533399 3723
rect 533341 3683 533399 3689
rect 533433 3723 533491 3729
rect 533433 3689 533445 3723
rect 533479 3720 533491 3723
rect 571426 3720 571432 3732
rect 533479 3692 571432 3720
rect 533479 3689 533491 3692
rect 533433 3683 533491 3689
rect 571426 3680 571432 3692
rect 571484 3680 571490 3732
rect 456334 3612 456340 3664
rect 456392 3652 456398 3664
rect 459646 3652 459652 3664
rect 456392 3624 459652 3652
rect 456392 3612 456398 3624
rect 459646 3612 459652 3624
rect 459704 3612 459710 3664
rect 460842 3612 460848 3664
rect 460900 3652 460906 3664
rect 485774 3652 485780 3664
rect 460900 3624 485780 3652
rect 460900 3612 460906 3624
rect 485774 3612 485780 3624
rect 485832 3612 485838 3664
rect 491202 3612 491208 3664
rect 491260 3652 491266 3664
rect 523862 3652 523868 3664
rect 491260 3624 523868 3652
rect 491260 3612 491266 3624
rect 523862 3612 523868 3624
rect 523920 3612 523926 3664
rect 532602 3612 532608 3664
rect 532660 3652 532666 3664
rect 573818 3652 573824 3664
rect 532660 3624 573824 3652
rect 532660 3612 532666 3624
rect 573818 3612 573824 3624
rect 573876 3612 573882 3664
rect 470318 3584 470324 3596
rect 456168 3556 470324 3584
rect 455969 3547 456027 3553
rect 470318 3544 470324 3556
rect 470376 3544 470382 3596
rect 470502 3544 470508 3596
rect 470560 3584 470566 3596
rect 498930 3584 498936 3596
rect 470560 3556 498936 3584
rect 470560 3544 470566 3556
rect 498930 3544 498936 3556
rect 498988 3544 498994 3596
rect 500862 3544 500868 3596
rect 500920 3584 500926 3596
rect 500920 3556 529152 3584
rect 500920 3544 500926 3556
rect 165948 3488 191236 3516
rect 165948 3476 165954 3488
rect 215846 3476 215852 3528
rect 215904 3516 215910 3528
rect 216582 3516 216588 3528
rect 215904 3488 216588 3516
rect 215904 3476 215910 3488
rect 216582 3476 216588 3488
rect 216640 3476 216646 3528
rect 217042 3476 217048 3528
rect 217100 3516 217106 3528
rect 217962 3516 217968 3528
rect 217100 3488 217968 3516
rect 217100 3476 217106 3488
rect 217962 3476 217968 3488
rect 218020 3476 218026 3528
rect 222930 3476 222936 3528
rect 222988 3516 222994 3528
rect 223482 3516 223488 3528
rect 222988 3488 223488 3516
rect 222988 3476 222994 3488
rect 223482 3476 223488 3488
rect 223540 3476 223546 3528
rect 225322 3476 225328 3528
rect 225380 3516 225386 3528
rect 226242 3516 226248 3528
rect 225380 3488 226248 3516
rect 225380 3476 225386 3488
rect 226242 3476 226248 3488
rect 226300 3476 226306 3528
rect 226518 3476 226524 3528
rect 226576 3516 226582 3528
rect 227622 3516 227628 3528
rect 226576 3488 227628 3516
rect 226576 3476 226582 3488
rect 227622 3476 227628 3488
rect 227680 3476 227686 3528
rect 231302 3476 231308 3528
rect 231360 3516 231366 3528
rect 231762 3516 231768 3528
rect 231360 3488 231768 3516
rect 231360 3476 231366 3488
rect 231762 3476 231768 3488
rect 231820 3476 231826 3528
rect 232498 3476 232504 3528
rect 232556 3516 232562 3528
rect 233142 3516 233148 3528
rect 232556 3488 233148 3516
rect 232556 3476 232562 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 233694 3476 233700 3528
rect 233752 3516 233758 3528
rect 234522 3516 234528 3528
rect 233752 3488 234528 3516
rect 233752 3476 233758 3488
rect 234522 3476 234528 3488
rect 234580 3476 234586 3528
rect 239582 3476 239588 3528
rect 239640 3516 239646 3528
rect 240042 3516 240048 3528
rect 239640 3488 240048 3516
rect 239640 3476 239646 3488
rect 240042 3476 240048 3488
rect 240100 3476 240106 3528
rect 240778 3476 240784 3528
rect 240836 3516 240842 3528
rect 241422 3516 241428 3528
rect 240836 3488 241428 3516
rect 240836 3476 240842 3488
rect 241422 3476 241428 3488
rect 241480 3476 241486 3528
rect 243170 3476 243176 3528
rect 243228 3516 243234 3528
rect 244182 3516 244188 3528
rect 243228 3488 244188 3516
rect 243228 3476 243234 3488
rect 244182 3476 244188 3488
rect 244240 3476 244246 3528
rect 244366 3476 244372 3528
rect 244424 3516 244430 3528
rect 245470 3516 245476 3528
rect 244424 3488 245476 3516
rect 244424 3476 244430 3488
rect 245470 3476 245476 3488
rect 245528 3476 245534 3528
rect 249150 3476 249156 3528
rect 249208 3516 249214 3528
rect 249702 3516 249708 3528
rect 249208 3488 249708 3516
rect 249208 3476 249214 3488
rect 249702 3476 249708 3488
rect 249760 3476 249766 3528
rect 250346 3476 250352 3528
rect 250404 3516 250410 3528
rect 251082 3516 251088 3528
rect 250404 3488 251088 3516
rect 250404 3476 250410 3488
rect 251082 3476 251088 3488
rect 251140 3476 251146 3528
rect 251450 3476 251456 3528
rect 251508 3516 251514 3528
rect 252462 3516 252468 3528
rect 251508 3488 252468 3516
rect 251508 3476 251514 3488
rect 252462 3476 252468 3488
rect 252520 3476 252526 3528
rect 257430 3476 257436 3528
rect 257488 3516 257494 3528
rect 257982 3516 257988 3528
rect 257488 3488 257988 3516
rect 257488 3476 257494 3488
rect 257982 3476 257988 3488
rect 258040 3476 258046 3528
rect 259822 3476 259828 3528
rect 259880 3516 259886 3528
rect 260742 3516 260748 3528
rect 259880 3488 260748 3516
rect 259880 3476 259886 3488
rect 260742 3476 260748 3488
rect 260800 3476 260806 3528
rect 262214 3476 262220 3528
rect 262272 3516 262278 3528
rect 263502 3516 263508 3528
rect 262272 3488 263508 3516
rect 262272 3476 262278 3488
rect 263502 3476 263508 3488
rect 263560 3476 263566 3528
rect 265802 3476 265808 3528
rect 265860 3516 265866 3528
rect 266262 3516 266268 3528
rect 265860 3488 266268 3516
rect 265860 3476 265866 3488
rect 266262 3476 266268 3488
rect 266320 3476 266326 3528
rect 269298 3476 269304 3528
rect 269356 3516 269362 3528
rect 270402 3516 270408 3528
rect 269356 3488 270408 3516
rect 269356 3476 269362 3488
rect 270402 3476 270408 3488
rect 270460 3476 270466 3528
rect 274082 3476 274088 3528
rect 274140 3516 274146 3528
rect 274542 3516 274548 3528
rect 274140 3488 274548 3516
rect 274140 3476 274146 3488
rect 274542 3476 274548 3488
rect 274600 3476 274606 3528
rect 275278 3476 275284 3528
rect 275336 3516 275342 3528
rect 275922 3516 275928 3528
rect 275336 3488 275928 3516
rect 275336 3476 275342 3488
rect 275922 3476 275928 3488
rect 275980 3476 275986 3528
rect 276474 3476 276480 3528
rect 276532 3516 276538 3528
rect 277302 3516 277308 3528
rect 276532 3488 277308 3516
rect 276532 3476 276538 3488
rect 277302 3476 277308 3488
rect 277360 3476 277366 3528
rect 277670 3476 277676 3528
rect 277728 3516 277734 3528
rect 278682 3516 278688 3528
rect 277728 3488 278688 3516
rect 277728 3476 277734 3488
rect 278682 3476 278688 3488
rect 278740 3476 278746 3528
rect 283650 3476 283656 3528
rect 283708 3516 283714 3528
rect 284202 3516 284208 3528
rect 283708 3488 284208 3516
rect 283708 3476 283714 3488
rect 284202 3476 284208 3488
rect 284260 3476 284266 3528
rect 284754 3476 284760 3528
rect 284812 3516 284818 3528
rect 285582 3516 285588 3528
rect 284812 3488 285588 3516
rect 284812 3476 284818 3488
rect 285582 3476 285588 3488
rect 285640 3476 285646 3528
rect 285950 3476 285956 3528
rect 286008 3516 286014 3528
rect 286962 3516 286968 3528
rect 286008 3488 286968 3516
rect 286008 3476 286014 3488
rect 286962 3476 286968 3488
rect 287020 3476 287026 3528
rect 291930 3476 291936 3528
rect 291988 3516 291994 3528
rect 292482 3516 292488 3528
rect 291988 3488 292488 3516
rect 291988 3476 291994 3488
rect 292482 3476 292488 3488
rect 292540 3476 292546 3528
rect 293126 3476 293132 3528
rect 293184 3516 293190 3528
rect 293862 3516 293868 3528
rect 293184 3488 293868 3516
rect 293184 3476 293190 3488
rect 293862 3476 293868 3488
rect 293920 3476 293926 3528
rect 294322 3476 294328 3528
rect 294380 3516 294386 3528
rect 295242 3516 295248 3528
rect 294380 3488 295248 3516
rect 294380 3476 294386 3488
rect 295242 3476 295248 3488
rect 295300 3476 295306 3528
rect 295518 3476 295524 3528
rect 295576 3516 295582 3528
rect 296622 3516 296628 3528
rect 295576 3488 296628 3516
rect 295576 3476 295582 3488
rect 296622 3476 296628 3488
rect 296680 3476 296686 3528
rect 301406 3476 301412 3528
rect 301464 3516 301470 3528
rect 302142 3516 302148 3528
rect 301464 3488 302148 3516
rect 301464 3476 301470 3488
rect 302142 3476 302148 3488
rect 302200 3476 302206 3528
rect 302602 3476 302608 3528
rect 302660 3516 302666 3528
rect 303522 3516 303528 3528
rect 302660 3488 303528 3516
rect 302660 3476 302666 3488
rect 303522 3476 303528 3488
rect 303580 3476 303586 3528
rect 303798 3476 303804 3528
rect 303856 3516 303862 3528
rect 304902 3516 304908 3528
rect 303856 3488 304908 3516
rect 303856 3476 303862 3488
rect 304902 3476 304908 3488
rect 304960 3476 304966 3528
rect 308582 3476 308588 3528
rect 308640 3516 308646 3528
rect 309042 3516 309048 3528
rect 308640 3488 309048 3516
rect 308640 3476 308646 3488
rect 309042 3476 309048 3488
rect 309100 3476 309106 3528
rect 309778 3476 309784 3528
rect 309836 3516 309842 3528
rect 310422 3516 310428 3528
rect 309836 3488 310428 3516
rect 309836 3476 309842 3488
rect 310422 3476 310428 3488
rect 310480 3476 310486 3528
rect 310974 3476 310980 3528
rect 311032 3516 311038 3528
rect 311802 3516 311808 3528
rect 311032 3488 311808 3516
rect 311032 3476 311038 3488
rect 311802 3476 311808 3488
rect 311860 3476 311866 3528
rect 312170 3476 312176 3528
rect 312228 3516 312234 3528
rect 313182 3516 313188 3528
rect 312228 3488 313188 3516
rect 312228 3476 312234 3488
rect 313182 3476 313188 3488
rect 313240 3476 313246 3528
rect 314562 3476 314568 3528
rect 314620 3516 314626 3528
rect 315298 3516 315304 3528
rect 314620 3488 315304 3516
rect 314620 3476 314626 3488
rect 315298 3476 315304 3488
rect 315356 3476 315362 3528
rect 318058 3476 318064 3528
rect 318116 3516 318122 3528
rect 319438 3516 319444 3528
rect 318116 3488 319444 3516
rect 318116 3476 318122 3488
rect 319438 3476 319444 3488
rect 319496 3476 319502 3528
rect 320450 3476 320456 3528
rect 320508 3516 320514 3528
rect 321462 3516 321468 3528
rect 320508 3488 321468 3516
rect 320508 3476 320514 3488
rect 321462 3476 321468 3488
rect 321520 3476 321526 3528
rect 321646 3476 321652 3528
rect 321704 3516 321710 3528
rect 322750 3516 322756 3528
rect 321704 3488 322756 3516
rect 321704 3476 321710 3488
rect 322750 3476 322756 3488
rect 322808 3476 322814 3528
rect 326430 3476 326436 3528
rect 326488 3516 326494 3528
rect 326982 3516 326988 3528
rect 326488 3488 326988 3516
rect 326488 3476 326494 3488
rect 326982 3476 326988 3488
rect 327040 3476 327046 3528
rect 327626 3476 327632 3528
rect 327684 3516 327690 3528
rect 328362 3516 328368 3528
rect 327684 3488 328368 3516
rect 327684 3476 327690 3488
rect 328362 3476 328368 3488
rect 328420 3476 328426 3528
rect 328822 3476 328828 3528
rect 328880 3516 328886 3528
rect 329926 3516 329932 3528
rect 328880 3488 329932 3516
rect 328880 3476 328886 3488
rect 329926 3476 329932 3488
rect 329984 3476 329990 3528
rect 340874 3476 340880 3528
rect 340932 3516 340938 3528
rect 341886 3516 341892 3528
rect 340932 3488 341892 3516
rect 340932 3476 340938 3488
rect 341886 3476 341892 3488
rect 341944 3476 341950 3528
rect 342162 3476 342168 3528
rect 342220 3516 342226 3528
rect 343082 3516 343088 3528
rect 342220 3488 343088 3516
rect 342220 3476 342226 3488
rect 343082 3476 343088 3488
rect 343140 3476 343146 3528
rect 349062 3476 349068 3528
rect 349120 3516 349126 3528
rect 350258 3516 350264 3528
rect 349120 3488 350264 3516
rect 349120 3476 349126 3488
rect 350258 3476 350264 3488
rect 350316 3476 350322 3528
rect 367002 3476 367008 3528
rect 367060 3516 367066 3528
rect 372798 3516 372804 3528
rect 367060 3488 372804 3516
rect 367060 3476 367066 3488
rect 372798 3476 372804 3488
rect 372856 3476 372862 3528
rect 376662 3476 376668 3528
rect 376720 3516 376726 3528
rect 384666 3516 384672 3528
rect 376720 3488 384672 3516
rect 376720 3476 376726 3488
rect 384666 3476 384672 3488
rect 384724 3476 384730 3528
rect 386230 3476 386236 3528
rect 386288 3516 386294 3528
rect 396626 3516 396632 3528
rect 386288 3488 396632 3516
rect 386288 3476 386294 3488
rect 396626 3476 396632 3488
rect 396684 3476 396690 3528
rect 402882 3476 402888 3528
rect 402940 3516 402946 3528
rect 416866 3516 416872 3528
rect 402940 3488 416872 3516
rect 402940 3476 402946 3488
rect 416866 3476 416872 3488
rect 416924 3476 416930 3528
rect 419350 3476 419356 3528
rect 419408 3516 419414 3528
rect 437014 3516 437020 3528
rect 419408 3488 437020 3516
rect 419408 3476 419414 3488
rect 437014 3476 437020 3488
rect 437072 3476 437078 3528
rect 440050 3476 440056 3528
rect 440108 3516 440114 3528
rect 456061 3519 456119 3525
rect 456061 3516 456073 3519
rect 440108 3488 456073 3516
rect 440108 3476 440114 3488
rect 456061 3485 456073 3488
rect 456107 3485 456119 3519
rect 456061 3479 456119 3485
rect 456153 3519 456211 3525
rect 456153 3485 456165 3519
rect 456199 3516 456211 3519
rect 463234 3516 463240 3528
rect 456199 3488 463240 3516
rect 456199 3485 456211 3488
rect 456153 3479 456211 3485
rect 463234 3476 463240 3488
rect 463292 3476 463298 3528
rect 463602 3476 463608 3528
rect 463660 3516 463666 3528
rect 465905 3519 465963 3525
rect 463660 3488 465764 3516
rect 463660 3476 463666 3488
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 65058 3448 65064 3460
rect 6512 3420 65064 3448
rect 6512 3408 6518 3420
rect 65058 3408 65064 3420
rect 65116 3408 65122 3460
rect 65153 3451 65211 3457
rect 65153 3417 65165 3451
rect 65199 3448 65211 3451
rect 71777 3451 71835 3457
rect 71777 3448 71789 3451
rect 65199 3420 71789 3448
rect 65199 3417 65211 3420
rect 65153 3411 65211 3417
rect 71777 3417 71789 3420
rect 71823 3417 71835 3451
rect 71777 3411 71835 3417
rect 71866 3408 71872 3460
rect 71924 3448 71930 3460
rect 115198 3448 115204 3460
rect 71924 3420 115204 3448
rect 71924 3408 71930 3420
rect 115198 3408 115204 3420
rect 115256 3408 115262 3460
rect 117130 3408 117136 3460
rect 117188 3448 117194 3460
rect 148689 3451 148747 3457
rect 117188 3420 148640 3448
rect 117188 3408 117194 3420
rect 29086 3340 29092 3392
rect 29144 3380 29150 3392
rect 30190 3380 30196 3392
rect 29144 3352 30196 3380
rect 29144 3340 29150 3352
rect 30190 3340 30196 3352
rect 30248 3340 30254 3392
rect 77754 3380 77760 3392
rect 30392 3352 77760 3380
rect 26694 3204 26700 3256
rect 26752 3244 26758 3256
rect 30392 3244 30420 3352
rect 77754 3340 77760 3352
rect 77812 3340 77818 3392
rect 77846 3340 77852 3392
rect 77904 3380 77910 3392
rect 82817 3383 82875 3389
rect 82817 3380 82829 3383
rect 77904 3352 82829 3380
rect 77904 3340 77910 3352
rect 82817 3349 82829 3352
rect 82863 3349 82875 3383
rect 82817 3343 82875 3349
rect 84930 3340 84936 3392
rect 84988 3380 84994 3392
rect 85482 3380 85488 3392
rect 84988 3352 85488 3380
rect 84988 3340 84994 3352
rect 85482 3340 85488 3352
rect 85540 3340 85546 3392
rect 86126 3340 86132 3392
rect 86184 3380 86190 3392
rect 86862 3380 86868 3392
rect 86184 3352 86868 3380
rect 86184 3340 86190 3352
rect 86862 3340 86868 3352
rect 86920 3340 86926 3392
rect 88518 3340 88524 3392
rect 88576 3380 88582 3392
rect 89622 3380 89628 3392
rect 88576 3352 89628 3380
rect 88576 3340 88582 3352
rect 89622 3340 89628 3352
rect 89680 3340 89686 3392
rect 104161 3383 104219 3389
rect 104161 3349 104173 3383
rect 104207 3380 104219 3383
rect 109678 3380 109684 3392
rect 104207 3352 109684 3380
rect 104207 3349 104219 3352
rect 104161 3343 104219 3349
rect 109678 3340 109684 3352
rect 109736 3340 109742 3392
rect 114738 3340 114744 3392
rect 114796 3380 114802 3392
rect 145558 3380 145564 3392
rect 114796 3352 145564 3380
rect 114796 3340 114802 3352
rect 145558 3340 145564 3352
rect 145616 3340 145622 3392
rect 146846 3340 146852 3392
rect 146904 3380 146910 3392
rect 147582 3380 147588 3392
rect 146904 3352 147588 3380
rect 146904 3340 146910 3352
rect 147582 3340 147588 3352
rect 147640 3340 147646 3392
rect 36170 3272 36176 3324
rect 36228 3312 36234 3324
rect 37182 3312 37188 3324
rect 36228 3284 37188 3312
rect 36228 3272 36234 3284
rect 37182 3272 37188 3284
rect 37240 3272 37246 3324
rect 37366 3272 37372 3324
rect 37424 3312 37430 3324
rect 38470 3312 38476 3324
rect 37424 3284 38476 3312
rect 37424 3272 37430 3284
rect 38470 3272 38476 3284
rect 38528 3272 38534 3324
rect 43346 3272 43352 3324
rect 43404 3312 43410 3324
rect 44082 3312 44088 3324
rect 43404 3284 44088 3312
rect 43404 3272 43410 3284
rect 44082 3272 44088 3284
rect 44140 3272 44146 3324
rect 45649 3315 45707 3321
rect 45649 3312 45661 3315
rect 44192 3284 45661 3312
rect 26752 3216 30420 3244
rect 26752 3204 26758 3216
rect 42150 3204 42156 3256
rect 42208 3244 42214 3256
rect 44192 3244 44220 3284
rect 45649 3281 45661 3284
rect 45695 3281 45707 3315
rect 45649 3275 45707 3281
rect 45738 3272 45744 3324
rect 45796 3312 45802 3324
rect 46842 3312 46848 3324
rect 45796 3284 46848 3312
rect 45796 3272 45802 3284
rect 46842 3272 46848 3284
rect 46900 3272 46906 3324
rect 50522 3272 50528 3324
rect 50580 3312 50586 3324
rect 50982 3312 50988 3324
rect 50580 3284 50988 3312
rect 50580 3272 50586 3284
rect 50982 3272 50988 3284
rect 51040 3272 51046 3324
rect 52822 3272 52828 3324
rect 52880 3312 52886 3324
rect 53742 3312 53748 3324
rect 52880 3284 53748 3312
rect 52880 3272 52886 3284
rect 53742 3272 53748 3284
rect 53800 3272 53806 3324
rect 98638 3312 98644 3324
rect 53852 3284 98644 3312
rect 42208 3216 44220 3244
rect 42208 3204 42214 3216
rect 44542 3204 44548 3256
rect 44600 3244 44606 3256
rect 45462 3244 45468 3256
rect 44600 3216 45468 3244
rect 44600 3204 44606 3216
rect 45462 3204 45468 3216
rect 45520 3204 45526 3256
rect 49326 3204 49332 3256
rect 49384 3244 49390 3256
rect 53852 3244 53880 3284
rect 98638 3272 98644 3284
rect 98696 3272 98702 3324
rect 107654 3272 107660 3324
rect 107712 3312 107718 3324
rect 135898 3312 135904 3324
rect 107712 3284 135904 3312
rect 107712 3272 107718 3284
rect 135898 3272 135904 3284
rect 135956 3272 135962 3324
rect 148612 3312 148640 3420
rect 148689 3417 148701 3451
rect 148735 3448 148747 3451
rect 152458 3448 152464 3460
rect 148735 3420 152464 3448
rect 148735 3417 148747 3420
rect 148689 3411 148747 3417
rect 152458 3408 152464 3420
rect 152516 3408 152522 3460
rect 156322 3408 156328 3460
rect 156380 3448 156386 3460
rect 157242 3448 157248 3460
rect 156380 3420 157248 3448
rect 156380 3408 156386 3420
rect 157242 3408 157248 3420
rect 157300 3408 157306 3460
rect 157518 3408 157524 3460
rect 157576 3448 157582 3460
rect 158622 3448 158628 3460
rect 157576 3420 158628 3448
rect 157576 3408 157582 3420
rect 158622 3408 158628 3420
rect 158680 3408 158686 3460
rect 162302 3408 162308 3460
rect 162360 3448 162366 3460
rect 192294 3448 192300 3460
rect 162360 3420 192300 3448
rect 162360 3408 162366 3420
rect 192294 3408 192300 3420
rect 192352 3408 192358 3460
rect 194410 3408 194416 3460
rect 194468 3448 194474 3460
rect 219526 3448 219532 3460
rect 194468 3420 219532 3448
rect 194468 3408 194474 3420
rect 219526 3408 219532 3420
rect 219584 3408 219590 3460
rect 227714 3408 227720 3460
rect 227772 3448 227778 3460
rect 229002 3448 229008 3460
rect 227772 3420 229008 3448
rect 227772 3408 227778 3420
rect 229002 3408 229008 3420
rect 229060 3408 229066 3460
rect 241974 3408 241980 3460
rect 242032 3448 242038 3460
rect 242802 3448 242808 3460
rect 242032 3420 242808 3448
rect 242032 3408 242038 3420
rect 242802 3408 242808 3420
rect 242860 3408 242866 3460
rect 266998 3408 267004 3460
rect 267056 3448 267062 3460
rect 267642 3448 267648 3460
rect 267056 3420 267648 3448
rect 267056 3408 267062 3420
rect 267642 3408 267648 3420
rect 267700 3408 267706 3460
rect 319254 3408 319260 3460
rect 319312 3448 319318 3460
rect 320082 3448 320088 3460
rect 319312 3420 320088 3448
rect 319312 3408 319318 3420
rect 320082 3408 320088 3420
rect 320140 3408 320146 3460
rect 346210 3408 346216 3460
rect 346268 3448 346274 3460
rect 347866 3448 347872 3460
rect 346268 3420 347872 3448
rect 346268 3408 346274 3420
rect 347866 3408 347872 3420
rect 347924 3408 347930 3460
rect 355962 3408 355968 3460
rect 356020 3448 356026 3460
rect 359734 3448 359740 3460
rect 356020 3420 359740 3448
rect 356020 3408 356026 3420
rect 359734 3408 359740 3420
rect 359792 3408 359798 3460
rect 372522 3408 372528 3460
rect 372580 3448 372586 3460
rect 379974 3448 379980 3460
rect 372580 3420 379980 3448
rect 372580 3408 372586 3420
rect 379974 3408 379980 3420
rect 380032 3408 380038 3460
rect 380158 3408 380164 3460
rect 380216 3448 380222 3460
rect 388254 3448 388260 3460
rect 380216 3420 388260 3448
rect 380216 3408 380222 3420
rect 388254 3408 388260 3420
rect 388312 3408 388318 3460
rect 388990 3408 388996 3460
rect 389048 3448 389054 3460
rect 400214 3448 400220 3460
rect 389048 3420 400220 3448
rect 389048 3408 389054 3420
rect 400214 3408 400220 3420
rect 400272 3408 400278 3460
rect 408402 3408 408408 3460
rect 408460 3448 408466 3460
rect 422754 3448 422760 3460
rect 408460 3420 422760 3448
rect 408460 3408 408466 3420
rect 422754 3408 422760 3420
rect 422812 3408 422818 3460
rect 423582 3408 423588 3460
rect 423640 3448 423646 3460
rect 441798 3448 441804 3460
rect 423640 3420 441804 3448
rect 423640 3408 423646 3420
rect 441798 3408 441804 3420
rect 441856 3408 441862 3460
rect 442810 3408 442816 3460
rect 442868 3448 442874 3460
rect 465626 3448 465632 3460
rect 442868 3420 465632 3448
rect 442868 3408 442874 3420
rect 465626 3408 465632 3420
rect 465684 3408 465690 3460
rect 465736 3448 465764 3488
rect 465905 3485 465917 3519
rect 465951 3516 465963 3519
rect 471514 3516 471520 3528
rect 465951 3488 471520 3516
rect 465951 3485 465963 3488
rect 465905 3479 465963 3485
rect 471514 3476 471520 3488
rect 471572 3476 471578 3528
rect 492950 3516 492956 3528
rect 475396 3488 492956 3516
rect 465813 3451 465871 3457
rect 465813 3448 465825 3451
rect 465736 3420 465825 3448
rect 465813 3417 465825 3420
rect 465859 3417 465871 3451
rect 465813 3411 465871 3417
rect 466362 3408 466368 3460
rect 466420 3448 466426 3460
rect 475396 3448 475424 3488
rect 492950 3476 492956 3488
rect 493008 3476 493014 3528
rect 493962 3476 493968 3528
rect 494020 3516 494026 3528
rect 527450 3516 527456 3528
rect 494020 3488 527456 3516
rect 494020 3476 494026 3488
rect 527450 3476 527456 3488
rect 527508 3476 527514 3528
rect 529124 3516 529152 3556
rect 529198 3544 529204 3596
rect 529256 3584 529262 3596
rect 532234 3584 532240 3596
rect 529256 3556 532240 3584
rect 529256 3544 529262 3556
rect 532234 3544 532240 3556
rect 532292 3544 532298 3596
rect 532881 3587 532939 3593
rect 532881 3553 532893 3587
rect 532927 3584 532939 3587
rect 532927 3556 534672 3584
rect 532927 3553 532939 3556
rect 532881 3547 532939 3553
rect 534534 3516 534540 3528
rect 529124 3488 534540 3516
rect 534534 3476 534540 3488
rect 534592 3476 534598 3528
rect 534644 3516 534672 3556
rect 535362 3544 535368 3596
rect 535420 3584 535426 3596
rect 576210 3584 576216 3596
rect 535420 3556 576216 3584
rect 535420 3544 535426 3556
rect 576210 3544 576216 3556
rect 576268 3544 576274 3596
rect 534644 3488 535868 3516
rect 466420 3420 475424 3448
rect 476117 3451 476175 3457
rect 466420 3408 466426 3420
rect 476117 3417 476129 3451
rect 476163 3448 476175 3451
rect 500126 3448 500132 3460
rect 476163 3420 500132 3448
rect 476163 3417 476175 3420
rect 476117 3411 476175 3417
rect 500126 3408 500132 3420
rect 500184 3408 500190 3460
rect 500770 3408 500776 3460
rect 500828 3448 500834 3460
rect 535730 3448 535736 3460
rect 500828 3420 535736 3448
rect 500828 3408 500834 3420
rect 535730 3408 535736 3420
rect 535788 3408 535794 3460
rect 535840 3448 535868 3488
rect 536742 3476 536748 3528
rect 536800 3516 536806 3528
rect 578602 3516 578608 3528
rect 536800 3488 578608 3516
rect 536800 3476 536806 3488
rect 578602 3476 578608 3488
rect 578660 3476 578666 3528
rect 538030 3448 538036 3460
rect 535840 3420 538036 3448
rect 538030 3408 538036 3420
rect 538088 3408 538094 3460
rect 538122 3408 538128 3460
rect 538180 3448 538186 3460
rect 579798 3448 579804 3460
rect 538180 3420 579804 3448
rect 538180 3408 538186 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 150434 3340 150440 3392
rect 150492 3380 150498 3392
rect 164878 3380 164884 3392
rect 150492 3352 164884 3380
rect 150492 3340 150498 3352
rect 164878 3340 164884 3352
rect 164936 3340 164942 3392
rect 174170 3340 174176 3392
rect 174228 3380 174234 3392
rect 175182 3380 175188 3392
rect 174228 3352 175188 3380
rect 174228 3340 174234 3352
rect 175182 3340 175188 3352
rect 175240 3340 175246 3392
rect 175366 3340 175372 3392
rect 175424 3380 175430 3392
rect 176562 3380 176568 3392
rect 175424 3352 176568 3380
rect 175424 3340 175430 3352
rect 176562 3340 176568 3352
rect 176620 3340 176626 3392
rect 181346 3340 181352 3392
rect 181404 3380 181410 3392
rect 182082 3380 182088 3392
rect 181404 3352 182088 3380
rect 181404 3340 181410 3352
rect 182082 3340 182088 3352
rect 182140 3340 182146 3392
rect 182542 3340 182548 3392
rect 182600 3380 182606 3392
rect 183462 3380 183468 3392
rect 182600 3352 183468 3380
rect 182600 3340 182606 3352
rect 183462 3340 183468 3352
rect 183520 3340 183526 3392
rect 192018 3340 192024 3392
rect 192076 3380 192082 3392
rect 193122 3380 193128 3392
rect 192076 3352 193128 3380
rect 192076 3340 192082 3352
rect 193122 3340 193128 3352
rect 193180 3340 193186 3392
rect 200390 3340 200396 3392
rect 200448 3380 200454 3392
rect 201402 3380 201408 3392
rect 200448 3352 201408 3380
rect 200448 3340 200454 3352
rect 201402 3340 201408 3352
rect 201460 3340 201466 3392
rect 325234 3340 325240 3392
rect 325292 3380 325298 3392
rect 326338 3380 326344 3392
rect 325292 3352 326344 3380
rect 325292 3340 325298 3352
rect 326338 3340 326344 3352
rect 326396 3340 326402 3392
rect 375282 3340 375288 3392
rect 375340 3380 375346 3392
rect 382366 3380 382372 3392
rect 375340 3352 382372 3380
rect 375340 3340 375346 3352
rect 382366 3340 382372 3352
rect 382424 3340 382430 3392
rect 391842 3340 391848 3392
rect 391900 3380 391906 3392
rect 402514 3380 402520 3392
rect 391900 3352 402520 3380
rect 391900 3340 391906 3352
rect 402514 3340 402520 3352
rect 402572 3340 402578 3392
rect 405642 3340 405648 3392
rect 405700 3380 405706 3392
rect 419166 3380 419172 3392
rect 405700 3352 419172 3380
rect 405700 3340 405706 3352
rect 419166 3340 419172 3352
rect 419224 3340 419230 3392
rect 419442 3340 419448 3392
rect 419500 3380 419506 3392
rect 435818 3380 435824 3392
rect 419500 3352 435824 3380
rect 419500 3340 419506 3352
rect 435818 3340 435824 3352
rect 435876 3340 435882 3392
rect 437382 3340 437388 3392
rect 437440 3380 437446 3392
rect 457254 3380 457260 3392
rect 437440 3352 457260 3380
rect 437440 3340 437446 3352
rect 457254 3340 457260 3352
rect 457312 3340 457318 3392
rect 457349 3383 457407 3389
rect 457349 3349 457361 3383
rect 457395 3380 457407 3383
rect 460845 3383 460903 3389
rect 460845 3380 460857 3383
rect 457395 3352 460857 3380
rect 457395 3349 457407 3352
rect 457349 3343 457407 3349
rect 460845 3349 460857 3352
rect 460891 3349 460903 3383
rect 460845 3343 460903 3349
rect 462133 3383 462191 3389
rect 462133 3349 462145 3383
rect 462179 3380 462191 3383
rect 481082 3380 481088 3392
rect 462179 3352 481088 3380
rect 462179 3349 462191 3352
rect 462133 3343 462191 3349
rect 481082 3340 481088 3352
rect 481140 3340 481146 3392
rect 482922 3340 482928 3392
rect 482980 3380 482986 3392
rect 513190 3380 513196 3392
rect 482980 3352 513196 3380
rect 482980 3340 482986 3352
rect 513190 3340 513196 3352
rect 513248 3340 513254 3392
rect 517422 3340 517428 3392
rect 517480 3380 517486 3392
rect 549809 3383 549867 3389
rect 549809 3380 549821 3383
rect 517480 3352 549821 3380
rect 517480 3340 517486 3352
rect 549809 3349 549821 3352
rect 549855 3349 549867 3383
rect 549809 3343 549867 3349
rect 549898 3340 549904 3392
rect 549956 3380 549962 3392
rect 553578 3380 553584 3392
rect 549956 3352 553584 3380
rect 549956 3340 549962 3352
rect 553578 3340 553584 3352
rect 553636 3340 553642 3392
rect 153838 3312 153844 3324
rect 148612 3284 153844 3312
rect 153838 3272 153844 3284
rect 153896 3272 153902 3324
rect 166261 3315 166319 3321
rect 166261 3281 166273 3315
rect 166307 3312 166319 3315
rect 172698 3312 172704 3324
rect 166307 3284 172704 3312
rect 166307 3281 166319 3284
rect 166261 3275 166319 3281
rect 172698 3272 172704 3284
rect 172756 3272 172762 3324
rect 234798 3272 234804 3324
rect 234856 3312 234862 3324
rect 235902 3312 235908 3324
rect 234856 3284 235908 3312
rect 234856 3272 234862 3284
rect 235902 3272 235908 3284
rect 235960 3272 235966 3324
rect 300302 3272 300308 3324
rect 300360 3312 300366 3324
rect 304258 3312 304264 3324
rect 300360 3284 304264 3312
rect 300360 3272 300366 3284
rect 304258 3272 304264 3284
rect 304316 3272 304322 3324
rect 330018 3272 330024 3324
rect 330076 3312 330082 3324
rect 331122 3312 331128 3324
rect 330076 3284 331128 3312
rect 330076 3272 330082 3284
rect 331122 3272 331128 3284
rect 331180 3272 331186 3324
rect 334066 3272 334072 3324
rect 334124 3312 334130 3324
rect 334710 3312 334716 3324
rect 334124 3284 334716 3312
rect 334124 3272 334130 3284
rect 334710 3272 334716 3284
rect 334768 3272 334774 3324
rect 358630 3272 358636 3324
rect 358688 3312 358694 3324
rect 362126 3312 362132 3324
rect 358688 3284 362132 3312
rect 358688 3272 358694 3284
rect 362126 3272 362132 3284
rect 362184 3272 362190 3324
rect 365622 3272 365628 3324
rect 365680 3312 365686 3324
rect 371602 3312 371608 3324
rect 365680 3284 371608 3312
rect 365680 3272 365686 3284
rect 371602 3272 371608 3284
rect 371660 3272 371666 3324
rect 374638 3272 374644 3324
rect 374696 3312 374702 3324
rect 378778 3312 378784 3324
rect 374696 3284 378784 3312
rect 374696 3272 374702 3284
rect 378778 3272 378784 3284
rect 378836 3272 378842 3324
rect 398742 3272 398748 3324
rect 398800 3312 398806 3324
rect 410886 3312 410892 3324
rect 398800 3284 410892 3312
rect 398800 3272 398806 3284
rect 410886 3272 410892 3284
rect 410944 3272 410950 3324
rect 416682 3272 416688 3324
rect 416740 3312 416746 3324
rect 432322 3312 432328 3324
rect 416740 3284 432328 3312
rect 416740 3272 416746 3284
rect 432322 3272 432328 3284
rect 432380 3272 432386 3324
rect 433150 3272 433156 3324
rect 433208 3312 433214 3324
rect 452470 3312 452476 3324
rect 433208 3284 452476 3312
rect 433208 3272 433214 3284
rect 452470 3272 452476 3284
rect 452528 3272 452534 3324
rect 455322 3272 455328 3324
rect 455380 3312 455386 3324
rect 455877 3315 455935 3321
rect 455877 3312 455889 3315
rect 455380 3284 455889 3312
rect 455380 3272 455386 3284
rect 455877 3281 455889 3284
rect 455923 3281 455935 3315
rect 455877 3275 455935 3281
rect 455969 3315 456027 3321
rect 455969 3281 455981 3315
rect 456015 3312 456027 3315
rect 475102 3312 475108 3324
rect 456015 3284 475108 3312
rect 456015 3281 456027 3284
rect 455969 3275 456027 3281
rect 475102 3272 475108 3284
rect 475160 3272 475166 3324
rect 478690 3312 478696 3324
rect 475212 3284 478696 3312
rect 49384 3216 53880 3244
rect 49384 3204 49390 3216
rect 54018 3204 54024 3256
rect 54076 3244 54082 3256
rect 102778 3244 102784 3256
rect 54076 3216 102784 3244
rect 54076 3204 54082 3216
rect 102778 3204 102784 3216
rect 102836 3204 102842 3256
rect 106366 3204 106372 3256
rect 106424 3244 106430 3256
rect 107562 3244 107568 3256
rect 106424 3216 107568 3244
rect 106424 3204 106430 3216
rect 107562 3204 107568 3216
rect 107620 3204 107626 3256
rect 128906 3244 128912 3256
rect 107672 3216 128912 3244
rect 35989 3179 36047 3185
rect 35989 3145 36001 3179
rect 36035 3176 36047 3179
rect 45373 3179 45431 3185
rect 45373 3176 45385 3179
rect 36035 3148 45385 3176
rect 36035 3145 36047 3148
rect 35989 3139 36047 3145
rect 45373 3145 45385 3148
rect 45419 3145 45431 3179
rect 45373 3139 45431 3145
rect 56410 3136 56416 3188
rect 56468 3176 56474 3188
rect 102870 3176 102876 3188
rect 56468 3148 102876 3176
rect 56468 3136 56474 3148
rect 102870 3136 102876 3148
rect 102928 3136 102934 3188
rect 103974 3136 103980 3188
rect 104032 3176 104038 3188
rect 107672 3176 107700 3216
rect 128906 3204 128912 3216
rect 128964 3204 128970 3256
rect 235994 3204 236000 3256
rect 236052 3244 236058 3256
rect 237282 3244 237288 3256
rect 236052 3216 237288 3244
rect 236052 3204 236058 3216
rect 237282 3204 237288 3216
rect 237340 3204 237346 3256
rect 261018 3204 261024 3256
rect 261076 3244 261082 3256
rect 262122 3244 262128 3256
rect 261076 3216 262128 3244
rect 261076 3204 261082 3216
rect 262122 3204 262128 3216
rect 262180 3204 262186 3256
rect 376570 3204 376576 3256
rect 376628 3244 376634 3256
rect 383562 3244 383568 3256
rect 376628 3216 383568 3244
rect 376628 3204 376634 3216
rect 383562 3204 383568 3216
rect 383620 3204 383626 3256
rect 394602 3204 394608 3256
rect 394660 3244 394666 3256
rect 406102 3244 406108 3256
rect 394660 3216 406108 3244
rect 394660 3204 394666 3216
rect 406102 3204 406108 3216
rect 406160 3204 406166 3256
rect 406930 3204 406936 3256
rect 406988 3244 406994 3256
rect 420362 3244 420368 3256
rect 406988 3216 420368 3244
rect 406988 3204 406994 3216
rect 420362 3204 420368 3216
rect 420420 3204 420426 3256
rect 424962 3204 424968 3256
rect 425020 3244 425026 3256
rect 442994 3244 443000 3256
rect 425020 3216 443000 3244
rect 425020 3204 425026 3216
rect 442994 3204 443000 3216
rect 443052 3204 443058 3256
rect 444282 3204 444288 3256
rect 444340 3244 444346 3256
rect 466822 3244 466828 3256
rect 444340 3216 466828 3244
rect 444340 3204 444346 3216
rect 466822 3204 466828 3216
rect 466880 3204 466886 3256
rect 469309 3247 469367 3253
rect 469309 3244 469321 3247
rect 467024 3216 469321 3244
rect 104032 3148 107700 3176
rect 104032 3136 104038 3148
rect 167086 3136 167092 3188
rect 167144 3176 167150 3188
rect 168282 3176 168288 3188
rect 167144 3148 168288 3176
rect 167144 3136 167150 3148
rect 168282 3136 168288 3148
rect 168340 3136 168346 3188
rect 355870 3136 355876 3188
rect 355928 3176 355934 3188
rect 358538 3176 358544 3188
rect 355928 3148 358544 3176
rect 355928 3136 355934 3148
rect 358538 3136 358544 3148
rect 358596 3136 358602 3188
rect 378042 3136 378048 3188
rect 378100 3176 378106 3188
rect 385862 3176 385868 3188
rect 378100 3148 385868 3176
rect 378100 3136 378106 3148
rect 385862 3136 385868 3148
rect 385920 3136 385926 3188
rect 411162 3136 411168 3188
rect 411220 3176 411226 3188
rect 426342 3176 426348 3188
rect 411220 3148 426348 3176
rect 411220 3136 411226 3148
rect 426342 3136 426348 3148
rect 426400 3136 426406 3188
rect 427722 3136 427728 3188
rect 427780 3176 427786 3188
rect 446582 3176 446588 3188
rect 427780 3148 446588 3176
rect 427780 3136 427786 3148
rect 446582 3136 446588 3148
rect 446640 3136 446646 3188
rect 446677 3179 446735 3185
rect 446677 3145 446689 3179
rect 446723 3176 446735 3179
rect 452562 3176 452568 3188
rect 446723 3148 452568 3176
rect 446723 3145 446735 3148
rect 446677 3139 446735 3145
rect 452562 3136 452568 3148
rect 452620 3136 452626 3188
rect 465721 3179 465779 3185
rect 465721 3176 465733 3179
rect 452672 3148 465733 3176
rect 27890 3068 27896 3120
rect 27948 3108 27954 3120
rect 69661 3111 69719 3117
rect 69661 3108 69673 3111
rect 27948 3080 69673 3108
rect 27948 3068 27954 3080
rect 69661 3077 69673 3080
rect 69707 3077 69719 3111
rect 69661 3071 69719 3077
rect 70394 3068 70400 3120
rect 70452 3108 70458 3120
rect 71038 3108 71044 3120
rect 70452 3080 71044 3108
rect 70452 3068 70458 3080
rect 71038 3068 71044 3080
rect 71096 3068 71102 3120
rect 99282 3068 99288 3120
rect 99340 3108 99346 3120
rect 119338 3108 119344 3120
rect 99340 3080 119344 3108
rect 99340 3068 99346 3080
rect 119338 3068 119344 3080
rect 119396 3068 119402 3120
rect 189626 3068 189632 3120
rect 189684 3108 189690 3120
rect 190362 3108 190368 3120
rect 189684 3080 190368 3108
rect 189684 3068 189690 3080
rect 190362 3068 190368 3080
rect 190420 3068 190426 3120
rect 206278 3068 206284 3120
rect 206336 3108 206342 3120
rect 206922 3108 206928 3120
rect 206336 3080 206928 3108
rect 206336 3068 206342 3080
rect 206922 3068 206928 3080
rect 206980 3068 206986 3120
rect 258626 3068 258632 3120
rect 258684 3108 258690 3120
rect 259362 3108 259368 3120
rect 258684 3080 259368 3108
rect 258684 3068 258690 3080
rect 259362 3068 259368 3080
rect 259420 3068 259426 3120
rect 368382 3068 368388 3120
rect 368440 3108 368446 3120
rect 373994 3108 374000 3120
rect 368440 3080 374000 3108
rect 368440 3068 368446 3080
rect 373994 3068 374000 3080
rect 374052 3068 374058 3120
rect 426250 3068 426256 3120
rect 426308 3108 426314 3120
rect 444190 3108 444196 3120
rect 426308 3080 444196 3108
rect 426308 3068 426314 3080
rect 444190 3068 444196 3080
rect 444248 3068 444254 3120
rect 446950 3068 446956 3120
rect 447008 3108 447014 3120
rect 448330 3108 448336 3120
rect 447008 3080 448336 3108
rect 447008 3068 447014 3080
rect 448330 3068 448336 3080
rect 448388 3068 448394 3120
rect 448422 3068 448428 3120
rect 448480 3108 448486 3120
rect 452672 3108 452700 3148
rect 465721 3145 465733 3148
rect 465767 3145 465779 3179
rect 465721 3139 465779 3145
rect 465813 3179 465871 3185
rect 465813 3145 465825 3179
rect 465859 3176 465871 3179
rect 467024 3176 467052 3216
rect 469309 3213 469321 3216
rect 469355 3213 469367 3247
rect 469309 3207 469367 3213
rect 471793 3247 471851 3253
rect 471793 3213 471805 3247
rect 471839 3244 471851 3247
rect 475212 3244 475240 3284
rect 478690 3272 478696 3284
rect 478748 3272 478754 3324
rect 480162 3272 480168 3324
rect 480220 3312 480226 3324
rect 509602 3312 509608 3324
rect 480220 3284 509608 3312
rect 480220 3272 480226 3284
rect 509602 3272 509608 3284
rect 509660 3272 509666 3324
rect 518802 3272 518808 3324
rect 518860 3312 518866 3324
rect 557166 3312 557172 3324
rect 518860 3284 557172 3312
rect 518860 3272 518866 3284
rect 557166 3272 557172 3284
rect 557224 3272 557230 3324
rect 471839 3216 475240 3244
rect 471839 3213 471851 3216
rect 471793 3207 471851 3213
rect 477402 3204 477408 3256
rect 477460 3244 477466 3256
rect 506014 3244 506020 3256
rect 477460 3216 506020 3244
rect 477460 3204 477466 3216
rect 506014 3204 506020 3216
rect 506072 3204 506078 3256
rect 521378 3204 521384 3256
rect 521436 3244 521442 3256
rect 559558 3244 559564 3256
rect 521436 3216 559564 3244
rect 521436 3204 521442 3216
rect 559558 3204 559564 3216
rect 559616 3204 559622 3256
rect 465859 3148 467052 3176
rect 465859 3145 465871 3148
rect 465813 3139 465871 3145
rect 469122 3136 469128 3188
rect 469180 3136 469186 3188
rect 474642 3136 474648 3188
rect 474700 3176 474706 3188
rect 503622 3176 503628 3188
rect 474700 3148 503628 3176
rect 474700 3136 474706 3148
rect 503622 3136 503628 3148
rect 503680 3136 503686 3188
rect 506382 3136 506388 3188
rect 506440 3176 506446 3188
rect 541710 3176 541716 3188
rect 506440 3148 541716 3176
rect 506440 3136 506446 3148
rect 541710 3136 541716 3148
rect 541768 3136 541774 3188
rect 541894 3136 541900 3188
rect 541952 3176 541958 3188
rect 541952 3148 545436 3176
rect 541952 3136 541958 3148
rect 448480 3080 452700 3108
rect 453761 3111 453819 3117
rect 448480 3068 448486 3080
rect 453761 3077 453773 3111
rect 453807 3108 453819 3111
rect 467926 3108 467932 3120
rect 453807 3080 467932 3108
rect 453807 3077 453819 3080
rect 453761 3071 453819 3077
rect 467926 3068 467932 3080
rect 467984 3068 467990 3120
rect 469140 3108 469168 3136
rect 496538 3108 496544 3120
rect 469140 3080 496544 3108
rect 496538 3068 496544 3080
rect 496596 3068 496602 3120
rect 509142 3068 509148 3120
rect 509200 3108 509206 3120
rect 545298 3108 545304 3120
rect 509200 3080 545304 3108
rect 509200 3068 509206 3080
rect 545298 3068 545304 3080
rect 545356 3068 545362 3120
rect 545408 3108 545436 3148
rect 545758 3136 545764 3188
rect 545816 3176 545822 3188
rect 546494 3176 546500 3188
rect 545816 3148 546500 3176
rect 545816 3136 545822 3148
rect 546494 3136 546500 3148
rect 546552 3136 546558 3188
rect 547138 3136 547144 3188
rect 547196 3176 547202 3188
rect 550082 3176 550088 3188
rect 547196 3148 550088 3176
rect 547196 3136 547202 3148
rect 550082 3136 550088 3148
rect 550140 3136 550146 3188
rect 552661 3179 552719 3185
rect 552661 3145 552673 3179
rect 552707 3176 552719 3179
rect 582190 3176 582196 3188
rect 552707 3148 582196 3176
rect 552707 3145 552719 3148
rect 552661 3139 552719 3145
rect 582190 3136 582196 3148
rect 582248 3136 582254 3188
rect 545408 3080 556108 3108
rect 39758 3000 39764 3052
rect 39816 3040 39822 3052
rect 82078 3040 82084 3052
rect 39816 3012 82084 3040
rect 39816 3000 39822 3012
rect 82078 3000 82084 3012
rect 82136 3000 82142 3052
rect 170582 3000 170588 3052
rect 170640 3040 170646 3052
rect 171042 3040 171048 3052
rect 170640 3012 171048 3040
rect 170640 3000 170646 3012
rect 171042 3000 171048 3012
rect 171100 3000 171106 3052
rect 171778 3000 171784 3052
rect 171836 3040 171842 3052
rect 172422 3040 172428 3052
rect 171836 3012 172428 3040
rect 171836 3000 171842 3012
rect 172422 3000 172428 3012
rect 172480 3000 172486 3052
rect 188430 3000 188436 3052
rect 188488 3040 188494 3052
rect 188982 3040 188988 3052
rect 188488 3012 188988 3040
rect 188488 3000 188494 3012
rect 188982 3000 188988 3012
rect 189040 3000 189046 3052
rect 224126 3000 224132 3052
rect 224184 3040 224190 3052
rect 224862 3040 224868 3052
rect 224184 3012 224868 3040
rect 224184 3000 224190 3012
rect 224862 3000 224868 3012
rect 224920 3000 224926 3052
rect 268102 3000 268108 3052
rect 268160 3040 268166 3052
rect 269022 3040 269028 3052
rect 268160 3012 269028 3040
rect 268160 3000 268166 3012
rect 269022 3000 269028 3012
rect 269080 3000 269086 3052
rect 351822 3000 351828 3052
rect 351880 3040 351886 3052
rect 353754 3040 353760 3052
rect 351880 3012 353760 3040
rect 351880 3000 351886 3012
rect 353754 3000 353760 3012
rect 353812 3000 353818 3052
rect 422202 3000 422208 3052
rect 422260 3040 422266 3052
rect 439406 3040 439412 3052
rect 422260 3012 439412 3040
rect 422260 3000 422266 3012
rect 439406 3000 439412 3012
rect 439464 3000 439470 3052
rect 440142 3000 440148 3052
rect 440200 3040 440206 3052
rect 445573 3043 445631 3049
rect 445573 3040 445585 3043
rect 440200 3012 445585 3040
rect 440200 3000 440206 3012
rect 445573 3009 445585 3012
rect 445619 3009 445631 3043
rect 445573 3003 445631 3009
rect 451182 3000 451188 3052
rect 451240 3040 451246 3052
rect 469122 3040 469128 3052
rect 451240 3012 469128 3040
rect 451240 3000 451246 3012
rect 469122 3000 469128 3012
rect 469180 3000 469186 3052
rect 495342 3040 495348 3052
rect 469232 3012 495348 3040
rect 24302 2932 24308 2984
rect 24360 2972 24366 2984
rect 70394 2972 70400 2984
rect 24360 2944 70400 2972
rect 24360 2932 24366 2944
rect 70394 2932 70400 2944
rect 70452 2932 70458 2984
rect 70670 2932 70676 2984
rect 70728 2972 70734 2984
rect 105538 2972 105544 2984
rect 70728 2944 105544 2972
rect 70728 2932 70734 2944
rect 105538 2932 105544 2944
rect 105596 2932 105602 2984
rect 139670 2932 139676 2984
rect 139728 2972 139734 2984
rect 140682 2972 140688 2984
rect 139728 2944 140688 2972
rect 139728 2932 139734 2944
rect 140682 2932 140688 2944
rect 140740 2932 140746 2984
rect 197998 2932 198004 2984
rect 198056 2972 198062 2984
rect 198642 2972 198648 2984
rect 198056 2944 198648 2972
rect 198056 2932 198062 2944
rect 198642 2932 198648 2944
rect 198700 2932 198706 2984
rect 209866 2932 209872 2984
rect 209924 2972 209930 2984
rect 210970 2972 210976 2984
rect 209924 2944 210976 2972
rect 209924 2932 209930 2944
rect 210970 2932 210976 2944
rect 211028 2932 211034 2984
rect 420822 2932 420828 2984
rect 420880 2972 420886 2984
rect 438210 2972 438216 2984
rect 420880 2944 438216 2972
rect 420880 2932 420886 2944
rect 438210 2932 438216 2944
rect 438268 2932 438274 2984
rect 442902 2932 442908 2984
rect 442960 2972 442966 2984
rect 464430 2972 464436 2984
rect 442960 2944 464436 2972
rect 442960 2932 442966 2944
rect 464430 2932 464436 2944
rect 464488 2932 464494 2984
rect 467742 2932 467748 2984
rect 467800 2972 467806 2984
rect 469232 2972 469260 3012
rect 495342 3000 495348 3012
rect 495400 3000 495406 3052
rect 509878 3000 509884 3052
rect 509936 3040 509942 3052
rect 510893 3043 510951 3049
rect 510893 3040 510905 3043
rect 509936 3012 510905 3040
rect 509936 3000 509942 3012
rect 510893 3009 510905 3012
rect 510939 3009 510951 3043
rect 510893 3003 510951 3009
rect 511902 3000 511908 3052
rect 511960 3040 511966 3052
rect 548886 3040 548892 3052
rect 511960 3012 548892 3040
rect 511960 3000 511966 3012
rect 548886 3000 548892 3012
rect 548944 3000 548950 3052
rect 549809 3043 549867 3049
rect 549809 3009 549821 3043
rect 549855 3040 549867 3043
rect 555970 3040 555976 3052
rect 549855 3012 555976 3040
rect 549855 3009 549867 3012
rect 549809 3003 549867 3009
rect 555970 3000 555976 3012
rect 556028 3000 556034 3052
rect 467800 2944 469260 2972
rect 469309 2975 469367 2981
rect 467800 2932 467806 2944
rect 469309 2941 469321 2975
rect 469355 2972 469367 2975
rect 489362 2972 489368 2984
rect 469355 2944 489368 2972
rect 469355 2941 469367 2944
rect 469309 2935 469367 2941
rect 489362 2932 489368 2944
rect 489420 2932 489426 2984
rect 498102 2932 498108 2984
rect 498160 2972 498166 2984
rect 531038 2972 531044 2984
rect 498160 2944 531044 2972
rect 498160 2932 498166 2944
rect 531038 2932 531044 2944
rect 531096 2932 531102 2984
rect 533338 2932 533344 2984
rect 533396 2972 533402 2984
rect 533396 2944 543044 2972
rect 533396 2932 533402 2944
rect 32674 2864 32680 2916
rect 32732 2904 32738 2916
rect 77294 2904 77300 2916
rect 32732 2876 77300 2904
rect 32732 2864 32738 2876
rect 77294 2864 77300 2876
rect 77352 2864 77358 2916
rect 102778 2864 102784 2916
rect 102836 2904 102842 2916
rect 122098 2904 122104 2916
rect 102836 2876 122104 2904
rect 102836 2864 102842 2876
rect 122098 2864 122104 2876
rect 122156 2864 122162 2916
rect 369670 2864 369676 2916
rect 369728 2904 369734 2916
rect 375190 2904 375196 2916
rect 369728 2876 375196 2904
rect 369728 2864 369734 2876
rect 375190 2864 375196 2876
rect 375248 2864 375254 2916
rect 436002 2864 436008 2916
rect 436060 2904 436066 2916
rect 456058 2904 456064 2916
rect 436060 2876 456064 2904
rect 436060 2864 436066 2876
rect 456058 2864 456064 2876
rect 456116 2864 456122 2916
rect 456153 2907 456211 2913
rect 456153 2873 456165 2907
rect 456199 2904 456211 2907
rect 479886 2904 479892 2916
rect 456199 2876 479892 2904
rect 456199 2873 456211 2876
rect 456153 2867 456211 2873
rect 479886 2864 479892 2876
rect 479944 2864 479950 2916
rect 491938 2864 491944 2916
rect 491996 2904 492002 2916
rect 517882 2904 517888 2916
rect 491996 2876 517888 2904
rect 491996 2864 492002 2876
rect 517882 2864 517888 2876
rect 517940 2864 517946 2916
rect 537478 2864 537484 2916
rect 537536 2904 537542 2916
rect 543016 2904 543044 2944
rect 544378 2932 544384 2984
rect 544436 2972 544442 2984
rect 552661 2975 552719 2981
rect 552661 2972 552673 2975
rect 544436 2944 552673 2972
rect 544436 2932 544442 2944
rect 552661 2941 552673 2944
rect 552707 2941 552719 2975
rect 556080 2972 556108 3080
rect 575014 2972 575020 2984
rect 556080 2944 575020 2972
rect 552661 2935 552719 2941
rect 575014 2932 575020 2944
rect 575072 2932 575078 2984
rect 566734 2904 566740 2916
rect 537536 2876 542768 2904
rect 543016 2876 566740 2904
rect 537536 2864 537542 2876
rect 46934 2796 46940 2848
rect 46992 2836 46998 2848
rect 91738 2836 91744 2848
rect 46992 2808 91744 2836
rect 46992 2796 46998 2808
rect 91738 2796 91744 2808
rect 91796 2796 91802 2848
rect 143261 2839 143319 2845
rect 143261 2805 143273 2839
rect 143307 2836 143319 2839
rect 143442 2836 143448 2848
rect 143307 2808 143448 2836
rect 143307 2805 143319 2808
rect 143261 2799 143319 2805
rect 143442 2796 143448 2808
rect 143500 2796 143506 2848
rect 213457 2839 213515 2845
rect 213457 2805 213469 2839
rect 213503 2836 213515 2839
rect 213822 2836 213828 2848
rect 213503 2808 213828 2836
rect 213503 2805 213515 2808
rect 213457 2799 213515 2805
rect 213822 2796 213828 2808
rect 213880 2796 213886 2848
rect 333609 2839 333667 2845
rect 333609 2805 333621 2839
rect 333655 2836 333667 2839
rect 333882 2836 333888 2848
rect 333655 2808 333888 2836
rect 333655 2805 333667 2808
rect 333609 2799 333667 2805
rect 333882 2796 333888 2808
rect 333940 2796 333946 2848
rect 433153 2839 433211 2845
rect 433153 2805 433165 2839
rect 433199 2836 433211 2839
rect 445481 2839 445539 2845
rect 445481 2836 445493 2839
rect 433199 2808 445493 2836
rect 433199 2805 433211 2808
rect 433153 2799 433211 2805
rect 445481 2805 445493 2808
rect 445527 2805 445539 2839
rect 445481 2799 445539 2805
rect 445573 2839 445631 2845
rect 445573 2805 445585 2839
rect 445619 2836 445631 2839
rect 445619 2808 452608 2836
rect 445619 2805 445631 2808
rect 445573 2799 445631 2805
rect 452580 2768 452608 2808
rect 452654 2796 452660 2848
rect 452712 2836 452718 2848
rect 453666 2836 453672 2848
rect 452712 2808 453672 2836
rect 452712 2796 452718 2808
rect 453666 2796 453672 2808
rect 453724 2796 453730 2848
rect 460750 2836 460756 2848
rect 453776 2808 460756 2836
rect 453776 2768 453804 2808
rect 460750 2796 460756 2808
rect 460808 2796 460814 2848
rect 460845 2839 460903 2845
rect 460845 2805 460857 2839
rect 460891 2836 460903 2839
rect 477494 2836 477500 2848
rect 460891 2808 477500 2836
rect 460891 2805 460903 2808
rect 460845 2799 460903 2805
rect 477494 2796 477500 2808
rect 477552 2796 477558 2848
rect 489178 2796 489184 2848
rect 489236 2836 489242 2848
rect 510798 2836 510804 2848
rect 489236 2808 510804 2836
rect 489236 2796 489242 2808
rect 510798 2796 510804 2808
rect 510856 2796 510862 2848
rect 510893 2839 510951 2845
rect 510893 2805 510905 2839
rect 510939 2836 510951 2839
rect 539318 2836 539324 2848
rect 510939 2808 539324 2836
rect 510939 2805 510951 2808
rect 510893 2799 510951 2805
rect 539318 2796 539324 2808
rect 539376 2796 539382 2848
rect 542740 2836 542768 2876
rect 566734 2864 566740 2876
rect 566792 2864 566798 2916
rect 570230 2836 570236 2848
rect 542740 2808 570236 2836
rect 570230 2796 570236 2808
rect 570288 2796 570294 2848
rect 452580 2740 453804 2768
rect 5258 552 5264 604
rect 5316 592 5322 604
rect 5442 592 5448 604
rect 5316 564 5448 592
rect 5316 552 5322 564
rect 5442 552 5448 564
rect 5500 552 5506 604
rect 14826 552 14832 604
rect 14884 592 14890 604
rect 15102 592 15108 604
rect 14884 564 15108 592
rect 14884 552 14890 564
rect 15102 552 15108 564
rect 15160 552 15166 604
rect 143258 592 143264 604
rect 143219 564 143264 592
rect 143258 552 143264 564
rect 143316 552 143322 604
rect 195606 592 195612 604
rect 195567 564 195612 592
rect 195606 552 195612 564
rect 195664 552 195670 604
rect 203702 552 203708 604
rect 203760 592 203766 604
rect 203886 592 203892 604
rect 203760 564 203892 592
rect 203760 552 203766 564
rect 203886 552 203892 564
rect 203944 552 203950 604
rect 212258 552 212264 604
rect 212316 592 212322 604
rect 212445 595 212503 601
rect 212445 592 212457 595
rect 212316 564 212457 592
rect 212316 552 212322 564
rect 212445 561 212457 564
rect 212491 561 212503 595
rect 213454 592 213460 604
rect 213415 564 213460 592
rect 212445 555 212503 561
rect 213454 552 213460 564
rect 213512 552 213518 604
rect 316954 552 316960 604
rect 317012 592 317018 604
rect 317322 592 317328 604
rect 317012 564 317328 592
rect 317012 552 317018 564
rect 317322 552 317328 564
rect 317380 552 317386 604
rect 333606 592 333612 604
rect 333567 564 333612 592
rect 333606 552 333612 564
rect 333664 552 333670 604
rect 369946 552 369952 604
rect 370004 592 370010 604
rect 370406 592 370412 604
rect 370004 564 370412 592
rect 370004 552 370010 564
rect 370406 552 370412 564
rect 370464 552 370470 604
rect 485958 552 485964 604
rect 486016 592 486022 604
rect 486970 592 486976 604
rect 486016 564 486976 592
rect 486016 552 486022 564
rect 486970 552 486976 564
rect 487028 552 487034 604
rect 501046 552 501052 604
rect 501104 592 501110 604
rect 501230 592 501236 604
rect 501104 564 501236 592
rect 501104 552 501110 564
rect 501230 552 501236 564
rect 501288 552 501294 604
rect 503714 552 503720 604
rect 503772 592 503778 604
rect 504818 592 504824 604
rect 503772 564 504824 592
rect 503772 552 503778 564
rect 504818 552 504824 564
rect 504876 552 504882 604
rect 507946 552 507952 604
rect 508004 592 508010 604
rect 508406 592 508412 604
rect 508004 564 508412 592
rect 508004 552 508010 564
rect 508406 552 508412 564
rect 508464 552 508470 604
rect 514754 552 514760 604
rect 514812 592 514818 604
rect 515582 592 515588 604
rect 514812 564 515588 592
rect 514812 552 514818 564
rect 515582 552 515588 564
rect 515640 552 515646 604
rect 521654 552 521660 604
rect 521712 592 521718 604
rect 522666 592 522672 604
rect 521712 564 522672 592
rect 521712 552 521718 564
rect 522666 552 522672 564
rect 522724 552 522730 604
rect 525794 552 525800 604
rect 525852 592 525858 604
rect 526254 592 526260 604
rect 525852 564 526260 592
rect 525852 552 525858 564
rect 526254 552 526260 564
rect 526312 552 526318 604
rect 542354 552 542360 604
rect 542412 592 542418 604
rect 542906 592 542912 604
rect 542412 564 542912 592
rect 542412 552 542418 564
rect 542906 552 542912 564
rect 542964 552 542970 604
rect 543734 552 543740 604
rect 543792 592 543798 604
rect 544102 592 544108 604
rect 543792 564 544108 592
rect 543792 552 543798 564
rect 544102 552 544108 564
rect 544160 552 544166 604
<< via1 >>
rect 154120 700952 154172 701004
rect 333980 700952 334032 701004
rect 137836 700884 137888 700936
rect 329840 700884 329892 700936
rect 269028 700816 269080 700868
rect 462320 700816 462372 700868
rect 273168 700748 273220 700800
rect 478512 700748 478564 700800
rect 105452 700680 105504 700732
rect 338120 700680 338172 700732
rect 89168 700612 89220 700664
rect 347872 700612 347924 700664
rect 72976 700544 73028 700596
rect 343640 700544 343692 700596
rect 255228 700476 255280 700528
rect 527180 700476 527232 700528
rect 259368 700408 259420 700460
rect 543464 700408 543516 700460
rect 40500 700340 40552 700392
rect 351920 700340 351972 700392
rect 24308 700272 24360 700324
rect 360200 700272 360252 700324
rect 170312 700204 170364 700256
rect 325700 700204 325752 700256
rect 285588 700136 285640 700188
rect 413652 700136 413704 700188
rect 281448 700068 281500 700120
rect 397460 700068 397512 700120
rect 202788 700000 202840 700052
rect 317420 700000 317472 700052
rect 218980 699932 219032 699984
rect 321560 699932 321612 699984
rect 348792 699864 348844 699916
rect 267648 699796 267700 699848
rect 298008 699796 298060 699848
rect 300124 699796 300176 699848
rect 300768 699796 300820 699848
rect 293868 699728 293920 699780
rect 332508 699728 332560 699780
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 283840 699660 283892 699712
rect 309140 699660 309192 699712
rect 305000 699592 305052 699644
rect 242808 696940 242860 696992
rect 580172 696940 580224 696992
rect 364340 692792 364392 692844
rect 365076 692792 365128 692844
rect 246948 685856 247000 685908
rect 580172 685856 580224 685908
rect 364340 683068 364392 683120
rect 364616 683068 364668 683120
rect 3516 681708 3568 681760
rect 364432 681708 364484 681760
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 364340 673548 364392 673600
rect 364616 673548 364668 673600
rect 238668 673480 238720 673532
rect 580172 673480 580224 673532
rect 364340 668584 364392 668636
rect 364524 668584 364576 668636
rect 3424 667904 3476 667956
rect 372620 667904 372672 667956
rect 494152 666544 494204 666596
rect 288900 663280 288952 663332
rect 364524 663280 364576 663332
rect 235908 663212 235960 663264
rect 314108 663212 314160 663264
rect 276204 663144 276256 663196
rect 429292 663144 429344 663196
rect 263600 663076 263652 663128
rect 494152 663076 494204 663128
rect 250996 663008 251048 663060
rect 559012 663008 559064 663060
rect 300768 662804 300820 662856
rect 301504 662804 301556 662856
rect 204628 662736 204680 662788
rect 539876 662736 539928 662788
rect 192024 662668 192076 662720
rect 539968 662668 540020 662720
rect 8852 662600 8904 662652
rect 394148 662600 394200 662652
rect 9588 662532 9640 662584
rect 406752 662532 406804 662584
rect 175188 662464 175240 662516
rect 577504 662464 577556 662516
rect 9496 662396 9548 662448
rect 432052 662396 432104 662448
rect 95240 662328 95292 662380
rect 232596 662328 232648 662380
rect 233884 662328 233936 662380
rect 398380 662328 398432 662380
rect 208860 662260 208912 662312
rect 381636 662260 381688 662312
rect 230664 662192 230716 662244
rect 419356 662192 419408 662244
rect 213828 662124 213880 662176
rect 448888 662124 448940 662176
rect 112076 662056 112128 662108
rect 369124 662056 369176 662108
rect 196256 661988 196308 662040
rect 540060 661988 540112 662040
rect 107844 661920 107896 661972
rect 169760 661920 169812 661972
rect 183652 661920 183704 661972
rect 541716 661920 541768 661972
rect 91008 661852 91060 661904
rect 165896 661852 165948 661904
rect 170956 661852 171008 661904
rect 541624 661852 541676 661904
rect 166816 661784 166868 661836
rect 540888 661784 540940 661836
rect 120448 661716 120500 661768
rect 158720 661716 158772 661768
rect 162584 661716 162636 661768
rect 538772 661716 538824 661768
rect 154120 661648 154172 661700
rect 540796 661648 540848 661700
rect 82544 661580 82596 661632
rect 155684 661580 155736 661632
rect 158352 661580 158404 661632
rect 548524 661580 548576 661632
rect 53104 661512 53156 661564
rect 444656 661512 444708 661564
rect 145748 661444 145800 661496
rect 540612 661444 540664 661496
rect 141516 661376 141568 661428
rect 540704 661376 540756 661428
rect 54484 661308 54536 661360
rect 457260 661308 457312 661360
rect 457536 661308 457588 661360
rect 495164 661308 495216 661360
rect 4068 661240 4120 661292
rect 436192 661240 436244 661292
rect 448520 661240 448572 661292
rect 528836 661240 528888 661292
rect 103612 661172 103664 661224
rect 540244 661172 540296 661224
rect 9404 661104 9456 661156
rect 461492 661104 461544 661156
rect 9128 661036 9180 661088
rect 486792 661036 486844 661088
rect 3884 660968 3936 661020
rect 213828 660968 213880 661020
rect 225696 660968 225748 661020
rect 538404 660968 538456 661020
rect 213092 660900 213144 660952
rect 538496 660900 538548 660952
rect 200488 660832 200540 660884
rect 538588 660832 538640 660884
rect 187792 660764 187844 660816
rect 538680 660764 538732 660816
rect 8208 660696 8260 660748
rect 377312 660696 377364 660748
rect 8116 660628 8168 660680
rect 389916 660628 389968 660680
rect 149980 660560 150032 660612
rect 539508 660560 539560 660612
rect 8024 660492 8076 660544
rect 402520 660492 402572 660544
rect 7932 660424 7984 660476
rect 415216 660424 415268 660476
rect 169760 660356 169812 660408
rect 580724 660356 580776 660408
rect 158720 660288 158772 660340
rect 580908 660288 580960 660340
rect 133052 660220 133104 660272
rect 540428 660220 540480 660272
rect 58716 660152 58768 660204
rect 474096 660152 474148 660204
rect 7840 660084 7892 660136
rect 427820 660084 427872 660136
rect 7748 660016 7800 660068
rect 440240 660016 440292 660068
rect 99656 659948 99708 660000
rect 539140 659948 539192 660000
rect 7656 659880 7708 659932
rect 452660 659880 452712 659932
rect 7564 659812 7616 659864
rect 465356 659812 465408 659864
rect 9220 659744 9272 659796
rect 478052 659744 478104 659796
rect 6184 659676 6236 659728
rect 490564 659676 490616 659728
rect 3332 659608 3384 659660
rect 230664 659608 230716 659660
rect 368572 659651 368624 659660
rect 368572 659617 368581 659651
rect 368581 659617 368615 659651
rect 368615 659617 368624 659651
rect 368572 659608 368624 659617
rect 369124 659651 369176 659660
rect 369124 659617 369133 659651
rect 369133 659617 369167 659651
rect 369167 659617 369176 659651
rect 369124 659608 369176 659617
rect 381268 659651 381320 659660
rect 381268 659617 381277 659651
rect 381277 659617 381311 659651
rect 381311 659617 381320 659651
rect 381268 659608 381320 659617
rect 381636 659651 381688 659660
rect 381636 659617 381645 659651
rect 381645 659617 381679 659651
rect 381679 659617 381688 659651
rect 381636 659608 381688 659617
rect 385316 659651 385368 659660
rect 385316 659617 385325 659651
rect 385325 659617 385359 659651
rect 385359 659617 385368 659651
rect 385316 659608 385368 659617
rect 410708 659651 410760 659660
rect 410708 659617 410717 659651
rect 410717 659617 410751 659651
rect 410751 659617 410760 659651
rect 410708 659608 410760 659617
rect 423220 659651 423272 659660
rect 423220 659617 423229 659651
rect 423229 659617 423263 659651
rect 423263 659617 423272 659651
rect 423220 659608 423272 659617
rect 469588 659651 469640 659660
rect 469588 659617 469597 659651
rect 469597 659617 469631 659651
rect 469631 659617 469640 659651
rect 469588 659608 469640 659617
rect 3240 659540 3292 659592
rect 233884 659540 233936 659592
rect 234528 659540 234580 659592
rect 541900 659540 541952 659592
rect 230296 659472 230348 659524
rect 539692 659472 539744 659524
rect 221832 659404 221884 659456
rect 541808 659404 541860 659456
rect 179696 659379 179748 659388
rect 179696 659345 179705 659379
rect 179705 659345 179739 659379
rect 179739 659345 179748 659379
rect 179696 659336 179748 659345
rect 217600 659336 217652 659388
rect 539784 659336 539836 659388
rect 116584 659311 116636 659320
rect 116584 659277 116593 659311
rect 116593 659277 116627 659311
rect 116627 659277 116636 659311
rect 116584 659268 116636 659277
rect 125048 659311 125100 659320
rect 125048 659277 125057 659311
rect 125057 659277 125091 659311
rect 125091 659277 125100 659311
rect 125048 659268 125100 659277
rect 129280 659311 129332 659320
rect 129280 659277 129289 659311
rect 129289 659277 129323 659311
rect 129323 659277 129332 659311
rect 129280 659268 129332 659277
rect 137560 659311 137612 659320
rect 137560 659277 137569 659311
rect 137569 659277 137603 659311
rect 137603 659277 137612 659311
rect 137560 659268 137612 659277
rect 165896 659268 165948 659320
rect 580632 659268 580684 659320
rect 540152 659200 540204 659252
rect 8668 659132 8720 659184
rect 580816 659132 580868 659184
rect 8760 659064 8812 659116
rect 580172 659064 580224 659116
rect 5080 658996 5132 659048
rect 539416 658928 539468 658980
rect 4988 658860 5040 658912
rect 540520 658792 540572 658844
rect 539324 658724 539376 658776
rect 4896 658656 4948 658708
rect 540336 658588 540388 658640
rect 9312 658520 9364 658572
rect 3148 653556 3200 653608
rect 8668 653556 8720 653608
rect 539692 651312 539744 651364
rect 580080 651312 580132 651364
rect 541900 640228 541952 640280
rect 580080 640228 580132 640280
rect 539600 627852 539652 627904
rect 580080 627852 580132 627904
rect 3148 624860 3200 624912
rect 8208 624860 8260 624912
rect 2780 610444 2832 610496
rect 5080 610444 5132 610496
rect 539784 604392 539836 604444
rect 580080 604392 580132 604444
rect 3148 596028 3200 596080
rect 8760 596028 8812 596080
rect 541808 593308 541860 593360
rect 580080 593308 580132 593360
rect 538496 580932 538548 580984
rect 580080 580932 580132 580984
rect 3148 567536 3200 567588
rect 8116 567536 8168 567588
rect 539876 557472 539928 557524
rect 580080 557472 580132 557524
rect 3240 538772 3292 538824
rect 8852 538772 8904 538824
rect 538588 534012 538640 534064
rect 580172 534012 580224 534064
rect 539968 510552 540020 510604
rect 579804 510552 579856 510604
rect 3240 510008 3292 510060
rect 8024 510008 8076 510060
rect 540060 499468 540112 499520
rect 579988 499468 580040 499520
rect 2780 496680 2832 496732
rect 4988 496680 5040 496732
rect 538680 487092 538732 487144
rect 580172 487092 580224 487144
rect 3240 481176 3292 481228
rect 9588 481176 9640 481228
rect 540152 463632 540204 463684
rect 579804 463632 579856 463684
rect 541716 452548 541768 452600
rect 579988 452548 580040 452600
rect 3240 452412 3292 452464
rect 7932 452412 7984 452464
rect 577504 440172 577556 440224
rect 579712 440172 579764 440224
rect 2780 438744 2832 438796
rect 4896 438744 4948 438796
rect 540888 416712 540940 416764
rect 579804 416712 579856 416764
rect 541624 405628 541676 405680
rect 579988 405628 580040 405680
rect 3332 395224 3384 395276
rect 7840 395224 7892 395276
rect 538772 393252 538824 393304
rect 580172 393252 580224 393304
rect 540796 369792 540848 369844
rect 579804 369792 579856 369844
rect 3148 366664 3200 366716
rect 9496 366664 9548 366716
rect 548524 358708 548576 358760
rect 579988 358708 580040 358760
rect 539508 346332 539560 346384
rect 580172 346332 580224 346384
rect 3332 337492 3384 337544
rect 7748 337492 7800 337544
rect 540704 322872 540756 322924
rect 579804 322872 579856 322924
rect 540612 311788 540664 311840
rect 579988 311788 580040 311840
rect 3056 309068 3108 309120
rect 53104 309068 53156 309120
rect 539416 299412 539468 299464
rect 580172 299412 580224 299464
rect 3148 294788 3200 294840
rect 7656 294788 7708 294840
rect 3332 280100 3384 280152
rect 9404 280100 9456 280152
rect 540520 275952 540572 276004
rect 579804 275952 579856 276004
rect 3332 266296 3384 266348
rect 54484 266296 54536 266348
rect 540428 264868 540480 264920
rect 579988 264868 580040 264920
rect 539324 252492 539376 252544
rect 580172 252492 580224 252544
rect 3332 252220 3384 252272
rect 7564 252220 7616 252272
rect 3332 237328 3384 237380
rect 58716 237328 58768 237380
rect 540336 229032 540388 229084
rect 579804 229032 579856 229084
rect 3332 223048 3384 223100
rect 9312 223048 9364 223100
rect 3332 208156 3384 208208
rect 9220 208156 9272 208208
rect 3332 194488 3384 194540
rect 9128 194488 9180 194540
rect 540244 182112 540296 182164
rect 580172 182112 580224 182164
rect 3332 179596 3384 179648
rect 9036 179596 9088 179648
rect 3056 165452 3108 165504
rect 6184 165452 6236 165504
rect 539140 158652 539192 158704
rect 580172 158652 580224 158704
rect 3332 122748 3384 122800
rect 25504 122748 25556 122800
rect 539232 111732 539284 111784
rect 580172 111732 580224 111784
rect 3332 93780 3384 93832
rect 58624 93780 58676 93832
rect 538956 88272 539008 88324
rect 580172 88272 580224 88324
rect 3148 79092 3200 79144
rect 8944 79092 8996 79144
rect 539048 64812 539100 64864
rect 579620 64812 579672 64864
rect 2780 64540 2832 64592
rect 4804 64540 4856 64592
rect 60740 57944 60792 57996
rect 61660 57944 61712 57996
rect 44088 57876 44140 57928
rect 95240 57876 95292 57928
rect 108948 57876 109000 57928
rect 41328 57808 41380 57860
rect 93216 57808 93268 57860
rect 100668 57808 100720 57860
rect 38476 57740 38528 57792
rect 90364 57740 90416 57792
rect 96528 57740 96580 57792
rect 104164 57808 104216 57860
rect 111892 57808 111944 57860
rect 113088 57876 113140 57928
rect 152004 57876 152056 57928
rect 152464 57876 152516 57928
rect 156972 57876 157024 57928
rect 158628 57876 158680 57928
rect 189264 57876 189316 57928
rect 190368 57876 190420 57928
rect 215668 57876 215720 57928
rect 242164 57876 242216 57928
rect 245568 57876 245620 57928
rect 261760 57876 261812 57928
rect 263508 57876 263560 57928
rect 275468 57876 275520 57928
rect 280068 57876 280120 57928
rect 289176 57876 289228 57928
rect 460572 57876 460624 57928
rect 485964 57876 486016 57928
rect 497832 57876 497884 57928
rect 529204 57876 529256 57928
rect 149060 57808 149112 57860
rect 150348 57808 150400 57860
rect 182364 57808 182416 57860
rect 183468 57808 183520 57860
rect 214748 57808 214800 57860
rect 215208 57808 215260 57860
rect 236276 57808 236328 57860
rect 240048 57808 240100 57860
rect 256884 57808 256936 57860
rect 259368 57808 259420 57860
rect 272524 57808 272576 57860
rect 274548 57808 274600 57860
rect 285220 57808 285272 57860
rect 319444 57808 319496 57860
rect 321468 57808 321520 57860
rect 480168 57808 480220 57860
rect 489184 57808 489236 57860
rect 519360 57808 519412 57860
rect 520188 57808 520240 57860
rect 520372 57808 520424 57860
rect 521568 57808 521620 57860
rect 527180 57808 527232 57860
rect 528468 57808 528520 57860
rect 38568 57672 38620 57724
rect 91284 57672 91336 57724
rect 93768 57672 93820 57724
rect 142252 57740 142304 57792
rect 142804 57740 142856 57792
rect 151084 57740 151136 57792
rect 153844 57740 153896 57792
rect 155960 57740 156012 57792
rect 185308 57740 185360 57792
rect 186228 57740 186280 57792
rect 212724 57740 212776 57792
rect 221556 57740 221608 57792
rect 222108 57740 222160 57792
rect 235264 57740 235316 57792
rect 237288 57740 237340 57792
rect 253940 57740 253992 57792
rect 257988 57740 258040 57792
rect 271512 57740 271564 57792
rect 275928 57740 275980 57792
rect 286232 57740 286284 57792
rect 326988 57740 327040 57792
rect 328368 57740 328420 57792
rect 347964 57740 348016 57792
rect 349068 57740 349120 57792
rect 371424 57740 371476 57792
rect 374644 57740 374696 57792
rect 482100 57740 482152 57792
rect 482928 57740 482980 57792
rect 483112 57740 483164 57792
rect 484308 57740 484360 57792
rect 489000 57740 489052 57792
rect 489828 57740 489880 57792
rect 498752 57740 498804 57792
rect 532700 57808 532752 57860
rect 533068 57808 533120 57860
rect 530124 57740 530176 57792
rect 531228 57740 531280 57792
rect 534080 57740 534132 57792
rect 535368 57740 535420 57792
rect 537024 57808 537076 57860
rect 538128 57808 538180 57860
rect 541624 57740 541676 57792
rect 30196 57604 30248 57656
rect 78036 57604 78088 57656
rect 81532 57604 81584 57656
rect 85488 57604 85540 57656
rect 138296 57672 138348 57724
rect 139124 57672 139176 57724
rect 136364 57604 136416 57656
rect 140688 57604 140740 57656
rect 147588 57672 147640 57724
rect 180432 57672 180484 57724
rect 182088 57672 182140 57724
rect 209780 57672 209832 57724
rect 213828 57672 213880 57724
rect 232320 57672 232372 57724
rect 233148 57672 233200 57724
rect 250996 57672 251048 57724
rect 255228 57672 255280 57724
rect 269580 57672 269632 57724
rect 271696 57672 271748 57724
rect 282276 57672 282328 57724
rect 284208 57672 284260 57724
rect 293040 57672 293092 57724
rect 296628 57672 296680 57724
rect 302884 57672 302936 57724
rect 310428 57672 310480 57724
rect 314660 57672 314712 57724
rect 321468 57672 321520 57724
rect 323492 57672 323544 57724
rect 466460 57672 466512 57724
rect 494244 57672 494296 57724
rect 31668 57536 31720 57588
rect 85396 57536 85448 57588
rect 89628 57536 89680 57588
rect 122472 57536 122524 57588
rect 130476 57536 130528 57588
rect 133420 57536 133472 57588
rect 147128 57536 147180 57588
rect 23388 57468 23440 57520
rect 78588 57468 78640 57520
rect 21916 57400 21968 57452
rect 76564 57400 76616 57452
rect 83464 57468 83516 57520
rect 86408 57468 86460 57520
rect 86868 57468 86920 57520
rect 82084 57400 82136 57452
rect 92296 57400 92348 57452
rect 129464 57468 129516 57520
rect 132408 57468 132460 57520
rect 145196 57468 145248 57520
rect 124128 57400 124180 57452
rect 136548 57400 136600 57452
rect 173624 57604 173676 57656
rect 176568 57604 176620 57656
rect 203984 57604 204036 57656
rect 204168 57604 204220 57656
rect 227444 57604 227496 57656
rect 229008 57604 229060 57656
rect 247040 57604 247092 57656
rect 252468 57604 252520 57656
rect 266636 57604 266688 57656
rect 267648 57604 267700 57656
rect 279332 57604 279384 57656
rect 281448 57604 281500 57656
rect 291108 57604 291160 57656
rect 311808 57604 311860 57656
rect 315580 57604 315632 57656
rect 316684 57604 316736 57656
rect 317604 57604 317656 57656
rect 322848 57604 322900 57656
rect 325424 57604 325476 57656
rect 328368 57604 328420 57656
rect 329288 57604 329340 57656
rect 344008 57604 344060 57656
rect 344928 57604 344980 57656
rect 346952 57604 347004 57656
rect 347964 57604 348016 57656
rect 350908 57604 350960 57656
rect 351828 57604 351880 57656
rect 357716 57604 357768 57656
rect 358636 57604 358688 57656
rect 360660 57604 360712 57656
rect 362224 57604 362276 57656
rect 367560 57604 367612 57656
rect 368388 57604 368440 57656
rect 368480 57604 368532 57656
rect 369676 57604 369728 57656
rect 374368 57604 374420 57656
rect 375288 57604 375340 57656
rect 375380 57604 375432 57656
rect 376576 57604 376628 57656
rect 379244 57604 379296 57656
rect 380164 57604 380216 57656
rect 381268 57604 381320 57656
rect 382096 57604 382148 57656
rect 388076 57604 388128 57656
rect 389088 57604 389140 57656
rect 391020 57604 391072 57656
rect 391848 57604 391900 57656
rect 392032 57604 392084 57656
rect 393228 57604 393280 57656
rect 394976 57604 395028 57656
rect 395896 57604 395948 57656
rect 397920 57604 397972 57656
rect 398748 57604 398800 57656
rect 398840 57604 398892 57656
rect 400036 57604 400088 57656
rect 401784 57604 401836 57656
rect 402796 57604 402848 57656
rect 404728 57604 404780 57656
rect 405648 57604 405700 57656
rect 408684 57604 408736 57656
rect 409696 57604 409748 57656
rect 411628 57604 411680 57656
rect 412456 57604 412508 57656
rect 418436 57604 418488 57656
rect 419448 57604 419500 57656
rect 421380 57604 421432 57656
rect 422208 57604 422260 57656
rect 422392 57604 422444 57656
rect 423496 57604 423548 57656
rect 425336 57604 425388 57656
rect 426256 57604 426308 57656
rect 428280 57604 428332 57656
rect 429108 57604 429160 57656
rect 432144 57604 432196 57656
rect 433156 57604 433208 57656
rect 435088 57604 435140 57656
rect 436008 57604 436060 57656
rect 439044 57604 439096 57656
rect 440148 57604 440200 57656
rect 441988 57604 442040 57656
rect 442908 57604 442960 57656
rect 448796 57604 448848 57656
rect 449716 57604 449768 57656
rect 451740 57604 451792 57656
rect 452568 57604 452620 57656
rect 452752 57604 452804 57656
rect 453948 57604 454000 57656
rect 455696 57604 455748 57656
rect 456708 57604 456760 57656
rect 458640 57604 458692 57656
rect 459468 57604 459520 57656
rect 459560 57604 459612 57656
rect 460848 57604 460900 57656
rect 462504 57604 462556 57656
rect 463608 57604 463660 57656
rect 465448 57604 465500 57656
rect 466368 57604 466420 57656
rect 469404 57604 469456 57656
rect 496912 57672 496964 57724
rect 512460 57672 512512 57724
rect 547144 57672 547196 57724
rect 496820 57604 496872 57656
rect 498108 57604 498160 57656
rect 499764 57604 499816 57656
rect 500868 57604 500920 57656
rect 502708 57604 502760 57656
rect 503628 57604 503680 57656
rect 505652 57604 505704 57656
rect 506388 57604 506440 57656
rect 513472 57604 513524 57656
rect 514576 57604 514628 57656
rect 515404 57604 515456 57656
rect 549904 57604 549956 57656
rect 176476 57536 176528 57588
rect 183376 57536 183428 57588
rect 184848 57536 184900 57588
rect 208860 57536 208912 57588
rect 211068 57536 211120 57588
rect 233332 57536 233384 57588
rect 237196 57536 237248 57588
rect 254860 57536 254912 57588
rect 256608 57536 256660 57588
rect 270592 57536 270644 57588
rect 273168 57536 273220 57588
rect 284300 57536 284352 57588
rect 286968 57536 287020 57588
rect 295064 57536 295116 57588
rect 309048 57536 309100 57588
rect 313648 57536 313700 57588
rect 317328 57536 317380 57588
rect 320548 57536 320600 57588
rect 322756 57536 322808 57588
rect 324412 57536 324464 57588
rect 349896 57536 349948 57588
rect 352012 57536 352064 57588
rect 361672 57536 361724 57588
rect 362776 57536 362828 57588
rect 364616 57536 364668 57588
rect 369952 57536 370004 57588
rect 378324 57536 378376 57588
rect 379428 57536 379480 57588
rect 429200 57536 429252 57588
rect 430488 57536 430540 57588
rect 473360 57536 473412 57588
rect 474556 57536 474608 57588
rect 475292 57536 475344 57588
rect 503720 57536 503772 57588
rect 506664 57536 506716 57588
rect 177488 57468 177540 57520
rect 15108 57332 15160 57384
rect 64972 57332 65024 57384
rect 65524 57332 65576 57384
rect 70768 57332 70820 57384
rect 71044 57332 71096 57384
rect 79508 57332 79560 57384
rect 12348 57264 12400 57316
rect 68744 57264 68796 57316
rect 71136 57264 71188 57316
rect 75644 57264 75696 57316
rect 75828 57264 75880 57316
rect 82728 57332 82780 57384
rect 79968 57264 80020 57316
rect 124588 57332 124640 57384
rect 13636 57196 13688 57248
rect 71688 57196 71740 57248
rect 73804 57196 73856 57248
rect 74632 57196 74684 57248
rect 75184 57196 75236 57248
rect 82452 57196 82504 57248
rect 115204 57196 115256 57248
rect 118700 57196 118752 57248
rect 126152 57332 126204 57384
rect 126244 57332 126296 57384
rect 139308 57332 139360 57384
rect 174544 57400 174596 57452
rect 175188 57400 175240 57452
rect 211804 57468 211856 57520
rect 218612 57468 218664 57520
rect 219256 57468 219308 57520
rect 240232 57468 240284 57520
rect 241428 57468 241480 57520
rect 257804 57468 257856 57520
rect 260748 57468 260800 57520
rect 273536 57468 273588 57520
rect 277308 57468 277360 57520
rect 287244 57468 287296 57520
rect 289728 57468 289780 57520
rect 298008 57468 298060 57520
rect 299388 57468 299440 57520
rect 305828 57468 305880 57520
rect 306288 57468 306340 57520
rect 311716 57468 311768 57520
rect 320088 57468 320140 57520
rect 322480 57468 322532 57520
rect 478236 57468 478288 57520
rect 507952 57468 508004 57520
rect 509516 57468 509568 57520
rect 538956 57536 539008 57588
rect 544384 57536 544436 57588
rect 542360 57468 542412 57520
rect 177948 57400 178000 57452
rect 205916 57400 205968 57452
rect 206744 57400 206796 57452
rect 229376 57400 229428 57452
rect 230480 57400 230532 57452
rect 248972 57400 249024 57452
rect 251088 57400 251140 57452
rect 265624 57400 265676 57452
rect 266268 57400 266320 57452
rect 278412 57400 278464 57452
rect 282828 57400 282880 57452
rect 292120 57400 292172 57452
rect 292488 57400 292540 57452
rect 299940 57400 299992 57452
rect 472348 57400 472400 57452
rect 501052 57400 501104 57452
rect 507584 57400 507636 57452
rect 543740 57400 543792 57452
rect 171600 57332 171652 57384
rect 179328 57332 179380 57384
rect 202972 57332 203024 57384
rect 205548 57332 205600 57384
rect 228456 57332 228508 57384
rect 125508 57196 125560 57248
rect 161848 57264 161900 57316
rect 168380 57264 168432 57316
rect 169300 57264 169352 57316
rect 194140 57264 194192 57316
rect 200028 57264 200080 57316
rect 223580 57264 223632 57316
rect 230388 57332 230440 57384
rect 231768 57332 231820 57384
rect 249984 57332 250036 57384
rect 253756 57332 253808 57384
rect 268568 57332 268620 57384
rect 271788 57332 271840 57384
rect 283288 57332 283340 57384
rect 285588 57332 285640 57384
rect 294052 57332 294104 57384
rect 295248 57332 295300 57384
rect 301872 57332 301924 57384
rect 304908 57332 304960 57384
rect 309692 57332 309744 57384
rect 384212 57332 384264 57384
rect 384948 57332 385000 57384
rect 414572 57332 414624 57384
rect 415308 57332 415360 57384
rect 444932 57332 444984 57384
rect 445668 57332 445720 57384
rect 457628 57332 457680 57384
rect 483112 57332 483164 57384
rect 484124 57332 484176 57384
rect 514760 57332 514812 57384
rect 516416 57332 516468 57384
rect 554872 57332 554924 57384
rect 228916 57264 228968 57316
rect 248052 57264 248104 57316
rect 248328 57264 248380 57316
rect 263692 57264 263744 57316
rect 264888 57264 264940 57316
rect 277400 57264 277452 57316
rect 278688 57264 278740 57316
rect 288164 57264 288216 57316
rect 288256 57264 288308 57316
rect 296996 57264 297048 57316
rect 298008 57264 298060 57316
rect 304816 57264 304868 57316
rect 306196 57264 306248 57316
rect 310704 57264 310756 57316
rect 463516 57264 463568 57316
rect 490104 57264 490156 57316
rect 492864 57264 492916 57316
rect 525800 57264 525852 57316
rect 528192 57264 528244 57316
rect 566464 57264 566516 57316
rect 160836 57196 160888 57248
rect 168196 57196 168248 57248
rect 198096 57196 198148 57248
rect 198648 57196 198700 57248
rect 222568 57196 222620 57248
rect 223488 57196 223540 57248
rect 243084 57196 243136 57248
rect 244188 57196 244240 57248
rect 259736 57196 259788 57248
rect 263416 57196 263468 57248
rect 276388 57196 276440 57248
rect 279976 57196 280028 57248
rect 290188 57196 290240 57248
rect 293868 57196 293920 57248
rect 300952 57196 301004 57248
rect 315948 57196 316000 57248
rect 319536 57196 319588 57248
rect 354772 57196 354824 57248
rect 355876 57196 355928 57248
rect 385132 57196 385184 57248
rect 386328 57196 386380 57248
rect 415492 57196 415544 57248
rect 416688 57196 416740 57248
rect 437112 57196 437164 57248
rect 458272 57196 458324 57248
rect 479156 57196 479208 57248
rect 480168 57196 480220 57248
rect 481180 57196 481232 57248
rect 512092 57196 512144 57248
rect 525248 57196 525300 57248
rect 564440 57196 564492 57248
rect 37188 57128 37240 57180
rect 89352 57128 89404 57180
rect 97172 57128 97224 57180
rect 102876 57128 102928 57180
rect 106004 57128 106056 57180
rect 107568 57128 107620 57180
rect 142068 57128 142120 57180
rect 153108 57128 153160 57180
rect 157248 57128 157300 57180
rect 188252 57128 188304 57180
rect 188988 57128 189040 57180
rect 220636 57128 220688 57180
rect 220728 57128 220780 57180
rect 241152 57128 241204 57180
rect 246948 57128 247000 57180
rect 262680 57128 262732 57180
rect 269028 57128 269080 57180
rect 280344 57128 280396 57180
rect 494888 57128 494940 57180
rect 526444 57128 526496 57180
rect 529112 57128 529164 57180
rect 537484 57128 537536 57180
rect 545764 57128 545816 57180
rect 45468 57060 45520 57112
rect 96160 57060 96212 57112
rect 112812 57060 112864 57112
rect 117228 57060 117280 57112
rect 154948 57060 155000 57112
rect 156604 57060 156656 57112
rect 159824 57060 159876 57112
rect 160008 57060 160060 57112
rect 191196 57060 191248 57112
rect 193128 57060 193180 57112
rect 217692 57060 217744 57112
rect 219348 57060 219400 57112
rect 239220 57060 239272 57112
rect 242808 57060 242860 57112
rect 258816 57060 258868 57112
rect 262128 57060 262180 57112
rect 274456 57060 274508 57112
rect 297916 57060 297968 57112
rect 303896 57060 303948 57112
rect 353852 57060 353904 57112
rect 356152 57060 356204 57112
rect 405740 57060 405792 57112
rect 406936 57060 406988 57112
rect 436100 57060 436152 57112
rect 437388 57060 437440 57112
rect 445852 57060 445904 57112
rect 446956 57060 447008 57112
rect 490012 57060 490064 57112
rect 521660 57060 521712 57112
rect 526168 57060 526220 57112
rect 533344 57060 533396 57112
rect 50988 56992 51040 57044
rect 101128 56992 101180 57044
rect 105544 56992 105596 57044
rect 117780 56992 117832 57044
rect 117964 56992 118016 57044
rect 119988 56992 120040 57044
rect 157892 56992 157944 57044
rect 159916 56992 159968 57044
rect 190276 56992 190328 57044
rect 197268 56992 197320 57044
rect 217968 56992 218020 57044
rect 238208 56992 238260 57044
rect 238668 56992 238720 57044
rect 255872 56992 255924 57044
rect 270408 56992 270460 57044
rect 281356 56992 281408 57044
rect 495808 56992 495860 57044
rect 528744 56992 528796 57044
rect 46848 56924 46900 56976
rect 91744 56924 91796 56976
rect 98184 56924 98236 56976
rect 108580 56924 108632 56976
rect 111064 56924 111116 56976
rect 121276 56924 121328 56976
rect 121368 56924 121420 56976
rect 158904 56924 158956 56976
rect 165528 56924 165580 56976
rect 195152 56924 195204 56976
rect 202696 56924 202748 56976
rect 225512 56924 225564 56976
rect 227628 56924 227680 56976
rect 246028 56924 246080 56976
rect 249708 56924 249760 56976
rect 264704 56924 264756 56976
rect 288348 56924 288400 56976
rect 295984 56924 296036 56976
rect 345020 56924 345072 56976
rect 346308 56924 346360 56976
rect 476212 56924 476264 56976
rect 477408 56924 477460 56976
rect 486056 56924 486108 56976
rect 491944 56924 491996 56976
rect 535000 56924 535052 56976
rect 538956 56924 539008 56976
rect 61384 56856 61436 56908
rect 62856 56856 62908 56908
rect 107016 56856 107068 56908
rect 114468 56856 114520 56908
rect 153016 56856 153068 56908
rect 164148 56856 164200 56908
rect 172428 56856 172480 56908
rect 201040 56856 201092 56908
rect 201408 56856 201460 56908
rect 224500 56856 224552 56908
rect 224868 56856 224920 56908
rect 244096 56856 244148 56908
rect 245476 56856 245528 56908
rect 260380 56856 260432 56908
rect 307668 56856 307720 56908
rect 312636 56856 312688 56908
rect 53748 56788 53800 56840
rect 103060 56788 103112 56840
rect 112444 56788 112496 56840
rect 135904 56788 135956 56840
rect 57888 56720 57940 56772
rect 64788 56720 64840 56772
rect 61476 56652 61528 56704
rect 66812 56652 66864 56704
rect 67548 56652 67600 56704
rect 60648 56584 60700 56636
rect 102784 56652 102836 56704
rect 104072 56652 104124 56704
rect 108304 56720 108356 56772
rect 109868 56720 109920 56772
rect 119344 56720 119396 56772
rect 141240 56720 141292 56772
rect 114836 56652 114888 56704
rect 120724 56652 120776 56704
rect 122104 56652 122156 56704
rect 109684 56584 109736 56636
rect 115756 56584 115808 56636
rect 122196 56584 122248 56636
rect 77944 56516 77996 56568
rect 135352 56584 135404 56636
rect 143448 56788 143500 56840
rect 168288 56788 168340 56840
rect 197084 56788 197136 56840
rect 209688 56788 209740 56840
rect 231400 56788 231452 56840
rect 234528 56788 234580 56840
rect 251916 56788 251968 56840
rect 253848 56788 253900 56840
rect 267372 56788 267424 56840
rect 536012 56788 536064 56840
rect 536748 56788 536800 56840
rect 171048 56720 171100 56772
rect 199660 56720 199712 56772
rect 144184 56652 144236 56704
rect 148140 56652 148192 56704
rect 169024 56652 169076 56704
rect 206928 56652 206980 56704
rect 145564 56584 145616 56636
rect 154028 56584 154080 56636
rect 160744 56584 160796 56636
rect 162768 56584 162820 56636
rect 164884 56584 164936 56636
rect 173164 56584 173216 56636
rect 192208 56584 192260 56636
rect 194508 56584 194560 56636
rect 212448 56720 212500 56772
rect 234344 56720 234396 56772
rect 235908 56720 235960 56772
rect 252928 56720 252980 56772
rect 302148 56720 302200 56772
rect 307760 56720 307812 56772
rect 313188 56720 313240 56772
rect 316592 56720 316644 56772
rect 208308 56652 208360 56704
rect 226248 56652 226300 56704
rect 245108 56652 245160 56704
rect 303528 56652 303580 56704
rect 308772 56652 308824 56704
rect 315304 56652 315356 56704
rect 318524 56652 318576 56704
rect 324228 56652 324280 56704
rect 326344 56652 326396 56704
rect 342996 56652 343048 56704
rect 343732 56652 343784 56704
rect 504088 56652 504140 56704
rect 509884 56652 509936 56704
rect 523316 56652 523368 56704
rect 524328 56652 524380 56704
rect 210976 56584 211028 56636
rect 216588 56584 216640 56636
rect 237012 56584 237064 56636
rect 291108 56584 291160 56636
rect 298928 56584 298980 56636
rect 304264 56584 304316 56636
rect 306840 56584 306892 56636
rect 327356 56584 327408 56636
rect 336740 56584 336792 56636
rect 337200 56584 337252 56636
rect 338120 56584 338172 56636
rect 338212 56584 338264 56636
rect 537944 56584 537996 56636
rect 540244 56584 540296 56636
rect 186320 56516 186372 56568
rect 326344 56516 326396 56568
rect 336740 56491 336792 56500
rect 336740 56457 336749 56491
rect 336749 56457 336783 56491
rect 336783 56457 336792 56491
rect 336740 56448 336792 56457
rect 165620 55836 165672 55888
rect 166356 55836 166408 55888
rect 334348 55564 334400 55616
rect 101220 52300 101272 52352
rect 121736 51552 121788 51604
rect 98552 48331 98604 48340
rect 98552 48297 98561 48331
rect 98561 48297 98595 48331
rect 98595 48297 98604 48331
rect 98552 48288 98604 48297
rect 100852 48331 100904 48340
rect 100852 48297 100861 48331
rect 100861 48297 100895 48331
rect 100895 48297 100904 48331
rect 100852 48288 100904 48297
rect 121552 48331 121604 48340
rect 121552 48297 121561 48331
rect 121561 48297 121595 48331
rect 121595 48297 121604 48331
rect 121552 48288 121604 48297
rect 129004 48288 129056 48340
rect 145196 48288 145248 48340
rect 145288 48288 145340 48340
rect 195888 48288 195940 48340
rect 212632 48288 212684 48340
rect 213460 48288 213512 48340
rect 334164 48331 334216 48340
rect 334164 48297 334173 48331
rect 334173 48297 334207 48331
rect 334207 48297 334216 48331
rect 334164 48288 334216 48297
rect 98644 48220 98696 48272
rect 100116 48220 100168 48272
rect 98552 46971 98604 46980
rect 98552 46937 98561 46971
rect 98561 46937 98595 46971
rect 98595 46937 98604 46971
rect 98552 46928 98604 46937
rect 336740 46971 336792 46980
rect 336740 46937 336749 46971
rect 336749 46937 336783 46971
rect 336783 46937 336792 46971
rect 336740 46928 336792 46937
rect 338120 46903 338172 46912
rect 338120 46869 338129 46903
rect 338129 46869 338163 46903
rect 338163 46869 338172 46903
rect 338120 46860 338172 46869
rect 121460 41352 121512 41404
rect 121644 41352 121696 41404
rect 212540 41352 212592 41404
rect 212724 41352 212776 41404
rect 145012 38632 145064 38684
rect 145104 38632 145156 38684
rect 101036 38607 101088 38616
rect 101036 38573 101045 38607
rect 101045 38573 101079 38607
rect 101079 38573 101088 38607
rect 101036 38564 101088 38573
rect 192116 38564 192168 38616
rect 195888 38607 195940 38616
rect 195888 38573 195897 38607
rect 195897 38573 195931 38607
rect 195931 38573 195940 38607
rect 195888 38564 195940 38573
rect 98276 37952 98328 38004
rect 98460 37952 98512 38004
rect 338120 37315 338172 37324
rect 338120 37281 338129 37315
rect 338129 37281 338163 37315
rect 338163 37281 338172 37315
rect 338120 37272 338172 37281
rect 128820 37204 128872 37256
rect 336740 37247 336792 37256
rect 336740 37213 336749 37247
rect 336749 37213 336783 37247
rect 336783 37213 336792 37247
rect 336740 37204 336792 37213
rect 145012 35751 145064 35760
rect 145012 35717 145021 35751
rect 145021 35717 145055 35751
rect 145055 35717 145064 35751
rect 145012 35708 145064 35717
rect 121644 31764 121696 31816
rect 333980 31764 334032 31816
rect 101220 31628 101272 31680
rect 121736 31628 121788 31680
rect 334072 31628 334124 31680
rect 145196 28976 145248 29028
rect 192024 29019 192076 29028
rect 192024 28985 192033 29019
rect 192033 28985 192067 29019
rect 192067 28985 192076 29019
rect 192024 28976 192076 28985
rect 195888 29019 195940 29028
rect 195888 28985 195897 29019
rect 195897 28985 195931 29019
rect 195931 28985 195940 29019
rect 195888 28976 195940 28985
rect 98000 28908 98052 28960
rect 98460 28908 98512 28960
rect 100760 28908 100812 28960
rect 101220 28908 101272 28960
rect 128636 27727 128688 27736
rect 128636 27693 128645 27727
rect 128645 27693 128679 27727
rect 128679 27693 128688 27727
rect 128636 27684 128688 27693
rect 336740 27659 336792 27668
rect 336740 27625 336749 27659
rect 336749 27625 336783 27659
rect 336783 27625 336792 27659
rect 336740 27616 336792 27625
rect 121736 27548 121788 27600
rect 128636 27548 128688 27600
rect 212540 27591 212592 27600
rect 212540 27557 212549 27591
rect 212549 27557 212583 27591
rect 212583 27557 212592 27591
rect 212540 27548 212592 27557
rect 338120 27591 338172 27600
rect 338120 27557 338129 27591
rect 338129 27557 338163 27591
rect 338163 27557 338172 27591
rect 338120 27548 338172 27557
rect 2872 22040 2924 22092
rect 538036 22040 538088 22092
rect 195888 19456 195940 19508
rect 145012 19320 145064 19372
rect 145104 19320 145156 19372
rect 195888 19320 195940 19372
rect 192208 19295 192260 19304
rect 192208 19261 192217 19295
rect 192217 19261 192251 19295
rect 192251 19261 192260 19295
rect 192208 19252 192260 19261
rect 128912 19227 128964 19236
rect 128912 19193 128921 19227
rect 128921 19193 128955 19227
rect 128955 19193 128964 19227
rect 128912 19184 128964 19193
rect 121644 18003 121696 18012
rect 121644 17969 121653 18003
rect 121653 17969 121687 18003
rect 121687 17969 121696 18003
rect 121644 17960 121696 17969
rect 212632 17960 212684 18012
rect 333980 17935 334032 17944
rect 333980 17901 333989 17935
rect 333989 17901 334023 17935
rect 334023 17901 334032 17935
rect 333980 17892 334032 17901
rect 336740 17935 336792 17944
rect 336740 17901 336749 17935
rect 336749 17901 336783 17935
rect 336783 17901 336792 17935
rect 336740 17892 336792 17901
rect 538864 17892 538916 17944
rect 579804 17892 579856 17944
rect 203708 13132 203760 13184
rect 204168 13132 204220 13184
rect 121644 12452 121696 12504
rect 128912 12452 128964 12504
rect 121552 12384 121604 12436
rect 128912 12316 128964 12368
rect 192300 9664 192352 9716
rect 338304 9664 338356 9716
rect 195888 9596 195940 9648
rect 212448 9639 212500 9648
rect 212448 9605 212457 9639
rect 212457 9605 212491 9639
rect 212491 9605 212500 9639
rect 212448 9596 212500 9605
rect 337108 9528 337160 9580
rect 334072 8304 334124 8356
rect 111064 6332 111116 6384
rect 94504 6196 94556 6248
rect 136640 6196 136692 6248
rect 87328 6128 87380 6180
rect 131212 6128 131264 6180
rect 51632 5448 51684 5500
rect 100944 5448 100996 5500
rect 105176 5448 105228 5500
rect 145104 5448 145156 5500
rect 521384 5448 521436 5500
rect 521568 5448 521620 5500
rect 58808 5380 58860 5432
rect 107752 5380 107804 5432
rect 48136 5312 48188 5364
rect 98184 5312 98236 5364
rect 101588 5312 101640 5364
rect 142344 5312 142396 5364
rect 30288 5244 30340 5296
rect 84292 5244 84344 5296
rect 90916 5244 90968 5296
rect 133880 5244 133932 5296
rect 12440 5176 12492 5228
rect 69020 5176 69072 5228
rect 76656 5176 76708 5228
rect 121552 5176 121604 5228
rect 155132 5176 155184 5228
rect 186412 5176 186464 5228
rect 502248 5176 502300 5228
rect 536932 5176 536984 5228
rect 22008 5108 22060 5160
rect 77392 5108 77444 5160
rect 80244 5108 80296 5160
rect 125600 5108 125652 5160
rect 148048 5108 148100 5160
rect 180800 5108 180852 5160
rect 505008 5108 505060 5160
rect 540520 5108 540572 5160
rect 17224 5040 17276 5092
rect 73160 5040 73212 5092
rect 83832 5040 83884 5092
rect 128452 5040 128504 5092
rect 134892 5040 134944 5092
rect 169760 5040 169812 5092
rect 510528 5040 510580 5092
rect 547696 5040 547748 5092
rect 2872 4972 2924 5024
rect 60740 4972 60792 5024
rect 69480 4972 69532 5024
rect 115940 4972 115992 5024
rect 131396 4972 131448 5024
rect 167000 4972 167052 5024
rect 514576 4972 514628 5024
rect 551192 4972 551244 5024
rect 7656 4904 7708 4956
rect 64972 4904 65024 4956
rect 73068 4904 73120 4956
rect 118792 4904 118844 4956
rect 132592 4904 132644 4956
rect 168472 4904 168524 4956
rect 520188 4904 520240 4956
rect 558368 4904 558420 4956
rect 572 4836 624 4888
rect 59360 4836 59412 4888
rect 65984 4836 66036 4888
rect 113180 4836 113232 4888
rect 127808 4836 127860 4888
rect 164240 4836 164292 4888
rect 522948 4836 523000 4888
rect 561956 4836 562008 4888
rect 1676 4768 1728 4820
rect 60832 4768 60884 4820
rect 62396 4768 62448 4820
rect 110420 4768 110472 4820
rect 129004 4768 129056 4820
rect 165712 4768 165764 4820
rect 487068 4768 487120 4820
rect 519084 4768 519136 4820
rect 531136 4768 531188 4820
rect 572628 4768 572680 4820
rect 55220 4700 55272 4752
rect 104992 4700 105044 4752
rect 98092 4632 98144 4684
rect 139400 4632 139452 4684
rect 356152 4224 356204 4276
rect 357348 4224 357400 4276
rect 61384 4156 61436 4208
rect 20720 4088 20772 4140
rect 21916 4088 21968 4140
rect 71136 4088 71188 4140
rect 74264 4088 74316 4140
rect 93308 4088 93360 4140
rect 93768 4088 93820 4140
rect 95700 4088 95752 4140
rect 96528 4088 96580 4140
rect 112352 4088 112404 4140
rect 113088 4088 113140 4140
rect 113548 4088 113600 4140
rect 114468 4088 114520 4140
rect 119436 4088 119488 4140
rect 119988 4088 120040 4140
rect 120632 4088 120684 4140
rect 121368 4088 121420 4140
rect 123024 4088 123076 4140
rect 124128 4088 124180 4140
rect 136088 4088 136140 4140
rect 136548 4088 136600 4140
rect 138480 4088 138532 4140
rect 139308 4088 139360 4140
rect 140872 4088 140924 4140
rect 145656 4088 145708 4140
rect 146208 4088 146260 4140
rect 453948 4156 454000 4208
rect 175372 4088 175424 4140
rect 193220 4088 193272 4140
rect 194508 4088 194560 4140
rect 196808 4088 196860 4140
rect 197268 4088 197320 4140
rect 199200 4088 199252 4140
rect 200028 4088 200080 4140
rect 201500 4088 201552 4140
rect 202696 4088 202748 4140
rect 205088 4088 205140 4140
rect 205548 4088 205600 4140
rect 207480 4088 207532 4140
rect 208308 4088 208360 4140
rect 208676 4088 208728 4140
rect 209688 4088 209740 4140
rect 214656 4088 214708 4140
rect 215208 4088 215260 4140
rect 332416 4088 332468 4140
rect 332692 4088 332744 4140
rect 335360 4088 335412 4140
rect 335912 4088 335964 4140
rect 339500 4088 339552 4140
rect 340696 4088 340748 4140
rect 344928 4088 344980 4140
rect 345480 4088 345532 4140
rect 353208 4088 353260 4140
rect 356152 4088 356204 4140
rect 357440 4088 357492 4140
rect 360936 4088 360988 4140
rect 362224 4088 362276 4140
rect 365720 4088 365772 4140
rect 379428 4088 379480 4140
rect 387064 4088 387116 4140
rect 397368 4088 397420 4140
rect 409604 4088 409656 4140
rect 409696 4088 409748 4140
rect 423956 4088 424008 4140
rect 430396 4088 430448 4140
rect 431868 4088 431920 4140
rect 451280 4088 451332 4140
rect 452568 4088 452620 4140
rect 476304 4088 476356 4140
rect 484308 4088 484360 4140
rect 514392 4088 514444 4140
rect 514668 4088 514720 4140
rect 552388 4088 552440 4140
rect 566464 4088 566516 4140
rect 569040 4088 569092 4140
rect 111156 4020 111208 4072
rect 142804 4020 142856 4072
rect 144460 4020 144512 4072
rect 178040 4020 178092 4072
rect 190828 4020 190880 4072
rect 362776 4020 362828 4072
rect 366916 4020 366968 4072
rect 384948 4020 385000 4072
rect 394240 4020 394292 4072
rect 395896 4020 395948 4072
rect 407304 4020 407356 4072
rect 412456 4020 412508 4072
rect 427544 4020 427596 4072
rect 430488 4020 430540 4072
rect 448980 4020 449032 4072
rect 449716 4020 449768 4072
rect 472716 4020 472768 4072
rect 474556 4020 474608 4072
rect 502432 4020 502484 4072
rect 503628 4020 503680 4072
rect 8852 3952 8904 4004
rect 61476 3952 61528 4004
rect 63592 3952 63644 4004
rect 104164 3952 104216 4004
rect 121828 3952 121880 4004
rect 156604 3952 156656 4004
rect 160744 3952 160796 4004
rect 161112 3952 161164 4004
rect 183744 3952 183796 4004
rect 209872 3952 209924 4004
rect 313372 3952 313424 4004
rect 316684 3952 316736 4004
rect 386328 3952 386380 4004
rect 395436 3952 395488 4004
rect 400036 3952 400088 4004
rect 412088 3952 412140 4004
rect 412548 3952 412600 4004
rect 428740 3952 428792 4004
rect 429108 3952 429160 4004
rect 447784 3952 447836 4004
rect 449808 3952 449860 4004
rect 473912 3952 473964 4004
rect 477316 3952 477368 4004
rect 507216 3952 507268 4004
rect 526444 3952 526496 4004
rect 528652 3952 528704 4004
rect 531228 4020 531280 4072
rect 538956 4020 539008 4072
rect 577412 4020 577464 4072
rect 563152 3952 563204 4004
rect 16028 3884 16080 3936
rect 33876 3884 33928 3936
rect 86960 3884 87012 3936
rect 92112 3884 92164 3936
rect 112444 3884 112496 3936
rect 118240 3884 118292 3936
rect 149244 3884 149296 3936
rect 150348 3884 150400 3936
rect 153936 3884 153988 3936
rect 169024 3884 169076 3936
rect 173164 3884 173216 3936
rect 198832 3884 198884 3936
rect 216680 3884 216732 3936
rect 382188 3884 382240 3936
rect 391756 3884 391808 3936
rect 393136 3884 393188 3936
rect 404912 3884 404964 3936
rect 407028 3884 407080 3936
rect 421564 3884 421616 3936
rect 423496 3884 423548 3936
rect 440608 3884 440660 3936
rect 441528 3884 441580 3936
rect 19524 3816 19576 3868
rect 34980 3816 35032 3868
rect 88340 3816 88392 3868
rect 93860 3816 93912 3868
rect 96896 3816 96948 3868
rect 126244 3816 126296 3868
rect 130200 3816 130252 3868
rect 165620 3816 165672 3868
rect 180156 3816 180208 3868
rect 207020 3816 207072 3868
rect 360108 3816 360160 3868
rect 364524 3816 364576 3868
rect 369768 3816 369820 3868
rect 376392 3816 376444 3868
rect 383568 3816 383620 3868
rect 393044 3816 393096 3868
rect 393228 3816 393280 3868
rect 403716 3816 403768 3868
rect 404268 3816 404320 3868
rect 417976 3816 418028 3868
rect 418068 3816 418120 3868
rect 434536 3816 434588 3868
rect 434628 3816 434680 3868
rect 454868 3816 454920 3868
rect 462044 3884 462096 3936
rect 464988 3884 465040 3936
rect 491760 3884 491812 3936
rect 492588 3884 492640 3936
rect 525064 3884 525116 3936
rect 528468 3884 528520 3936
rect 567844 3884 567896 3936
rect 456708 3816 456760 3868
rect 462228 3816 462280 3868
rect 488172 3816 488224 3868
rect 489828 3816 489880 3868
rect 521476 3816 521528 3868
rect 524328 3816 524380 3868
rect 564348 3816 564400 3868
rect 25504 3748 25556 3800
rect 80060 3748 80112 3800
rect 10048 3680 10100 3732
rect 11244 3544 11296 3596
rect 12348 3544 12400 3596
rect 18328 3680 18380 3732
rect 75184 3680 75236 3732
rect 89720 3748 89772 3800
rect 122196 3748 122248 3800
rect 133788 3748 133840 3800
rect 168380 3748 168432 3800
rect 172980 3748 173032 3800
rect 201684 3748 201736 3800
rect 371148 3748 371200 3800
rect 377588 3748 377640 3800
rect 380808 3748 380860 3800
rect 389456 3748 389508 3800
rect 390468 3748 390520 3800
rect 401324 3748 401376 3800
rect 401508 3748 401560 3800
rect 414480 3748 414532 3800
rect 415308 3748 415360 3800
rect 431132 3748 431184 3800
rect 433248 3748 433300 3800
rect 82636 3680 82688 3732
rect 115296 3680 115348 3732
rect 115940 3680 115992 3732
rect 117228 3680 117280 3732
rect 124220 3680 124272 3732
rect 125508 3680 125560 3732
rect 137284 3680 137336 3732
rect 176476 3680 176528 3732
rect 204260 3680 204312 3732
rect 364248 3680 364300 3732
rect 369216 3680 369268 3732
rect 389088 3680 389140 3732
rect 399024 3680 399076 3732
rect 400128 3680 400180 3732
rect 413284 3680 413336 3732
rect 413928 3680 413980 3732
rect 429936 3680 429988 3732
rect 445668 3748 445720 3800
rect 453856 3748 453908 3800
rect 471888 3748 471940 3800
rect 485688 3748 485740 3800
rect 516784 3748 516836 3800
rect 521568 3748 521620 3800
rect 560760 3748 560812 3800
rect 447048 3680 447100 3732
rect 55312 3612 55364 3664
rect 64696 3612 64748 3664
rect 67824 3544 67876 3596
rect 108304 3612 108356 3664
rect 109960 3612 110012 3664
rect 149152 3612 149204 3664
rect 151544 3612 151596 3664
rect 183560 3612 183612 3664
rect 187240 3612 187292 3664
rect 212724 3612 212776 3664
rect 362868 3612 362920 3664
rect 368020 3612 368072 3664
rect 387708 3612 387760 3664
rect 397828 3612 397880 3664
rect 402796 3612 402848 3664
rect 415676 3612 415728 3664
rect 416596 3612 416648 3664
rect 433524 3612 433576 3664
rect 438768 3612 438820 3664
rect 456064 3612 456116 3664
rect 71780 3544 71832 3596
rect 73804 3544 73856 3596
rect 77300 3544 77352 3596
rect 77944 3544 77996 3596
rect 79048 3544 79100 3596
rect 79968 3544 80020 3596
rect 81440 3544 81492 3596
rect 82728 3544 82780 3596
rect 117964 3544 118016 3596
rect 125416 3544 125468 3596
rect 158720 3544 158772 3596
rect 159916 3544 159968 3596
rect 169392 3544 169444 3596
rect 4068 3476 4120 3528
rect 60004 3476 60056 3528
rect 60648 3476 60700 3528
rect 61200 3476 61252 3528
rect 68284 3476 68336 3528
rect 126612 3476 126664 3528
rect 162952 3476 163004 3528
rect 163504 3476 163556 3528
rect 164148 3476 164200 3528
rect 164700 3476 164752 3528
rect 165528 3476 165580 3528
rect 165896 3476 165948 3528
rect 196072 3544 196124 3596
rect 218152 3544 218204 3596
rect 219348 3544 219400 3596
rect 252652 3544 252704 3596
rect 253848 3544 253900 3596
rect 270500 3544 270552 3596
rect 271696 3544 271748 3596
rect 278872 3544 278924 3596
rect 280068 3544 280120 3596
rect 287152 3544 287204 3596
rect 288348 3544 288400 3596
rect 296720 3544 296772 3596
rect 297916 3544 297968 3596
rect 305000 3544 305052 3596
rect 306196 3544 306248 3596
rect 348976 3544 349028 3596
rect 351368 3544 351420 3596
rect 351736 3544 351788 3596
rect 354956 3544 355008 3596
rect 358728 3544 358780 3596
rect 363328 3544 363380 3596
rect 373908 3544 373960 3596
rect 381176 3544 381228 3596
rect 382096 3544 382148 3596
rect 390652 3544 390704 3596
rect 395988 3544 396040 3596
rect 408500 3544 408552 3596
rect 409788 3544 409840 3596
rect 425152 3544 425204 3596
rect 426348 3544 426400 3596
rect 445392 3544 445444 3596
rect 450176 3544 450228 3596
rect 451188 3544 451240 3596
rect 459468 3680 459520 3732
rect 484584 3680 484636 3732
rect 488448 3680 488500 3732
rect 520280 3680 520332 3732
rect 524236 3680 524288 3732
rect 571432 3680 571484 3732
rect 456340 3612 456392 3664
rect 459652 3612 459704 3664
rect 460848 3612 460900 3664
rect 485780 3612 485832 3664
rect 491208 3612 491260 3664
rect 523868 3612 523920 3664
rect 532608 3612 532660 3664
rect 573824 3612 573876 3664
rect 470324 3544 470376 3596
rect 470508 3544 470560 3596
rect 498936 3544 498988 3596
rect 500868 3544 500920 3596
rect 215852 3476 215904 3528
rect 216588 3476 216640 3528
rect 217048 3476 217100 3528
rect 217968 3476 218020 3528
rect 222936 3476 222988 3528
rect 223488 3476 223540 3528
rect 225328 3476 225380 3528
rect 226248 3476 226300 3528
rect 226524 3476 226576 3528
rect 227628 3476 227680 3528
rect 231308 3476 231360 3528
rect 231768 3476 231820 3528
rect 232504 3476 232556 3528
rect 233148 3476 233200 3528
rect 233700 3476 233752 3528
rect 234528 3476 234580 3528
rect 239588 3476 239640 3528
rect 240048 3476 240100 3528
rect 240784 3476 240836 3528
rect 241428 3476 241480 3528
rect 243176 3476 243228 3528
rect 244188 3476 244240 3528
rect 244372 3476 244424 3528
rect 245476 3476 245528 3528
rect 249156 3476 249208 3528
rect 249708 3476 249760 3528
rect 250352 3476 250404 3528
rect 251088 3476 251140 3528
rect 251456 3476 251508 3528
rect 252468 3476 252520 3528
rect 257436 3476 257488 3528
rect 257988 3476 258040 3528
rect 259828 3476 259880 3528
rect 260748 3476 260800 3528
rect 262220 3476 262272 3528
rect 263508 3476 263560 3528
rect 265808 3476 265860 3528
rect 266268 3476 266320 3528
rect 269304 3476 269356 3528
rect 270408 3476 270460 3528
rect 274088 3476 274140 3528
rect 274548 3476 274600 3528
rect 275284 3476 275336 3528
rect 275928 3476 275980 3528
rect 276480 3476 276532 3528
rect 277308 3476 277360 3528
rect 277676 3476 277728 3528
rect 278688 3476 278740 3528
rect 283656 3476 283708 3528
rect 284208 3476 284260 3528
rect 284760 3476 284812 3528
rect 285588 3476 285640 3528
rect 285956 3476 286008 3528
rect 286968 3476 287020 3528
rect 291936 3476 291988 3528
rect 292488 3476 292540 3528
rect 293132 3476 293184 3528
rect 293868 3476 293920 3528
rect 294328 3476 294380 3528
rect 295248 3476 295300 3528
rect 295524 3476 295576 3528
rect 296628 3476 296680 3528
rect 301412 3476 301464 3528
rect 302148 3476 302200 3528
rect 302608 3476 302660 3528
rect 303528 3476 303580 3528
rect 303804 3476 303856 3528
rect 304908 3476 304960 3528
rect 308588 3476 308640 3528
rect 309048 3476 309100 3528
rect 309784 3476 309836 3528
rect 310428 3476 310480 3528
rect 310980 3476 311032 3528
rect 311808 3476 311860 3528
rect 312176 3476 312228 3528
rect 313188 3476 313240 3528
rect 314568 3476 314620 3528
rect 315304 3476 315356 3528
rect 318064 3476 318116 3528
rect 319444 3476 319496 3528
rect 320456 3476 320508 3528
rect 321468 3476 321520 3528
rect 321652 3476 321704 3528
rect 322756 3476 322808 3528
rect 326436 3476 326488 3528
rect 326988 3476 327040 3528
rect 327632 3476 327684 3528
rect 328368 3476 328420 3528
rect 328828 3476 328880 3528
rect 329932 3476 329984 3528
rect 340880 3476 340932 3528
rect 341892 3476 341944 3528
rect 342168 3476 342220 3528
rect 343088 3476 343140 3528
rect 349068 3476 349120 3528
rect 350264 3476 350316 3528
rect 367008 3476 367060 3528
rect 372804 3476 372856 3528
rect 376668 3476 376720 3528
rect 384672 3476 384724 3528
rect 386236 3476 386288 3528
rect 396632 3476 396684 3528
rect 402888 3476 402940 3528
rect 416872 3476 416924 3528
rect 419356 3476 419408 3528
rect 437020 3476 437072 3528
rect 440056 3476 440108 3528
rect 463240 3476 463292 3528
rect 463608 3476 463660 3528
rect 6460 3408 6512 3460
rect 65064 3408 65116 3460
rect 71872 3408 71924 3460
rect 115204 3408 115256 3460
rect 117136 3408 117188 3460
rect 29092 3340 29144 3392
rect 30196 3340 30248 3392
rect 26700 3204 26752 3256
rect 77760 3340 77812 3392
rect 77852 3340 77904 3392
rect 84936 3340 84988 3392
rect 85488 3340 85540 3392
rect 86132 3340 86184 3392
rect 86868 3340 86920 3392
rect 88524 3340 88576 3392
rect 89628 3340 89680 3392
rect 109684 3340 109736 3392
rect 114744 3340 114796 3392
rect 145564 3340 145616 3392
rect 146852 3340 146904 3392
rect 147588 3340 147640 3392
rect 36176 3272 36228 3324
rect 37188 3272 37240 3324
rect 37372 3272 37424 3324
rect 38476 3272 38528 3324
rect 43352 3272 43404 3324
rect 44088 3272 44140 3324
rect 42156 3204 42208 3256
rect 45744 3272 45796 3324
rect 46848 3272 46900 3324
rect 50528 3272 50580 3324
rect 50988 3272 51040 3324
rect 52828 3272 52880 3324
rect 53748 3272 53800 3324
rect 44548 3204 44600 3256
rect 45468 3204 45520 3256
rect 49332 3204 49384 3256
rect 98644 3272 98696 3324
rect 107660 3272 107712 3324
rect 135904 3272 135956 3324
rect 152464 3408 152516 3460
rect 156328 3408 156380 3460
rect 157248 3408 157300 3460
rect 157524 3408 157576 3460
rect 158628 3408 158680 3460
rect 162308 3408 162360 3460
rect 192300 3408 192352 3460
rect 194416 3408 194468 3460
rect 219532 3408 219584 3460
rect 227720 3408 227772 3460
rect 229008 3408 229060 3460
rect 241980 3408 242032 3460
rect 242808 3408 242860 3460
rect 267004 3408 267056 3460
rect 267648 3408 267700 3460
rect 319260 3408 319312 3460
rect 320088 3408 320140 3460
rect 346216 3408 346268 3460
rect 347872 3408 347924 3460
rect 355968 3408 356020 3460
rect 359740 3408 359792 3460
rect 372528 3408 372580 3460
rect 379980 3408 380032 3460
rect 380164 3408 380216 3460
rect 388260 3408 388312 3460
rect 388996 3408 389048 3460
rect 400220 3408 400272 3460
rect 408408 3408 408460 3460
rect 422760 3408 422812 3460
rect 423588 3408 423640 3460
rect 441804 3408 441856 3460
rect 442816 3408 442868 3460
rect 465632 3408 465684 3460
rect 471520 3476 471572 3528
rect 466368 3408 466420 3460
rect 492956 3476 493008 3528
rect 493968 3476 494020 3528
rect 527456 3476 527508 3528
rect 529204 3544 529256 3596
rect 532240 3544 532292 3596
rect 534540 3476 534592 3528
rect 535368 3544 535420 3596
rect 576216 3544 576268 3596
rect 500132 3408 500184 3460
rect 500776 3408 500828 3460
rect 535736 3408 535788 3460
rect 536748 3476 536800 3528
rect 578608 3476 578660 3528
rect 538036 3408 538088 3460
rect 538128 3408 538180 3460
rect 579804 3408 579856 3460
rect 150440 3340 150492 3392
rect 164884 3340 164936 3392
rect 174176 3340 174228 3392
rect 175188 3340 175240 3392
rect 175372 3340 175424 3392
rect 176568 3340 176620 3392
rect 181352 3340 181404 3392
rect 182088 3340 182140 3392
rect 182548 3340 182600 3392
rect 183468 3340 183520 3392
rect 192024 3340 192076 3392
rect 193128 3340 193180 3392
rect 200396 3340 200448 3392
rect 201408 3340 201460 3392
rect 325240 3340 325292 3392
rect 326344 3340 326396 3392
rect 375288 3340 375340 3392
rect 382372 3340 382424 3392
rect 391848 3340 391900 3392
rect 402520 3340 402572 3392
rect 405648 3340 405700 3392
rect 419172 3340 419224 3392
rect 419448 3340 419500 3392
rect 435824 3340 435876 3392
rect 437388 3340 437440 3392
rect 457260 3340 457312 3392
rect 481088 3340 481140 3392
rect 482928 3340 482980 3392
rect 513196 3340 513248 3392
rect 517428 3340 517480 3392
rect 549904 3340 549956 3392
rect 553584 3340 553636 3392
rect 153844 3272 153896 3324
rect 172704 3272 172756 3324
rect 234804 3272 234856 3324
rect 235908 3272 235960 3324
rect 300308 3272 300360 3324
rect 304264 3272 304316 3324
rect 330024 3272 330076 3324
rect 331128 3272 331180 3324
rect 334072 3272 334124 3324
rect 334716 3272 334768 3324
rect 358636 3272 358688 3324
rect 362132 3272 362184 3324
rect 365628 3272 365680 3324
rect 371608 3272 371660 3324
rect 374644 3272 374696 3324
rect 378784 3272 378836 3324
rect 398748 3272 398800 3324
rect 410892 3272 410944 3324
rect 416688 3272 416740 3324
rect 432328 3272 432380 3324
rect 433156 3272 433208 3324
rect 452476 3272 452528 3324
rect 455328 3272 455380 3324
rect 475108 3272 475160 3324
rect 54024 3204 54076 3256
rect 102784 3204 102836 3256
rect 106372 3204 106424 3256
rect 107568 3204 107620 3256
rect 56416 3136 56468 3188
rect 102876 3136 102928 3188
rect 103980 3136 104032 3188
rect 128912 3204 128964 3256
rect 236000 3204 236052 3256
rect 237288 3204 237340 3256
rect 261024 3204 261076 3256
rect 262128 3204 262180 3256
rect 376576 3204 376628 3256
rect 383568 3204 383620 3256
rect 394608 3204 394660 3256
rect 406108 3204 406160 3256
rect 406936 3204 406988 3256
rect 420368 3204 420420 3256
rect 424968 3204 425020 3256
rect 443000 3204 443052 3256
rect 444288 3204 444340 3256
rect 466828 3204 466880 3256
rect 167092 3136 167144 3188
rect 168288 3136 168340 3188
rect 355876 3136 355928 3188
rect 358544 3136 358596 3188
rect 378048 3136 378100 3188
rect 385868 3136 385920 3188
rect 411168 3136 411220 3188
rect 426348 3136 426400 3188
rect 427728 3136 427780 3188
rect 446588 3136 446640 3188
rect 452568 3136 452620 3188
rect 27896 3068 27948 3120
rect 70400 3068 70452 3120
rect 71044 3068 71096 3120
rect 99288 3068 99340 3120
rect 119344 3068 119396 3120
rect 189632 3068 189684 3120
rect 190368 3068 190420 3120
rect 206284 3068 206336 3120
rect 206928 3068 206980 3120
rect 258632 3068 258684 3120
rect 259368 3068 259420 3120
rect 368388 3068 368440 3120
rect 374000 3068 374052 3120
rect 426256 3068 426308 3120
rect 444196 3068 444248 3120
rect 446956 3068 447008 3120
rect 448336 3068 448388 3120
rect 448428 3068 448480 3120
rect 478696 3272 478748 3324
rect 480168 3272 480220 3324
rect 509608 3272 509660 3324
rect 518808 3272 518860 3324
rect 557172 3272 557224 3324
rect 477408 3204 477460 3256
rect 506020 3204 506072 3256
rect 521384 3204 521436 3256
rect 559564 3204 559616 3256
rect 469128 3136 469180 3188
rect 474648 3136 474700 3188
rect 503628 3136 503680 3188
rect 506388 3136 506440 3188
rect 541716 3136 541768 3188
rect 541900 3136 541952 3188
rect 467932 3068 467984 3120
rect 496544 3068 496596 3120
rect 509148 3068 509200 3120
rect 545304 3068 545356 3120
rect 545764 3136 545816 3188
rect 546500 3136 546552 3188
rect 547144 3136 547196 3188
rect 550088 3136 550140 3188
rect 582196 3136 582248 3188
rect 39764 3000 39816 3052
rect 82084 3000 82136 3052
rect 170588 3000 170640 3052
rect 171048 3000 171100 3052
rect 171784 3000 171836 3052
rect 172428 3000 172480 3052
rect 188436 3000 188488 3052
rect 188988 3000 189040 3052
rect 224132 3000 224184 3052
rect 224868 3000 224920 3052
rect 268108 3000 268160 3052
rect 269028 3000 269080 3052
rect 351828 3000 351880 3052
rect 353760 3000 353812 3052
rect 422208 3000 422260 3052
rect 439412 3000 439464 3052
rect 440148 3000 440200 3052
rect 451188 3000 451240 3052
rect 469128 3000 469180 3052
rect 24308 2932 24360 2984
rect 70400 2932 70452 2984
rect 70676 2932 70728 2984
rect 105544 2932 105596 2984
rect 139676 2932 139728 2984
rect 140688 2932 140740 2984
rect 198004 2932 198056 2984
rect 198648 2932 198700 2984
rect 209872 2932 209924 2984
rect 210976 2932 211028 2984
rect 420828 2932 420880 2984
rect 438216 2932 438268 2984
rect 442908 2932 442960 2984
rect 464436 2932 464488 2984
rect 467748 2932 467800 2984
rect 495348 3000 495400 3052
rect 509884 3000 509936 3052
rect 511908 3000 511960 3052
rect 548892 3000 548944 3052
rect 555976 3000 556028 3052
rect 489368 2932 489420 2984
rect 498108 2932 498160 2984
rect 531044 2932 531096 2984
rect 533344 2932 533396 2984
rect 32680 2864 32732 2916
rect 77300 2864 77352 2916
rect 102784 2864 102836 2916
rect 122104 2864 122156 2916
rect 369676 2864 369728 2916
rect 375196 2864 375248 2916
rect 436008 2864 436060 2916
rect 456064 2864 456116 2916
rect 479892 2864 479944 2916
rect 491944 2864 491996 2916
rect 517888 2864 517940 2916
rect 537484 2864 537536 2916
rect 544384 2932 544436 2984
rect 575020 2932 575072 2984
rect 46940 2796 46992 2848
rect 91744 2796 91796 2848
rect 143448 2796 143500 2848
rect 213828 2796 213880 2848
rect 333888 2796 333940 2848
rect 452660 2796 452712 2848
rect 453672 2796 453724 2848
rect 460756 2796 460808 2848
rect 477500 2796 477552 2848
rect 489184 2796 489236 2848
rect 510804 2796 510856 2848
rect 539324 2796 539376 2848
rect 566740 2864 566792 2916
rect 570236 2796 570288 2848
rect 5264 552 5316 604
rect 5448 552 5500 604
rect 14832 552 14884 604
rect 15108 552 15160 604
rect 143264 595 143316 604
rect 143264 561 143273 595
rect 143273 561 143307 595
rect 143307 561 143316 595
rect 143264 552 143316 561
rect 195612 595 195664 604
rect 195612 561 195621 595
rect 195621 561 195655 595
rect 195655 561 195664 595
rect 195612 552 195664 561
rect 203708 552 203760 604
rect 203892 552 203944 604
rect 212264 552 212316 604
rect 213460 595 213512 604
rect 213460 561 213469 595
rect 213469 561 213503 595
rect 213503 561 213512 595
rect 213460 552 213512 561
rect 316960 552 317012 604
rect 317328 552 317380 604
rect 333612 595 333664 604
rect 333612 561 333621 595
rect 333621 561 333655 595
rect 333655 561 333664 595
rect 333612 552 333664 561
rect 369952 552 370004 604
rect 370412 552 370464 604
rect 485964 552 486016 604
rect 486976 552 487028 604
rect 501052 552 501104 604
rect 501236 552 501288 604
rect 503720 552 503772 604
rect 504824 552 504876 604
rect 507952 552 508004 604
rect 508412 552 508464 604
rect 514760 552 514812 604
rect 515588 552 515640 604
rect 521660 552 521712 604
rect 522672 552 522724 604
rect 525800 552 525852 604
rect 526260 552 526312 604
rect 542360 552 542412 604
rect 542912 552 542964 604
rect 543740 552 543792 604
rect 544108 552 544160 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700369 8156 703520
rect 8114 700360 8170 700369
rect 24320 700330 24348 703520
rect 40512 700398 40540 703520
rect 72988 700602 73016 703520
rect 89180 700670 89208 703520
rect 105464 700738 105492 703520
rect 137848 700942 137876 703520
rect 154132 701010 154160 703520
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 137836 700936 137888 700942
rect 137836 700878 137888 700884
rect 105452 700732 105504 700738
rect 105452 700674 105504 700680
rect 89168 700664 89220 700670
rect 89168 700606 89220 700612
rect 72976 700596 73028 700602
rect 72976 700538 73028 700544
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 8114 700295 8170 700304
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 202800 700058 202828 703520
rect 202788 700052 202840 700058
rect 202788 699994 202840 700000
rect 218992 699990 219020 703520
rect 218980 699984 219032 699990
rect 218980 699926 219032 699932
rect 235184 699718 235212 703520
rect 255228 700528 255280 700534
rect 255228 700470 255280 700476
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 235920 663270 235948 699654
rect 242808 696992 242860 696998
rect 242808 696934 242860 696940
rect 238668 673532 238720 673538
rect 238668 673474 238720 673480
rect 235908 663264 235960 663270
rect 235908 663206 235960 663212
rect 204628 662788 204680 662794
rect 204628 662730 204680 662736
rect 192024 662720 192076 662726
rect 192024 662662 192076 662668
rect 8852 662652 8904 662658
rect 8852 662594 8904 662600
rect 3974 661872 4030 661881
rect 3974 661807 4030 661816
rect 3790 661736 3846 661745
rect 3790 661671 3846 661680
rect 3606 661328 3662 661337
rect 3606 661263 3662 661272
rect 3422 661056 3478 661065
rect 3422 660991 3478 661000
rect 3332 659660 3384 659666
rect 3332 659602 3384 659608
rect 3240 659592 3292 659598
rect 3240 659534 3292 659540
rect 3148 653608 3200 653614
rect 3146 653576 3148 653585
rect 3200 653576 3202 653585
rect 3146 653511 3202 653520
rect 3148 624912 3200 624918
rect 3146 624880 3148 624889
rect 3200 624880 3202 624889
rect 3146 624815 3202 624824
rect 2780 610496 2832 610502
rect 2778 610464 2780 610473
rect 2832 610464 2834 610473
rect 2778 610399 2834 610408
rect 3148 596080 3200 596086
rect 3146 596048 3148 596057
rect 3200 596048 3202 596057
rect 3146 595983 3202 595992
rect 3148 567588 3200 567594
rect 3148 567530 3200 567536
rect 3160 567361 3188 567530
rect 3146 567352 3202 567361
rect 3146 567287 3202 567296
rect 3252 553081 3280 659534
rect 3238 553072 3294 553081
rect 3238 553007 3294 553016
rect 3240 538824 3292 538830
rect 3240 538766 3292 538772
rect 3252 538665 3280 538766
rect 3238 538656 3294 538665
rect 3238 538591 3294 538600
rect 3240 510060 3292 510066
rect 3240 510002 3292 510008
rect 3252 509969 3280 510002
rect 3238 509960 3294 509969
rect 3238 509895 3294 509904
rect 2780 496732 2832 496738
rect 2780 496674 2832 496680
rect 2792 495553 2820 496674
rect 2778 495544 2834 495553
rect 2778 495479 2834 495488
rect 3240 481228 3292 481234
rect 3240 481170 3292 481176
rect 3252 481137 3280 481170
rect 3238 481128 3294 481137
rect 3238 481063 3294 481072
rect 3240 452464 3292 452470
rect 3238 452432 3240 452441
rect 3292 452432 3294 452441
rect 3238 452367 3294 452376
rect 2780 438796 2832 438802
rect 2780 438738 2832 438744
rect 2792 438025 2820 438738
rect 2778 438016 2834 438025
rect 2778 437951 2834 437960
rect 3344 423745 3372 659602
rect 3330 423736 3386 423745
rect 3330 423671 3386 423680
rect 3332 395276 3384 395282
rect 3332 395218 3384 395224
rect 3344 395049 3372 395218
rect 3330 395040 3386 395049
rect 3330 394975 3386 394984
rect 3148 366716 3200 366722
rect 3148 366658 3200 366664
rect 3160 366217 3188 366658
rect 3146 366208 3202 366217
rect 3146 366143 3202 366152
rect 3332 337544 3384 337550
rect 3330 337512 3332 337521
rect 3384 337512 3386 337521
rect 3330 337447 3386 337456
rect 3056 309120 3108 309126
rect 3056 309062 3108 309068
rect 3068 308825 3096 309062
rect 3054 308816 3110 308825
rect 3054 308751 3110 308760
rect 3148 294840 3200 294846
rect 3148 294782 3200 294788
rect 3160 294409 3188 294782
rect 3146 294400 3202 294409
rect 3146 294335 3202 294344
rect 3332 280152 3384 280158
rect 3330 280120 3332 280129
rect 3384 280120 3386 280129
rect 3330 280055 3386 280064
rect 3332 266348 3384 266354
rect 3332 266290 3384 266296
rect 3344 265713 3372 266290
rect 3330 265704 3386 265713
rect 3330 265639 3386 265648
rect 3332 252272 3384 252278
rect 3332 252214 3384 252220
rect 3344 251297 3372 252214
rect 3330 251288 3386 251297
rect 3330 251223 3386 251232
rect 3332 237380 3384 237386
rect 3332 237322 3384 237328
rect 3344 237017 3372 237322
rect 3330 237008 3386 237017
rect 3330 236943 3386 236952
rect 3332 223100 3384 223106
rect 3332 223042 3384 223048
rect 3344 222601 3372 223042
rect 3330 222592 3386 222601
rect 3330 222527 3386 222536
rect 3332 208208 3384 208214
rect 3330 208176 3332 208185
rect 3384 208176 3386 208185
rect 3330 208111 3386 208120
rect 3332 194540 3384 194546
rect 3332 194482 3384 194488
rect 3344 193905 3372 194482
rect 3330 193896 3386 193905
rect 3330 193831 3386 193840
rect 3332 179648 3384 179654
rect 3332 179590 3384 179596
rect 3344 179489 3372 179590
rect 3330 179480 3386 179489
rect 3330 179415 3386 179424
rect 3056 165504 3108 165510
rect 3056 165446 3108 165452
rect 3068 165073 3096 165446
rect 3054 165064 3110 165073
rect 3054 164999 3110 165008
rect 3332 122800 3384 122806
rect 3332 122742 3384 122748
rect 3344 122097 3372 122742
rect 3330 122088 3386 122097
rect 3330 122023 3386 122032
rect 3332 93832 3384 93838
rect 3332 93774 3384 93780
rect 3344 93265 3372 93774
rect 3330 93256 3386 93265
rect 3330 93191 3386 93200
rect 3148 79144 3200 79150
rect 3148 79086 3200 79092
rect 3160 78985 3188 79086
rect 3146 78976 3202 78985
rect 3146 78911 3202 78920
rect 2780 64592 2832 64598
rect 2778 64560 2780 64569
rect 2832 64560 2834 64569
rect 2778 64495 2834 64504
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 2884 21457 2912 22034
rect 2870 21448 2926 21457
rect 2870 21383 2926 21392
rect 3436 7177 3464 660991
rect 3514 659016 3570 659025
rect 3514 658951 3570 658960
rect 3528 35873 3556 658951
rect 3620 50153 3648 661263
rect 3698 658880 3754 658889
rect 3698 658815 3754 658824
rect 3712 136377 3740 658815
rect 3698 136368 3754 136377
rect 3698 136303 3754 136312
rect 3804 107681 3832 661671
rect 3884 661020 3936 661026
rect 3884 660962 3936 660968
rect 3896 323105 3924 660962
rect 3882 323096 3938 323105
rect 3882 323031 3938 323040
rect 3988 150793 4016 661807
rect 4068 661292 4120 661298
rect 4068 661234 4120 661240
rect 4080 380633 4108 661234
rect 4802 661192 4858 661201
rect 4802 661127 4858 661136
rect 4066 380624 4122 380633
rect 4066 380559 4122 380568
rect 3974 150784 4030 150793
rect 3974 150719 4030 150728
rect 3790 107672 3846 107681
rect 3790 107607 3846 107616
rect 4816 64598 4844 661127
rect 8208 660748 8260 660754
rect 8208 660690 8260 660696
rect 8116 660680 8168 660686
rect 8116 660622 8168 660628
rect 8024 660544 8076 660550
rect 8024 660486 8076 660492
rect 7932 660476 7984 660482
rect 7932 660418 7984 660424
rect 7840 660136 7892 660142
rect 7840 660078 7892 660084
rect 7748 660068 7800 660074
rect 7748 660010 7800 660016
rect 7656 659932 7708 659938
rect 7656 659874 7708 659880
rect 7564 659864 7616 659870
rect 7564 659806 7616 659812
rect 6184 659728 6236 659734
rect 6184 659670 6236 659676
rect 5080 659048 5132 659054
rect 5080 658990 5132 658996
rect 4988 658912 5040 658918
rect 4988 658854 5040 658860
rect 4896 658708 4948 658714
rect 4896 658650 4948 658656
rect 4908 438802 4936 658650
rect 5000 496738 5028 658854
rect 5092 610502 5120 658990
rect 5080 610496 5132 610502
rect 5080 610438 5132 610444
rect 4988 496732 5040 496738
rect 4988 496674 5040 496680
rect 4896 438796 4948 438802
rect 4896 438738 4948 438744
rect 6196 165510 6224 659670
rect 7576 252278 7604 659806
rect 7668 294846 7696 659874
rect 7760 337550 7788 660010
rect 7852 395282 7880 660078
rect 7944 452470 7972 660418
rect 8036 510066 8064 660486
rect 8128 567594 8156 660622
rect 8220 624918 8248 660690
rect 8668 659184 8720 659190
rect 8668 659126 8720 659132
rect 8680 653614 8708 659126
rect 8760 659116 8812 659122
rect 8760 659058 8812 659064
rect 8668 653608 8720 653614
rect 8668 653550 8720 653556
rect 8208 624912 8260 624918
rect 8208 624854 8260 624860
rect 8772 596086 8800 659058
rect 8760 596080 8812 596086
rect 8760 596022 8812 596028
rect 8116 567588 8168 567594
rect 8116 567530 8168 567536
rect 8864 538830 8892 662594
rect 9588 662584 9640 662590
rect 9588 662526 9640 662532
rect 9496 662448 9548 662454
rect 9496 662390 9548 662396
rect 9034 662008 9090 662017
rect 9034 661943 9090 661952
rect 8942 658336 8998 658345
rect 8942 658271 8998 658280
rect 8852 538824 8904 538830
rect 8852 538766 8904 538772
rect 8024 510060 8076 510066
rect 8024 510002 8076 510008
rect 7932 452464 7984 452470
rect 7932 452406 7984 452412
rect 7840 395276 7892 395282
rect 7840 395218 7892 395224
rect 7748 337544 7800 337550
rect 7748 337486 7800 337492
rect 7656 294840 7708 294846
rect 7656 294782 7708 294788
rect 7564 252272 7616 252278
rect 7564 252214 7616 252220
rect 6184 165504 6236 165510
rect 6184 165446 6236 165452
rect 8956 79150 8984 658271
rect 9048 179654 9076 661943
rect 9404 661156 9456 661162
rect 9404 661098 9456 661104
rect 9128 661088 9180 661094
rect 9128 661030 9180 661036
rect 9140 194546 9168 661030
rect 9220 659796 9272 659802
rect 9220 659738 9272 659744
rect 9232 208214 9260 659738
rect 9312 658572 9364 658578
rect 9312 658514 9364 658520
rect 9324 223106 9352 658514
rect 9416 280158 9444 661098
rect 9508 366722 9536 662390
rect 9600 481234 9628 662526
rect 175188 662516 175240 662522
rect 175188 662458 175240 662464
rect 95240 662380 95292 662386
rect 95240 662322 95292 662328
rect 58622 662144 58678 662153
rect 58622 662079 58678 662088
rect 53104 661564 53156 661570
rect 53104 661506 53156 661512
rect 25502 659832 25558 659841
rect 25502 659767 25558 659776
rect 9588 481228 9640 481234
rect 9588 481170 9640 481176
rect 9496 366716 9548 366722
rect 9496 366658 9548 366664
rect 9404 280152 9456 280158
rect 9404 280094 9456 280100
rect 9312 223100 9364 223106
rect 9312 223042 9364 223048
rect 9220 208208 9272 208214
rect 9220 208150 9272 208156
rect 9128 194540 9180 194546
rect 9128 194482 9180 194488
rect 9036 179648 9088 179654
rect 9036 179590 9088 179596
rect 25516 122806 25544 659767
rect 53116 309126 53144 661506
rect 54484 661360 54536 661366
rect 54484 661302 54536 661308
rect 53104 309120 53156 309126
rect 53104 309062 53156 309068
rect 54496 266354 54524 661302
rect 54484 266348 54536 266354
rect 54484 266290 54536 266296
rect 25504 122800 25556 122806
rect 25504 122742 25556 122748
rect 58636 93838 58664 662079
rect 91008 661904 91060 661910
rect 91008 661846 91060 661852
rect 82544 661632 82596 661638
rect 69938 661600 69994 661609
rect 82544 661574 82596 661580
rect 69938 661535 69994 661544
rect 65706 661464 65762 661473
rect 65706 661399 65762 661408
rect 58716 660204 58768 660210
rect 58716 660146 58768 660152
rect 58728 237386 58756 660146
rect 65720 659940 65748 661399
rect 69952 659940 69980 661535
rect 74354 659968 74410 659977
rect 74198 659926 74354 659954
rect 82556 659940 82584 661574
rect 86774 660104 86830 660113
rect 86774 660039 86830 660048
rect 86788 659940 86816 660039
rect 91020 659940 91048 661846
rect 95252 659940 95280 662322
rect 112076 662108 112128 662114
rect 112076 662050 112128 662056
rect 107844 661972 107896 661978
rect 107844 661914 107896 661920
rect 103612 661224 103664 661230
rect 103612 661166 103664 661172
rect 99656 660000 99708 660006
rect 99406 659948 99656 659954
rect 99406 659942 99708 659948
rect 99406 659926 99696 659942
rect 103624 659940 103652 661166
rect 107856 659940 107884 661914
rect 112088 659940 112116 662050
rect 169760 661972 169812 661978
rect 169760 661914 169812 661920
rect 165896 661904 165948 661910
rect 165896 661846 165948 661852
rect 120448 661768 120500 661774
rect 120448 661710 120500 661716
rect 158720 661768 158772 661774
rect 158720 661710 158772 661716
rect 162584 661768 162636 661774
rect 162584 661710 162636 661716
rect 120460 659940 120488 661710
rect 154120 661700 154172 661706
rect 154120 661642 154172 661648
rect 145748 661496 145800 661502
rect 145748 661438 145800 661444
rect 141516 661428 141568 661434
rect 141516 661370 141568 661376
rect 133052 660272 133104 660278
rect 133052 660214 133104 660220
rect 133064 659940 133092 660214
rect 141528 659940 141556 661370
rect 145760 659940 145788 661438
rect 149980 660612 150032 660618
rect 149980 660554 150032 660560
rect 149992 659940 150020 660554
rect 154132 659940 154160 661642
rect 155684 661632 155736 661638
rect 155684 661574 155736 661580
rect 158352 661632 158404 661638
rect 158352 661574 158404 661580
rect 74354 659903 74410 659912
rect 61934 659696 61990 659705
rect 61594 659654 61934 659682
rect 61934 659631 61990 659640
rect 155696 659433 155724 661574
rect 158364 659940 158392 661574
rect 158732 660346 158760 661710
rect 158720 660340 158772 660346
rect 158720 660282 158772 660288
rect 162596 659940 162624 661710
rect 78586 659424 78642 659433
rect 78430 659382 78586 659410
rect 78586 659359 78642 659368
rect 155682 659424 155738 659433
rect 155682 659359 155738 659368
rect 165908 659326 165936 661846
rect 166816 661836 166868 661842
rect 166816 661778 166868 661784
rect 166828 659940 166856 661778
rect 169772 660414 169800 661914
rect 170956 661904 171008 661910
rect 170956 661846 171008 661852
rect 169760 660408 169812 660414
rect 169760 660350 169812 660356
rect 170968 659940 170996 661846
rect 175200 659940 175228 662458
rect 183652 661972 183704 661978
rect 183652 661914 183704 661920
rect 183664 659940 183692 661914
rect 187792 660816 187844 660822
rect 187792 660758 187844 660764
rect 187804 659940 187832 660758
rect 192036 659940 192064 662662
rect 196256 662040 196308 662046
rect 196256 661982 196308 661988
rect 196268 659940 196296 661982
rect 200488 660884 200540 660890
rect 200488 660826 200540 660832
rect 200500 659940 200528 660826
rect 204640 659940 204668 662730
rect 232596 662380 232648 662386
rect 232596 662322 232648 662328
rect 233884 662380 233936 662386
rect 233884 662322 233936 662328
rect 208860 662312 208912 662318
rect 208860 662254 208912 662260
rect 208872 659940 208900 662254
rect 230664 662244 230716 662250
rect 230664 662186 230716 662192
rect 213828 662176 213880 662182
rect 213828 662118 213880 662124
rect 213840 661026 213868 662118
rect 213828 661020 213880 661026
rect 213828 660962 213880 660968
rect 225696 661020 225748 661026
rect 225696 660962 225748 660968
rect 213092 660952 213144 660958
rect 213092 660894 213144 660900
rect 213104 659940 213132 660894
rect 225708 659940 225736 660962
rect 230676 659666 230704 662186
rect 232608 660249 232636 662322
rect 232594 660240 232650 660249
rect 232594 660175 232650 660184
rect 230664 659660 230716 659666
rect 230664 659602 230716 659608
rect 233896 659598 233924 662322
rect 238680 659954 238708 673474
rect 242820 659954 242848 696934
rect 246948 685908 247000 685914
rect 246948 685850 247000 685856
rect 246960 659954 246988 685850
rect 250996 663060 251048 663066
rect 250996 663002 251048 663008
rect 238418 659926 238708 659954
rect 242558 659926 242848 659954
rect 246790 659926 246988 659954
rect 251008 659940 251036 663002
rect 255240 659940 255268 700470
rect 259368 700460 259420 700466
rect 259368 700402 259420 700408
rect 259380 659940 259408 700402
rect 267660 699854 267688 703520
rect 269028 700868 269080 700874
rect 269028 700810 269080 700816
rect 267648 699848 267700 699854
rect 267648 699790 267700 699796
rect 263600 663128 263652 663134
rect 263600 663070 263652 663076
rect 263612 659940 263640 663070
rect 269040 660090 269068 700810
rect 273168 700800 273220 700806
rect 273168 700742 273220 700748
rect 273180 660090 273208 700742
rect 281448 700120 281500 700126
rect 281448 700062 281500 700068
rect 276204 663196 276256 663202
rect 276204 663138 276256 663144
rect 268396 660062 269068 660090
rect 272628 660062 273208 660090
rect 268396 659818 268424 660062
rect 272628 659818 272656 660062
rect 276216 659940 276244 663138
rect 281460 660090 281488 700062
rect 283852 699718 283880 703520
rect 285588 700188 285640 700194
rect 285588 700130 285640 700136
rect 283840 699712 283892 699718
rect 283840 699654 283892 699660
rect 280908 660062 281488 660090
rect 280908 659818 280936 660062
rect 285600 659818 285628 700130
rect 300136 699854 300164 703520
rect 329840 700936 329892 700942
rect 329840 700878 329892 700884
rect 325700 700256 325752 700262
rect 325700 700198 325752 700204
rect 317420 700052 317472 700058
rect 317420 699994 317472 700000
rect 298008 699848 298060 699854
rect 298008 699790 298060 699796
rect 300124 699848 300176 699854
rect 300124 699790 300176 699796
rect 300768 699848 300820 699854
rect 300768 699790 300820 699796
rect 293868 699780 293920 699786
rect 293868 699722 293920 699728
rect 288900 663332 288952 663338
rect 288900 663274 288952 663280
rect 288912 659940 288940 663274
rect 293880 659818 293908 699722
rect 298020 659818 298048 699790
rect 300780 662862 300808 699790
rect 309140 699712 309192 699718
rect 309140 699654 309192 699660
rect 305000 699644 305052 699650
rect 305000 699586 305052 699592
rect 300768 662856 300820 662862
rect 300768 662798 300820 662804
rect 301504 662856 301556 662862
rect 301504 662798 301556 662804
rect 301516 659940 301544 662798
rect 305012 660090 305040 699586
rect 305012 660062 305316 660090
rect 267858 659790 268424 659818
rect 272090 659790 272656 659818
rect 280462 659790 280936 659818
rect 284694 659790 285628 659818
rect 293066 659790 293908 659818
rect 297298 659790 298048 659818
rect 305288 659818 305316 660062
rect 309152 659818 309180 699654
rect 314108 663264 314160 663270
rect 314108 663206 314160 663212
rect 314120 659940 314148 663206
rect 317432 659818 317460 699994
rect 321560 699984 321612 699990
rect 321560 699926 321612 699932
rect 321572 660090 321600 699926
rect 325712 660090 325740 700198
rect 329852 660090 329880 700878
rect 332520 699786 332548 703520
rect 333980 701004 334032 701010
rect 333980 700946 334032 700952
rect 332508 699780 332560 699786
rect 332508 699722 332560 699728
rect 333992 660090 334020 700946
rect 338120 700732 338172 700738
rect 338120 700674 338172 700680
rect 338132 660090 338160 700674
rect 347872 700664 347924 700670
rect 347872 700606 347924 700612
rect 343640 700596 343692 700602
rect 343640 700538 343692 700544
rect 321572 660062 322060 660090
rect 325712 660062 326292 660090
rect 329852 660062 330524 660090
rect 333992 660062 334756 660090
rect 338132 660062 338988 660090
rect 322032 659818 322060 660062
rect 326264 659818 326292 660062
rect 330496 659818 330524 660062
rect 334728 659818 334756 660062
rect 338960 659818 338988 660062
rect 343652 659940 343680 700538
rect 347884 659954 347912 700606
rect 348804 699922 348832 703520
rect 364996 703474 365024 703520
rect 364996 703446 365116 703474
rect 351920 700392 351972 700398
rect 351920 700334 351972 700340
rect 356058 700360 356114 700369
rect 348792 699916 348844 699922
rect 348792 699858 348844 699864
rect 347806 659926 347912 659954
rect 351932 659954 351960 700334
rect 356058 700295 356114 700304
rect 360200 700324 360252 700330
rect 356072 659954 356100 700295
rect 360200 700266 360252 700272
rect 360212 659954 360240 700266
rect 365088 692850 365116 703446
rect 397472 700126 397500 703520
rect 413664 700194 413692 703520
rect 413652 700188 413704 700194
rect 413652 700130 413704 700136
rect 397460 700120 397512 700126
rect 397460 700062 397512 700068
rect 364340 692844 364392 692850
rect 364340 692786 364392 692792
rect 365076 692844 365128 692850
rect 365076 692786 365128 692792
rect 364352 683126 364380 692786
rect 429856 688922 429884 703520
rect 462332 700874 462360 703520
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 478524 700806 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 429580 688894 429884 688922
rect 429580 688650 429608 688894
rect 429488 688622 429608 688650
rect 364340 683120 364392 683126
rect 364340 683062 364392 683068
rect 364616 683120 364668 683126
rect 364616 683062 364668 683068
rect 364432 681760 364484 681766
rect 364432 681702 364484 681708
rect 364340 673600 364392 673606
rect 364340 673542 364392 673548
rect 364352 668642 364380 673542
rect 364340 668636 364392 668642
rect 364340 668578 364392 668584
rect 364444 659954 364472 681702
rect 364628 673606 364656 683062
rect 364616 673600 364668 673606
rect 364616 673542 364668 673548
rect 429488 669338 429516 688622
rect 494900 686089 494928 703446
rect 527192 700534 527220 703520
rect 527180 700528 527232 700534
rect 527180 700470 527232 700476
rect 543476 700466 543504 703520
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 559668 688786 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 559300 688758 559696 688786
rect 559300 688650 559328 688758
rect 559208 688622 559328 688650
rect 494886 686080 494942 686089
rect 494886 686015 494942 686024
rect 494242 685944 494298 685953
rect 494242 685879 494298 685888
rect 494256 678994 494284 685879
rect 494072 678966 494284 678994
rect 494072 676190 494100 678966
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 559208 669338 559236 688622
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 580172 685850 580224 685856
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 429304 669310 429516 669338
rect 559024 669310 559236 669338
rect 364524 668636 364576 668642
rect 364524 668578 364576 668584
rect 364536 663338 364564 668578
rect 372620 667956 372672 667962
rect 372620 667898 372672 667904
rect 364524 663332 364576 663338
rect 364524 663274 364576 663280
rect 369124 662108 369176 662114
rect 369124 662050 369176 662056
rect 351932 659926 352038 659954
rect 356072 659926 356270 659954
rect 360212 659926 360502 659954
rect 364444 659926 364642 659954
rect 305288 659790 305762 659818
rect 309152 659790 309994 659818
rect 317432 659790 318366 659818
rect 322032 659790 322598 659818
rect 326264 659790 326830 659818
rect 330496 659790 330970 659818
rect 334728 659790 335202 659818
rect 338960 659790 339434 659818
rect 368584 659666 368874 659682
rect 369136 659666 369164 662050
rect 372632 659818 372660 667898
rect 429304 663202 429332 669310
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 429292 663196 429344 663202
rect 429292 663138 429344 663144
rect 494164 663134 494192 666538
rect 494152 663128 494204 663134
rect 494152 663070 494204 663076
rect 559024 663066 559052 669310
rect 559012 663060 559064 663066
rect 559012 663002 559064 663008
rect 539876 662788 539928 662794
rect 539876 662730 539928 662736
rect 394148 662652 394200 662658
rect 394148 662594 394200 662600
rect 381636 662312 381688 662318
rect 381636 662254 381688 662260
rect 377312 660748 377364 660754
rect 377312 660690 377364 660696
rect 377324 659940 377352 660690
rect 372632 659790 373106 659818
rect 381280 659666 381570 659682
rect 381648 659666 381676 662254
rect 389916 660680 389968 660686
rect 389916 660622 389968 660628
rect 389928 659940 389956 660622
rect 394160 659940 394188 662594
rect 406752 662584 406804 662590
rect 406752 662526 406804 662532
rect 398380 662380 398432 662386
rect 398380 662322 398432 662328
rect 398392 659940 398420 662322
rect 402520 660544 402572 660550
rect 402520 660486 402572 660492
rect 402532 659940 402560 660486
rect 406764 659940 406792 662526
rect 432052 662448 432104 662454
rect 432052 662390 432104 662396
rect 419356 662244 419408 662250
rect 419356 662186 419408 662192
rect 415216 660476 415268 660482
rect 415216 660418 415268 660424
rect 415228 659940 415256 660418
rect 419368 659940 419396 662186
rect 427820 660136 427872 660142
rect 427820 660078 427872 660084
rect 427832 659940 427860 660078
rect 432064 659940 432092 662390
rect 448888 662176 448940 662182
rect 448888 662118 448940 662124
rect 507766 662144 507822 662153
rect 444656 661564 444708 661570
rect 444656 661506 444708 661512
rect 436192 661292 436244 661298
rect 436192 661234 436244 661240
rect 436204 659940 436232 661234
rect 440240 660068 440292 660074
rect 440240 660010 440292 660016
rect 440252 659954 440280 660010
rect 440252 659926 440450 659954
rect 444668 659940 444696 661506
rect 448520 661292 448572 661298
rect 448520 661234 448572 661240
rect 385328 659666 385710 659682
rect 410720 659666 411010 659682
rect 423232 659666 423614 659682
rect 368572 659660 368874 659666
rect 368624 659654 368874 659660
rect 369124 659660 369176 659666
rect 368572 659602 368624 659608
rect 369124 659602 369176 659608
rect 381268 659660 381570 659666
rect 381320 659654 381570 659660
rect 381636 659660 381688 659666
rect 381268 659602 381320 659608
rect 381636 659602 381688 659608
rect 385316 659660 385710 659666
rect 385368 659654 385710 659660
rect 410708 659660 411010 659666
rect 385316 659602 385368 659608
rect 410760 659654 411010 659660
rect 423220 659660 423614 659666
rect 410708 659602 410760 659608
rect 423272 659654 423614 659660
rect 423220 659602 423272 659608
rect 233884 659592 233936 659598
rect 229954 659530 230336 659546
rect 234528 659592 234580 659598
rect 233884 659534 233936 659540
rect 234186 659540 234528 659546
rect 234186 659534 234580 659540
rect 229954 659524 230348 659530
rect 229954 659518 230296 659524
rect 234186 659518 234568 659534
rect 230296 659466 230348 659472
rect 221832 659456 221884 659462
rect 179446 659394 179736 659410
rect 217350 659394 217640 659410
rect 221582 659404 221832 659410
rect 448532 659433 448560 661234
rect 448900 659940 448928 662118
rect 507766 662079 507822 662088
rect 482558 662008 482614 662017
rect 482558 661943 482614 661952
rect 457260 661360 457312 661366
rect 457260 661302 457312 661308
rect 457536 661360 457588 661366
rect 457536 661302 457588 661308
rect 452672 659938 453054 659954
rect 457272 659940 457300 661302
rect 452660 659932 453054 659938
rect 452712 659926 453054 659932
rect 452660 659874 452712 659880
rect 457548 659433 457576 661302
rect 461492 661156 461544 661162
rect 461492 661098 461544 661104
rect 461504 659940 461532 661098
rect 474096 660204 474148 660210
rect 474096 660146 474148 660152
rect 474108 659940 474136 660146
rect 482572 659940 482600 661943
rect 499394 661872 499450 661881
rect 499394 661807 499450 661816
rect 495164 661360 495216 661366
rect 495164 661302 495216 661308
rect 486792 661088 486844 661094
rect 486792 661030 486844 661036
rect 486804 659940 486832 661030
rect 495176 659940 495204 661302
rect 499408 659940 499436 661807
rect 507780 659940 507808 662079
rect 538772 661768 538824 661774
rect 511998 661736 512054 661745
rect 538772 661710 538824 661716
rect 511998 661671 512054 661680
rect 512012 659940 512040 661671
rect 520462 661328 520518 661337
rect 520462 661263 520518 661272
rect 528836 661292 528888 661298
rect 520476 659940 520504 661263
rect 528836 661234 528888 661240
rect 524602 661192 524658 661201
rect 524602 661127 524658 661136
rect 524616 659940 524644 661127
rect 528848 659940 528876 661234
rect 533066 661056 533122 661065
rect 533066 660991 533122 661000
rect 538404 661020 538456 661026
rect 533080 659940 533108 660991
rect 538404 660962 538456 660968
rect 465356 659864 465408 659870
rect 503258 659832 503314 659841
rect 465408 659812 465750 659818
rect 465356 659806 465750 659812
rect 465368 659790 465750 659806
rect 478064 659802 478354 659818
rect 478052 659796 478354 659802
rect 478104 659790 478354 659796
rect 503314 659790 503654 659818
rect 503258 659767 503314 659776
rect 478052 659738 478104 659744
rect 490564 659728 490616 659734
rect 469600 659666 469982 659682
rect 490616 659676 490958 659682
rect 490564 659670 490958 659676
rect 469588 659660 469982 659666
rect 469640 659654 469982 659660
rect 490576 659654 490958 659670
rect 469588 659602 469640 659608
rect 221582 659398 221884 659404
rect 448518 659424 448574 659433
rect 179446 659388 179748 659394
rect 179446 659382 179696 659388
rect 217350 659388 217652 659394
rect 217350 659382 217600 659388
rect 179696 659330 179748 659336
rect 221582 659382 221872 659398
rect 448518 659359 448574 659368
rect 457534 659424 457590 659433
rect 457534 659359 457590 659368
rect 516138 659424 516194 659433
rect 516194 659382 516258 659410
rect 516138 659359 516194 659368
rect 217600 659330 217652 659336
rect 116584 659320 116636 659326
rect 116242 659268 116584 659274
rect 125048 659320 125100 659326
rect 116242 659262 116636 659268
rect 124706 659268 125048 659274
rect 129280 659320 129332 659326
rect 124706 659262 125100 659268
rect 128938 659268 129280 659274
rect 137560 659320 137612 659326
rect 128938 659262 129332 659268
rect 137310 659268 137560 659274
rect 137310 659262 137612 659268
rect 165896 659320 165948 659326
rect 165896 659262 165948 659268
rect 116242 659246 116624 659262
rect 124706 659246 125088 659262
rect 128938 659246 129320 659262
rect 137310 659246 137600 659262
rect 537326 659246 538076 659274
rect 58716 237380 58768 237386
rect 58716 237322 58768 237328
rect 58624 93832 58676 93838
rect 58624 93774 58676 93780
rect 8944 79144 8996 79150
rect 8944 79086 8996 79092
rect 4804 64592 4856 64598
rect 4804 64534 4856 64540
rect 101232 60166 102074 60194
rect 121748 60166 122682 60194
rect 145300 60166 146142 60194
rect 192312 60166 193154 60194
rect 334360 60166 335202 60194
rect 59372 60030 60030 60058
rect 60844 60030 60950 60058
rect 61672 60030 61962 60058
rect 44088 57928 44140 57934
rect 44088 57870 44140 57876
rect 41328 57860 41380 57866
rect 41328 57802 41380 57808
rect 38476 57792 38528 57798
rect 38476 57734 38528 57740
rect 30196 57656 30248 57662
rect 30196 57598 30248 57604
rect 23388 57520 23440 57526
rect 23388 57462 23440 57468
rect 21916 57452 21968 57458
rect 21916 57394 21968 57400
rect 15108 57384 15160 57390
rect 15108 57326 15160 57332
rect 12348 57316 12400 57322
rect 12348 57258 12400 57264
rect 5446 57216 5502 57225
rect 5446 57151 5502 57160
rect 3606 50144 3662 50153
rect 3606 50079 3662 50088
rect 3514 35864 3570 35873
rect 3514 35799 3570 35808
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 572 4888 624 4894
rect 572 4830 624 4836
rect 584 480 612 4830
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 480 1716 4762
rect 2884 480 2912 4966
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4080 480 4108 3470
rect 5460 610 5488 57151
rect 7656 4956 7708 4962
rect 7656 4898 7708 4904
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 5264 604 5316 610
rect 5264 546 5316 552
rect 5448 604 5500 610
rect 5448 546 5500 552
rect 5276 480 5304 546
rect 6472 480 6500 3402
rect 7668 480 7696 4898
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 8864 480 8892 3946
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10060 480 10088 3674
rect 12360 3602 12388 57258
rect 13636 57248 13688 57254
rect 13636 57190 13688 57196
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 11256 480 11284 3538
rect 12452 480 12480 5170
rect 13648 480 13676 57190
rect 15120 610 15148 57326
rect 17224 5092 17276 5098
rect 17224 5034 17276 5040
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 14832 604 14884 610
rect 14832 546 14884 552
rect 15108 604 15160 610
rect 15108 546 15160 552
rect 14844 480 14872 546
rect 16040 480 16068 3878
rect 17236 480 17264 5034
rect 21928 4146 21956 57394
rect 22008 5160 22060 5166
rect 22008 5102 22060 5108
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 21916 4140 21968 4146
rect 21916 4082 21968 4088
rect 19524 3868 19576 3874
rect 19524 3810 19576 3816
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18340 480 18368 3674
rect 19536 480 19564 3810
rect 20732 480 20760 4082
rect 22020 2666 22048 5102
rect 23400 3482 23428 57462
rect 25504 3800 25556 3806
rect 25504 3742 25556 3748
rect 21928 2638 22048 2666
rect 23124 3454 23428 3482
rect 21928 480 21956 2638
rect 23124 480 23152 3454
rect 24308 2984 24360 2990
rect 24308 2926 24360 2932
rect 24320 480 24348 2926
rect 25516 480 25544 3742
rect 30208 3398 30236 57598
rect 31668 57588 31720 57594
rect 31668 57530 31720 57536
rect 30288 5296 30340 5302
rect 30288 5238 30340 5244
rect 29092 3392 29144 3398
rect 29092 3334 29144 3340
rect 30196 3392 30248 3398
rect 30196 3334 30248 3340
rect 26700 3256 26752 3262
rect 26700 3198 26752 3204
rect 26712 480 26740 3198
rect 27896 3120 27948 3126
rect 27896 3062 27948 3068
rect 27908 480 27936 3062
rect 29104 480 29132 3334
rect 30300 480 30328 5238
rect 31680 3482 31708 57530
rect 37188 57180 37240 57186
rect 37188 57122 37240 57128
rect 33876 3936 33928 3942
rect 33876 3878 33928 3884
rect 31496 3454 31708 3482
rect 31496 480 31524 3454
rect 32680 2916 32732 2922
rect 32680 2858 32732 2864
rect 32692 480 32720 2858
rect 33888 480 33916 3878
rect 34980 3868 35032 3874
rect 34980 3810 35032 3816
rect 34992 480 35020 3810
rect 37200 3330 37228 57122
rect 38488 3330 38516 57734
rect 38568 57724 38620 57730
rect 38568 57666 38620 57672
rect 36176 3324 36228 3330
rect 36176 3266 36228 3272
rect 37188 3324 37240 3330
rect 37188 3266 37240 3272
rect 37372 3324 37424 3330
rect 37372 3266 37424 3272
rect 38476 3324 38528 3330
rect 38476 3266 38528 3272
rect 36188 480 36216 3266
rect 37384 480 37412 3266
rect 38580 480 38608 57666
rect 41340 3482 41368 57802
rect 40972 3454 41368 3482
rect 39764 3052 39816 3058
rect 39764 2994 39816 3000
rect 39776 480 39804 2994
rect 40972 480 41000 3454
rect 44100 3330 44128 57870
rect 45468 57112 45520 57118
rect 45468 57054 45520 57060
rect 43352 3324 43404 3330
rect 43352 3266 43404 3272
rect 44088 3324 44140 3330
rect 44088 3266 44140 3272
rect 42156 3256 42208 3262
rect 42156 3198 42208 3204
rect 42168 480 42196 3198
rect 43364 480 43392 3266
rect 45480 3262 45508 57054
rect 50988 57044 51040 57050
rect 50988 56986 51040 56992
rect 46848 56976 46900 56982
rect 46848 56918 46900 56924
rect 46860 3330 46888 56918
rect 48136 5364 48188 5370
rect 48136 5306 48188 5312
rect 45744 3324 45796 3330
rect 45744 3266 45796 3272
rect 46848 3324 46900 3330
rect 46848 3266 46900 3272
rect 44548 3256 44600 3262
rect 44548 3198 44600 3204
rect 45468 3256 45520 3262
rect 45468 3198 45520 3204
rect 44560 480 44588 3198
rect 45756 480 45784 3266
rect 46940 2848 46992 2854
rect 46940 2790 46992 2796
rect 46952 480 46980 2790
rect 48148 480 48176 5306
rect 51000 3330 51028 56986
rect 53748 56840 53800 56846
rect 53748 56782 53800 56788
rect 51632 5500 51684 5506
rect 51632 5442 51684 5448
rect 50528 3324 50580 3330
rect 50528 3266 50580 3272
rect 50988 3324 51040 3330
rect 50988 3266 51040 3272
rect 49332 3256 49384 3262
rect 49332 3198 49384 3204
rect 49344 480 49372 3198
rect 50540 480 50568 3266
rect 51644 480 51672 5442
rect 53760 3330 53788 56782
rect 57888 56772 57940 56778
rect 57888 56714 57940 56720
rect 55220 4752 55272 4758
rect 55220 4694 55272 4700
rect 52828 3324 52880 3330
rect 52828 3266 52880 3272
rect 53748 3324 53800 3330
rect 53748 3266 53800 3272
rect 52840 480 52868 3266
rect 54024 3256 54076 3262
rect 54024 3198 54076 3204
rect 54036 480 54064 3198
rect 55232 480 55260 4694
rect 55312 3664 55364 3670
rect 55310 3632 55312 3641
rect 55364 3632 55366 3641
rect 55310 3567 55366 3576
rect 56416 3188 56468 3194
rect 56416 3130 56468 3136
rect 56428 480 56456 3130
rect 57900 626 57928 56714
rect 58808 5432 58860 5438
rect 58808 5374 58860 5380
rect 57624 598 57928 626
rect 57624 480 57652 598
rect 58820 480 58848 5374
rect 59372 4894 59400 60030
rect 60740 57996 60792 58002
rect 60740 57938 60792 57944
rect 60648 56636 60700 56642
rect 60648 56578 60700 56584
rect 59360 4888 59412 4894
rect 59360 4830 59412 4836
rect 60660 3534 60688 56578
rect 60752 5030 60780 57938
rect 60740 5024 60792 5030
rect 60740 4966 60792 4972
rect 60844 4826 60872 60030
rect 61672 58002 61700 60030
rect 61660 57996 61712 58002
rect 61660 57938 61712 57944
rect 62868 56914 62896 60044
rect 63880 57225 63908 60044
rect 64906 60030 65104 60058
rect 64972 57384 65024 57390
rect 64972 57326 65024 57332
rect 63866 57216 63922 57225
rect 63866 57151 63922 57160
rect 61384 56908 61436 56914
rect 61384 56850 61436 56856
rect 62856 56908 62908 56914
rect 62856 56850 62908 56856
rect 60832 4820 60884 4826
rect 60832 4762 60884 4768
rect 61396 4214 61424 56850
rect 64788 56772 64840 56778
rect 64788 56714 64840 56720
rect 61476 56704 61528 56710
rect 61476 56646 61528 56652
rect 61384 4208 61436 4214
rect 61384 4150 61436 4156
rect 61488 4010 61516 56646
rect 62396 4820 62448 4826
rect 62396 4762 62448 4768
rect 61476 4004 61528 4010
rect 61476 3946 61528 3952
rect 60004 3528 60056 3534
rect 60004 3470 60056 3476
rect 60648 3528 60700 3534
rect 60648 3470 60700 3476
rect 61200 3528 61252 3534
rect 61200 3470 61252 3476
rect 60016 480 60044 3470
rect 61212 480 61240 3470
rect 62408 480 62436 4762
rect 63592 4004 63644 4010
rect 63592 3946 63644 3952
rect 63604 480 63632 3946
rect 64696 3664 64748 3670
rect 64694 3632 64696 3641
rect 64748 3632 64750 3641
rect 64694 3567 64750 3576
rect 64800 480 64828 56714
rect 64984 4962 65012 57326
rect 64972 4956 65024 4962
rect 64972 4898 65024 4904
rect 65076 3466 65104 60030
rect 65536 60030 65826 60058
rect 65536 57390 65564 60030
rect 65524 57384 65576 57390
rect 65524 57326 65576 57332
rect 66824 56710 66852 60044
rect 66812 56704 66864 56710
rect 66812 56646 66864 56652
rect 67548 56704 67600 56710
rect 67548 56646 67600 56652
rect 65984 4888 66036 4894
rect 65984 4830 66036 4836
rect 65064 3460 65116 3466
rect 65064 3402 65116 3408
rect 65996 480 66024 4830
rect 67560 626 67588 56646
rect 67836 3602 67864 60044
rect 68756 57322 68784 60044
rect 69032 60030 69782 60058
rect 68744 57316 68796 57322
rect 68744 57258 68796 57264
rect 69032 5234 69060 60030
rect 70780 57390 70808 60044
rect 70768 57384 70820 57390
rect 70768 57326 70820 57332
rect 71044 57384 71096 57390
rect 71044 57326 71096 57332
rect 69020 5228 69072 5234
rect 69020 5170 69072 5176
rect 69480 5024 69532 5030
rect 69480 4966 69532 4972
rect 67824 3596 67876 3602
rect 67824 3538 67876 3544
rect 68284 3528 68336 3534
rect 68284 3470 68336 3476
rect 67192 598 67588 626
rect 67192 480 67220 598
rect 68296 480 68324 3470
rect 69492 480 69520 4966
rect 71056 3126 71084 57326
rect 71136 57316 71188 57322
rect 71136 57258 71188 57264
rect 71148 4146 71176 57258
rect 71700 57254 71728 60044
rect 71792 60030 72726 60058
rect 73172 60030 73738 60058
rect 71688 57248 71740 57254
rect 71688 57190 71740 57196
rect 71136 4140 71188 4146
rect 71136 4082 71188 4088
rect 71792 3602 71820 60030
rect 73172 5098 73200 60030
rect 74644 57254 74672 60044
rect 75656 57322 75684 60044
rect 76576 57458 76604 60044
rect 77404 60030 77602 60058
rect 76564 57452 76616 57458
rect 76564 57394 76616 57400
rect 75644 57316 75696 57322
rect 75644 57258 75696 57264
rect 75828 57316 75880 57322
rect 75828 57258 75880 57264
rect 73804 57248 73856 57254
rect 73804 57190 73856 57196
rect 74632 57248 74684 57254
rect 74632 57190 74684 57196
rect 75184 57248 75236 57254
rect 75184 57190 75236 57196
rect 73160 5092 73212 5098
rect 73160 5034 73212 5040
rect 73068 4956 73120 4962
rect 73068 4898 73120 4904
rect 71780 3596 71832 3602
rect 71780 3538 71832 3544
rect 71872 3460 71924 3466
rect 71872 3402 71924 3408
rect 70400 3120 70452 3126
rect 70400 3062 70452 3068
rect 71044 3120 71096 3126
rect 71044 3062 71096 3068
rect 70412 2990 70440 3062
rect 70400 2984 70452 2990
rect 70400 2926 70452 2932
rect 70676 2984 70728 2990
rect 70676 2926 70728 2932
rect 70688 480 70716 2926
rect 71884 480 71912 3402
rect 73080 480 73108 4898
rect 73816 3602 73844 57190
rect 74264 4140 74316 4146
rect 74264 4082 74316 4088
rect 73804 3596 73856 3602
rect 73804 3538 73856 3544
rect 74276 480 74304 4082
rect 75196 3738 75224 57190
rect 75184 3732 75236 3738
rect 75184 3674 75236 3680
rect 75840 626 75868 57258
rect 76656 5228 76708 5234
rect 76656 5170 76708 5176
rect 75472 598 75868 626
rect 75472 480 75500 598
rect 76668 480 76696 5170
rect 77404 5166 77432 60030
rect 78036 57656 78088 57662
rect 78036 57598 78088 57604
rect 77944 56568 77996 56574
rect 77944 56510 77996 56516
rect 77392 5160 77444 5166
rect 77392 5102 77444 5108
rect 77956 3602 77984 56510
rect 77300 3596 77352 3602
rect 77300 3538 77352 3544
rect 77944 3596 77996 3602
rect 77944 3538 77996 3544
rect 77312 2922 77340 3538
rect 78048 3482 78076 57598
rect 78600 57526 78628 60044
rect 78588 57520 78640 57526
rect 78588 57462 78640 57468
rect 79520 57390 79548 60044
rect 80072 60030 80546 60058
rect 79508 57384 79560 57390
rect 79508 57326 79560 57332
rect 79968 57316 80020 57322
rect 79968 57258 80020 57264
rect 79980 3602 80008 57258
rect 80072 3806 80100 60030
rect 81544 57662 81572 60044
rect 81532 57656 81584 57662
rect 81532 57598 81584 57604
rect 82084 57452 82136 57458
rect 82084 57394 82136 57400
rect 80244 5160 80296 5166
rect 80244 5102 80296 5108
rect 80060 3800 80112 3806
rect 80060 3742 80112 3748
rect 79048 3596 79100 3602
rect 79048 3538 79100 3544
rect 79968 3596 80020 3602
rect 79968 3538 80020 3544
rect 77772 3454 78076 3482
rect 77772 3398 77800 3454
rect 77760 3392 77812 3398
rect 77760 3334 77812 3340
rect 77852 3392 77904 3398
rect 77852 3334 77904 3340
rect 77300 2916 77352 2922
rect 77300 2858 77352 2864
rect 77864 480 77892 3334
rect 79060 480 79088 3538
rect 80256 480 80284 5102
rect 81440 3596 81492 3602
rect 81440 3538 81492 3544
rect 81452 480 81480 3538
rect 82096 3058 82124 57394
rect 82464 57254 82492 60044
rect 83476 57526 83504 60044
rect 84304 60030 84502 60058
rect 83464 57520 83516 57526
rect 83464 57462 83516 57468
rect 82728 57384 82780 57390
rect 82728 57326 82780 57332
rect 82452 57248 82504 57254
rect 82452 57190 82504 57196
rect 82636 3732 82688 3738
rect 82636 3674 82688 3680
rect 82084 3052 82136 3058
rect 82084 2994 82136 3000
rect 82648 480 82676 3674
rect 82740 3602 82768 57326
rect 84304 5302 84332 60030
rect 85408 57594 85436 60044
rect 85488 57656 85540 57662
rect 85488 57598 85540 57604
rect 85396 57588 85448 57594
rect 85396 57530 85448 57536
rect 84292 5296 84344 5302
rect 84292 5238 84344 5244
rect 83832 5092 83884 5098
rect 83832 5034 83884 5040
rect 82728 3596 82780 3602
rect 82728 3538 82780 3544
rect 83844 480 83872 5034
rect 85500 3398 85528 57598
rect 86420 57526 86448 60044
rect 86972 60030 87446 60058
rect 86408 57520 86460 57526
rect 86408 57462 86460 57468
rect 86868 57520 86920 57526
rect 86868 57462 86920 57468
rect 86880 3398 86908 57462
rect 86972 3942 87000 60030
rect 87328 6180 87380 6186
rect 87328 6122 87380 6128
rect 86960 3936 87012 3942
rect 86960 3878 87012 3884
rect 84936 3392 84988 3398
rect 84936 3334 84988 3340
rect 85488 3392 85540 3398
rect 85488 3334 85540 3340
rect 86132 3392 86184 3398
rect 86132 3334 86184 3340
rect 86868 3392 86920 3398
rect 86868 3334 86920 3340
rect 84948 480 84976 3334
rect 86144 480 86172 3334
rect 87340 480 87368 6122
rect 88352 3874 88380 60044
rect 89364 57186 89392 60044
rect 90376 57798 90404 60044
rect 90364 57792 90416 57798
rect 90364 57734 90416 57740
rect 91296 57730 91324 60044
rect 91284 57724 91336 57730
rect 91284 57666 91336 57672
rect 89628 57588 89680 57594
rect 89628 57530 89680 57536
rect 89352 57180 89404 57186
rect 89352 57122 89404 57128
rect 88340 3868 88392 3874
rect 88340 3810 88392 3816
rect 89640 3398 89668 57530
rect 92308 57458 92336 60044
rect 93228 57866 93256 60044
rect 93872 60030 94254 60058
rect 93216 57860 93268 57866
rect 93216 57802 93268 57808
rect 93768 57724 93820 57730
rect 93768 57666 93820 57672
rect 92296 57452 92348 57458
rect 92296 57394 92348 57400
rect 91744 56976 91796 56982
rect 91744 56918 91796 56924
rect 90916 5296 90968 5302
rect 90916 5238 90968 5244
rect 89720 3800 89772 3806
rect 89720 3742 89772 3748
rect 88524 3392 88576 3398
rect 88524 3334 88576 3340
rect 89628 3392 89680 3398
rect 89628 3334 89680 3340
rect 88536 480 88564 3334
rect 89732 480 89760 3742
rect 90928 480 90956 5238
rect 91756 2854 91784 56918
rect 93780 4146 93808 57666
rect 93308 4140 93360 4146
rect 93308 4082 93360 4088
rect 93768 4140 93820 4146
rect 93768 4082 93820 4088
rect 92112 3936 92164 3942
rect 92112 3878 92164 3884
rect 91744 2848 91796 2854
rect 91744 2790 91796 2796
rect 92124 480 92152 3878
rect 93320 480 93348 4082
rect 93872 3874 93900 60030
rect 95252 57934 95280 60044
rect 95240 57928 95292 57934
rect 95240 57870 95292 57876
rect 96172 57118 96200 60044
rect 96528 57792 96580 57798
rect 96528 57734 96580 57740
rect 96160 57112 96212 57118
rect 96160 57054 96212 57060
rect 94504 6248 94556 6254
rect 94504 6190 94556 6196
rect 93860 3868 93912 3874
rect 93860 3810 93912 3816
rect 94516 480 94544 6190
rect 96540 4146 96568 57734
rect 97184 57186 97212 60044
rect 97172 57180 97224 57186
rect 97172 57122 97224 57128
rect 98196 56982 98224 60044
rect 99116 58177 99144 60044
rect 99102 58168 99158 58177
rect 99102 58103 99158 58112
rect 98458 58032 98514 58041
rect 98514 57990 98592 58018
rect 98458 57967 98514 57976
rect 98184 56976 98236 56982
rect 98184 56918 98236 56924
rect 98564 48346 98592 57990
rect 98552 48340 98604 48346
rect 98552 48282 98604 48288
rect 100128 48278 100156 60044
rect 100668 57860 100720 57866
rect 100668 57802 100720 57808
rect 98644 48272 98696 48278
rect 98644 48214 98696 48220
rect 100116 48272 100168 48278
rect 100116 48214 100168 48220
rect 98552 46980 98604 46986
rect 98552 46922 98604 46928
rect 98564 46866 98592 46922
rect 98472 46838 98592 46866
rect 98472 38010 98500 46838
rect 98276 38004 98328 38010
rect 98276 37946 98328 37952
rect 98460 38004 98512 38010
rect 98460 37946 98512 37952
rect 98288 29073 98316 37946
rect 98274 29064 98330 29073
rect 98274 28999 98330 29008
rect 98458 29064 98514 29073
rect 98458 28999 98514 29008
rect 98472 28966 98500 28999
rect 98000 28960 98052 28966
rect 98000 28902 98052 28908
rect 98460 28960 98512 28966
rect 98460 28902 98512 28908
rect 98012 12458 98040 28902
rect 98012 12430 98224 12458
rect 98196 5370 98224 12430
rect 98184 5364 98236 5370
rect 98184 5306 98236 5312
rect 98092 4684 98144 4690
rect 98092 4626 98144 4632
rect 95700 4140 95752 4146
rect 95700 4082 95752 4088
rect 96528 4140 96580 4146
rect 96528 4082 96580 4088
rect 95712 480 95740 4082
rect 96896 3868 96948 3874
rect 96896 3810 96948 3816
rect 96908 480 96936 3810
rect 98104 480 98132 4626
rect 98656 3330 98684 48214
rect 98644 3324 98696 3330
rect 98644 3266 98696 3272
rect 99288 3120 99340 3126
rect 99288 3062 99340 3068
rect 99300 480 99328 3062
rect 100680 626 100708 57802
rect 101140 57050 101168 60044
rect 101128 57044 101180 57050
rect 101128 56986 101180 56992
rect 101232 52358 101260 60166
rect 102876 57180 102928 57186
rect 102876 57122 102928 57128
rect 102784 56704 102836 56710
rect 102784 56646 102836 56652
rect 101220 52352 101272 52358
rect 101220 52294 101272 52300
rect 100852 48340 100904 48346
rect 100852 48282 100904 48288
rect 100864 43466 100892 48282
rect 100864 43438 101076 43466
rect 101048 38622 101076 43438
rect 101036 38616 101088 38622
rect 101036 38558 101088 38564
rect 101220 31680 101272 31686
rect 101220 31622 101272 31628
rect 101232 28966 101260 31622
rect 100760 28960 100812 28966
rect 100760 28902 100812 28908
rect 101220 28960 101272 28966
rect 101220 28902 101272 28908
rect 100772 12458 100800 28902
rect 100772 12430 100984 12458
rect 100956 5506 100984 12430
rect 100944 5500 100996 5506
rect 100944 5442 100996 5448
rect 101588 5364 101640 5370
rect 101588 5306 101640 5312
rect 100496 598 100708 626
rect 100496 480 100524 598
rect 101600 480 101628 5306
rect 102796 3262 102824 56646
rect 102784 3256 102836 3262
rect 102784 3198 102836 3204
rect 102888 3194 102916 57122
rect 103072 56846 103100 60044
rect 103060 56840 103112 56846
rect 103060 56782 103112 56788
rect 104084 56710 104112 60044
rect 104164 57860 104216 57866
rect 104164 57802 104216 57808
rect 104072 56704 104124 56710
rect 104072 56646 104124 56652
rect 104176 4010 104204 57802
rect 105004 4758 105032 60044
rect 106016 57186 106044 60044
rect 106004 57180 106056 57186
rect 106004 57122 106056 57128
rect 105544 57044 105596 57050
rect 105544 56986 105596 56992
rect 105176 5500 105228 5506
rect 105176 5442 105228 5448
rect 104992 4752 105044 4758
rect 104992 4694 105044 4700
rect 104164 4004 104216 4010
rect 104164 3946 104216 3952
rect 102876 3188 102928 3194
rect 102876 3130 102928 3136
rect 103980 3188 104032 3194
rect 103980 3130 104032 3136
rect 102784 2916 102836 2922
rect 102784 2858 102836 2864
rect 102796 480 102824 2858
rect 103992 480 104020 3130
rect 105188 480 105216 5442
rect 105556 2990 105584 56986
rect 107028 56914 107056 60044
rect 107764 60030 107962 60058
rect 108592 60030 108974 60058
rect 107568 57180 107620 57186
rect 107568 57122 107620 57128
rect 107016 56908 107068 56914
rect 107016 56850 107068 56856
rect 107580 3262 107608 57122
rect 107764 5438 107792 60030
rect 108592 56982 108620 60030
rect 108948 57928 109000 57934
rect 108948 57870 109000 57876
rect 108580 56976 108632 56982
rect 108580 56918 108632 56924
rect 108304 56772 108356 56778
rect 108304 56714 108356 56720
rect 107752 5432 107804 5438
rect 107752 5374 107804 5380
rect 108316 3670 108344 56714
rect 108304 3664 108356 3670
rect 108304 3606 108356 3612
rect 107660 3324 107712 3330
rect 107660 3266 107712 3272
rect 106372 3256 106424 3262
rect 106372 3198 106424 3204
rect 107568 3256 107620 3262
rect 107568 3198 107620 3204
rect 105544 2984 105596 2990
rect 105544 2926 105596 2932
rect 106384 480 106412 3198
rect 107672 3108 107700 3266
rect 107580 3080 107700 3108
rect 107580 480 107608 3080
rect 108960 626 108988 57870
rect 109880 56778 109908 60044
rect 110432 60030 110906 60058
rect 109868 56772 109920 56778
rect 109868 56714 109920 56720
rect 109684 56636 109736 56642
rect 109684 56578 109736 56584
rect 109696 3398 109724 56578
rect 110432 4826 110460 60030
rect 111904 57866 111932 60044
rect 111892 57860 111944 57866
rect 111892 57802 111944 57808
rect 112824 57118 112852 60044
rect 113192 60030 113850 60058
rect 113088 57928 113140 57934
rect 113088 57870 113140 57876
rect 112812 57112 112864 57118
rect 112812 57054 112864 57060
rect 111064 56976 111116 56982
rect 111064 56918 111116 56924
rect 111076 6390 111104 56918
rect 112444 56840 112496 56846
rect 112444 56782 112496 56788
rect 111064 6384 111116 6390
rect 111064 6326 111116 6332
rect 110420 4820 110472 4826
rect 110420 4762 110472 4768
rect 112352 4140 112404 4146
rect 112352 4082 112404 4088
rect 111156 4072 111208 4078
rect 111156 4014 111208 4020
rect 109960 3664 110012 3670
rect 109960 3606 110012 3612
rect 109684 3392 109736 3398
rect 109684 3334 109736 3340
rect 108776 598 108988 626
rect 108776 480 108804 598
rect 109972 480 110000 3606
rect 111168 480 111196 4014
rect 112364 480 112392 4082
rect 112456 3942 112484 56782
rect 113100 4146 113128 57870
rect 113192 4894 113220 60030
rect 114468 56908 114520 56914
rect 114468 56850 114520 56856
rect 113180 4888 113232 4894
rect 113180 4830 113232 4836
rect 114480 4146 114508 56850
rect 114848 56710 114876 60044
rect 115204 57248 115256 57254
rect 115204 57190 115256 57196
rect 115294 57216 115350 57225
rect 114836 56704 114888 56710
rect 114836 56646 114888 56652
rect 113088 4140 113140 4146
rect 113088 4082 113140 4088
rect 113548 4140 113600 4146
rect 113548 4082 113600 4088
rect 114468 4140 114520 4146
rect 114468 4082 114520 4088
rect 112444 3936 112496 3942
rect 112444 3878 112496 3884
rect 113560 480 113588 4082
rect 115216 3466 115244 57190
rect 115294 57151 115350 57160
rect 115308 3738 115336 57151
rect 115768 56642 115796 60044
rect 115952 60030 116794 60058
rect 115756 56636 115808 56642
rect 115756 56578 115808 56584
rect 115952 5030 115980 60030
rect 117228 57112 117280 57118
rect 117228 57054 117280 57060
rect 115940 5024 115992 5030
rect 115940 4966 115992 4972
rect 117240 3738 117268 57054
rect 117792 57050 117820 60044
rect 118712 57254 118740 60044
rect 118804 60030 119738 60058
rect 118700 57248 118752 57254
rect 118700 57190 118752 57196
rect 117780 57044 117832 57050
rect 117780 56986 117832 56992
rect 117964 57044 118016 57050
rect 117964 56986 118016 56992
rect 115296 3732 115348 3738
rect 115296 3674 115348 3680
rect 115940 3732 115992 3738
rect 115940 3674 115992 3680
rect 117228 3732 117280 3738
rect 117228 3674 117280 3680
rect 115204 3460 115256 3466
rect 115204 3402 115256 3408
rect 114744 3392 114796 3398
rect 114744 3334 114796 3340
rect 114756 480 114784 3334
rect 115952 480 115980 3674
rect 117976 3602 118004 56986
rect 118804 4962 118832 60030
rect 119988 57044 120040 57050
rect 119988 56986 120040 56992
rect 119344 56772 119396 56778
rect 119344 56714 119396 56720
rect 118792 4956 118844 4962
rect 118792 4898 118844 4904
rect 118240 3936 118292 3942
rect 118240 3878 118292 3884
rect 117964 3596 118016 3602
rect 117964 3538 118016 3544
rect 117136 3460 117188 3466
rect 117136 3402 117188 3408
rect 117148 480 117176 3402
rect 118252 480 118280 3878
rect 119356 3126 119384 56714
rect 120000 4146 120028 56986
rect 120736 56710 120764 60044
rect 121472 60030 121670 60058
rect 121472 57066 121500 60030
rect 121288 57038 121500 57066
rect 121288 56982 121316 57038
rect 121276 56976 121328 56982
rect 121276 56918 121328 56924
rect 121368 56976 121420 56982
rect 121368 56918 121420 56924
rect 120724 56704 120776 56710
rect 120724 56646 120776 56652
rect 121380 4146 121408 56918
rect 121748 51610 121776 60166
rect 122852 60030 123694 60058
rect 122852 57610 122880 60030
rect 122484 57594 122880 57610
rect 122472 57588 122880 57594
rect 122524 57582 122880 57588
rect 122472 57530 122524 57536
rect 124128 57452 124180 57458
rect 124128 57394 124180 57400
rect 122104 56704 122156 56710
rect 122104 56646 122156 56652
rect 121736 51604 121788 51610
rect 121736 51546 121788 51552
rect 121552 48340 121604 48346
rect 121552 48282 121604 48288
rect 121564 41426 121592 48282
rect 121472 41410 121592 41426
rect 121460 41404 121592 41410
rect 121512 41398 121592 41404
rect 121644 41404 121696 41410
rect 121460 41346 121512 41352
rect 121644 41346 121696 41352
rect 121656 31822 121684 41346
rect 121644 31816 121696 31822
rect 121644 31758 121696 31764
rect 121736 31680 121788 31686
rect 121736 31622 121788 31628
rect 121748 27606 121776 31622
rect 121736 27600 121788 27606
rect 121736 27542 121788 27548
rect 121644 18012 121696 18018
rect 121644 17954 121696 17960
rect 121656 12510 121684 17954
rect 121644 12504 121696 12510
rect 121644 12446 121696 12452
rect 121552 12436 121604 12442
rect 121552 12378 121604 12384
rect 121564 5234 121592 12378
rect 121552 5228 121604 5234
rect 121552 5170 121604 5176
rect 119436 4140 119488 4146
rect 119436 4082 119488 4088
rect 119988 4140 120040 4146
rect 119988 4082 120040 4088
rect 120632 4140 120684 4146
rect 120632 4082 120684 4088
rect 121368 4140 121420 4146
rect 121368 4082 121420 4088
rect 119344 3120 119396 3126
rect 119344 3062 119396 3068
rect 119448 480 119476 4082
rect 120644 480 120672 4082
rect 121828 4004 121880 4010
rect 121828 3946 121880 3952
rect 121840 480 121868 3946
rect 122116 2922 122144 56646
rect 122196 56636 122248 56642
rect 122196 56578 122248 56584
rect 122208 3806 122236 56578
rect 124140 4146 124168 57394
rect 124600 57390 124628 60044
rect 124588 57384 124640 57390
rect 124588 57326 124640 57332
rect 125508 57248 125560 57254
rect 125508 57190 125560 57196
rect 123024 4140 123076 4146
rect 123024 4082 123076 4088
rect 124128 4140 124180 4146
rect 124128 4082 124180 4088
rect 122196 3800 122248 3806
rect 122196 3742 122248 3748
rect 122104 2916 122156 2922
rect 122104 2858 122156 2864
rect 123036 480 123064 4082
rect 125520 3738 125548 57190
rect 125612 5166 125640 60044
rect 126164 60030 126546 60058
rect 126164 57390 126192 60030
rect 126152 57384 126204 57390
rect 126152 57326 126204 57332
rect 126244 57384 126296 57390
rect 126244 57326 126296 57332
rect 125600 5160 125652 5166
rect 125600 5102 125652 5108
rect 126256 3874 126284 57326
rect 127544 57225 127572 60044
rect 128464 60030 128570 60058
rect 127530 57216 127586 57225
rect 127530 57151 127586 57160
rect 128464 5098 128492 60030
rect 129476 57526 129504 60044
rect 130488 57594 130516 60044
rect 131224 60030 131514 60058
rect 130476 57588 130528 57594
rect 130476 57530 130528 57536
rect 129464 57520 129516 57526
rect 129464 57462 129516 57468
rect 129004 48340 129056 48346
rect 129004 48282 129056 48288
rect 129016 41426 129044 48282
rect 128832 41398 129044 41426
rect 128832 37262 128860 41398
rect 128820 37256 128872 37262
rect 128820 37198 128872 37204
rect 128636 27736 128688 27742
rect 128636 27678 128688 27684
rect 128648 27606 128676 27678
rect 128636 27600 128688 27606
rect 128636 27542 128688 27548
rect 128912 19236 128964 19242
rect 128912 19178 128964 19184
rect 128924 12510 128952 19178
rect 128912 12504 128964 12510
rect 128912 12446 128964 12452
rect 128912 12368 128964 12374
rect 128912 12310 128964 12316
rect 128452 5092 128504 5098
rect 128452 5034 128504 5040
rect 127808 4888 127860 4894
rect 127808 4830 127860 4836
rect 126244 3868 126296 3874
rect 126244 3810 126296 3816
rect 124220 3732 124272 3738
rect 124220 3674 124272 3680
rect 125508 3732 125560 3738
rect 125508 3674 125560 3680
rect 124232 480 124260 3674
rect 125416 3596 125468 3602
rect 125416 3538 125468 3544
rect 125428 480 125456 3538
rect 126612 3528 126664 3534
rect 126612 3470 126664 3476
rect 126624 480 126652 3470
rect 127820 480 127848 4830
rect 128924 3262 128952 12310
rect 131224 6186 131252 60030
rect 132420 57526 132448 60044
rect 133432 57594 133460 60044
rect 133892 60030 134458 60058
rect 133420 57588 133472 57594
rect 133420 57530 133472 57536
rect 132408 57520 132460 57526
rect 132408 57462 132460 57468
rect 131212 6180 131264 6186
rect 131212 6122 131264 6128
rect 133892 5302 133920 60030
rect 135364 56642 135392 60044
rect 136376 57662 136404 60044
rect 136652 60030 137402 60058
rect 136364 57656 136416 57662
rect 136364 57598 136416 57604
rect 136548 57452 136600 57458
rect 136548 57394 136600 57400
rect 135904 56840 135956 56846
rect 135904 56782 135956 56788
rect 135352 56636 135404 56642
rect 135352 56578 135404 56584
rect 133880 5296 133932 5302
rect 133880 5238 133932 5244
rect 134892 5092 134944 5098
rect 134892 5034 134944 5040
rect 131396 5024 131448 5030
rect 131396 4966 131448 4972
rect 129004 4820 129056 4826
rect 129004 4762 129056 4768
rect 128912 3256 128964 3262
rect 128912 3198 128964 3204
rect 129016 480 129044 4762
rect 130200 3868 130252 3874
rect 130200 3810 130252 3816
rect 130212 480 130240 3810
rect 131408 480 131436 4966
rect 132592 4956 132644 4962
rect 132592 4898 132644 4904
rect 132604 480 132632 4898
rect 133788 3800 133840 3806
rect 133788 3742 133840 3748
rect 133800 480 133828 3742
rect 134904 480 134932 5034
rect 135916 3330 135944 56782
rect 136560 4146 136588 57394
rect 136652 6254 136680 60030
rect 138308 57730 138336 60044
rect 138296 57724 138348 57730
rect 138296 57666 138348 57672
rect 139124 57724 139176 57730
rect 139124 57666 139176 57672
rect 139136 54346 139164 57666
rect 139320 57390 139348 60044
rect 139412 60030 140346 60058
rect 139308 57384 139360 57390
rect 139308 57326 139360 57332
rect 139136 54318 139348 54346
rect 136640 6248 136692 6254
rect 136640 6190 136692 6196
rect 139320 4146 139348 54318
rect 139412 4690 139440 60030
rect 140688 57656 140740 57662
rect 140688 57598 140740 57604
rect 139400 4684 139452 4690
rect 139400 4626 139452 4632
rect 136088 4140 136140 4146
rect 136088 4082 136140 4088
rect 136548 4140 136600 4146
rect 136548 4082 136600 4088
rect 138480 4140 138532 4146
rect 138480 4082 138532 4088
rect 139308 4140 139360 4146
rect 139308 4082 139360 4088
rect 135904 3324 135956 3330
rect 135904 3266 135956 3272
rect 136100 480 136128 4082
rect 137284 3732 137336 3738
rect 137284 3674 137336 3680
rect 137296 480 137324 3674
rect 138492 480 138520 4082
rect 140700 2990 140728 57598
rect 141252 56778 141280 60044
rect 142264 57798 142292 60044
rect 142356 60030 143198 60058
rect 142252 57792 142304 57798
rect 142252 57734 142304 57740
rect 142068 57180 142120 57186
rect 142068 57122 142120 57128
rect 141240 56772 141292 56778
rect 141240 56714 141292 56720
rect 140872 4140 140924 4146
rect 140872 4082 140924 4088
rect 139676 2984 139728 2990
rect 139676 2926 139728 2932
rect 140688 2984 140740 2990
rect 140688 2926 140740 2932
rect 139688 480 139716 2926
rect 140884 480 140912 4082
rect 142080 480 142108 57122
rect 142356 5370 142384 60030
rect 142804 57792 142856 57798
rect 142804 57734 142856 57740
rect 142344 5364 142396 5370
rect 142344 5306 142396 5312
rect 142816 4078 142844 57734
rect 143448 56840 143500 56846
rect 143448 56782 143500 56788
rect 142804 4072 142856 4078
rect 142804 4014 142856 4020
rect 143460 2854 143488 56782
rect 144196 56710 144224 60044
rect 145208 57526 145236 60044
rect 145196 57520 145248 57526
rect 145196 57462 145248 57468
rect 144184 56704 144236 56710
rect 144184 56646 144236 56652
rect 145300 48346 145328 60166
rect 147140 57594 147168 60044
rect 147588 57724 147640 57730
rect 147588 57666 147640 57672
rect 147128 57588 147180 57594
rect 147128 57530 147180 57536
rect 146206 57216 146262 57225
rect 146206 57151 146262 57160
rect 145564 56636 145616 56642
rect 145564 56578 145616 56584
rect 145196 48340 145248 48346
rect 145196 48282 145248 48288
rect 145288 48340 145340 48346
rect 145288 48282 145340 48288
rect 145208 41562 145236 48282
rect 145116 41534 145236 41562
rect 145116 38690 145144 41534
rect 145012 38684 145064 38690
rect 145012 38626 145064 38632
rect 145104 38684 145156 38690
rect 145104 38626 145156 38632
rect 145024 35766 145052 38626
rect 145012 35760 145064 35766
rect 145012 35702 145064 35708
rect 145196 29028 145248 29034
rect 145196 28970 145248 28976
rect 145208 22250 145236 28970
rect 145116 22222 145236 22250
rect 145116 19378 145144 22222
rect 145012 19372 145064 19378
rect 145012 19314 145064 19320
rect 145104 19372 145156 19378
rect 145104 19314 145156 19320
rect 145024 12458 145052 19314
rect 145024 12430 145144 12458
rect 145116 5506 145144 12430
rect 145104 5500 145156 5506
rect 145104 5442 145156 5448
rect 144460 4072 144512 4078
rect 144460 4014 144512 4020
rect 143448 2848 143500 2854
rect 143448 2790 143500 2796
rect 143264 604 143316 610
rect 143264 546 143316 552
rect 143276 480 143304 546
rect 144472 480 144500 4014
rect 145576 3398 145604 56578
rect 146220 4146 146248 57151
rect 145656 4140 145708 4146
rect 145656 4082 145708 4088
rect 146208 4140 146260 4146
rect 146208 4082 146260 4088
rect 145564 3392 145616 3398
rect 145564 3334 145616 3340
rect 145668 480 145696 4082
rect 147600 3398 147628 57666
rect 148152 56710 148180 60044
rect 149072 57866 149100 60044
rect 149164 60030 150098 60058
rect 149060 57860 149112 57866
rect 149060 57802 149112 57808
rect 148140 56704 148192 56710
rect 148140 56646 148192 56652
rect 148048 5160 148100 5166
rect 148048 5102 148100 5108
rect 146852 3392 146904 3398
rect 146852 3334 146904 3340
rect 147588 3392 147640 3398
rect 147588 3334 147640 3340
rect 146864 480 146892 3334
rect 148060 480 148088 5102
rect 149164 3670 149192 60030
rect 150348 57860 150400 57866
rect 150348 57802 150400 57808
rect 150360 3942 150388 57802
rect 151096 57798 151124 60044
rect 152016 57934 152044 60044
rect 152004 57928 152056 57934
rect 152004 57870 152056 57876
rect 152464 57928 152516 57934
rect 152464 57870 152516 57876
rect 151084 57792 151136 57798
rect 151084 57734 151136 57740
rect 149244 3936 149296 3942
rect 149244 3878 149296 3884
rect 150348 3936 150400 3942
rect 150348 3878 150400 3884
rect 149152 3664 149204 3670
rect 149152 3606 149204 3612
rect 149256 480 149284 3878
rect 151544 3664 151596 3670
rect 151544 3606 151596 3612
rect 150440 3392 150492 3398
rect 150440 3334 150492 3340
rect 150452 480 150480 3334
rect 151556 480 151584 3606
rect 152476 3466 152504 57870
rect 153028 56914 153056 60044
rect 153844 57792 153896 57798
rect 153844 57734 153896 57740
rect 153108 57180 153160 57186
rect 153108 57122 153160 57128
rect 153016 56908 153068 56914
rect 153016 56850 153068 56856
rect 152464 3460 152516 3466
rect 152464 3402 152516 3408
rect 153120 3346 153148 57122
rect 152752 3318 153148 3346
rect 153856 3330 153884 57734
rect 154040 56642 154068 60044
rect 154960 57118 154988 60044
rect 155972 57798 156000 60044
rect 156984 57934 157012 60044
rect 156972 57928 157024 57934
rect 156972 57870 157024 57876
rect 155960 57792 156012 57798
rect 155960 57734 156012 57740
rect 157248 57180 157300 57186
rect 157248 57122 157300 57128
rect 154948 57112 155000 57118
rect 154948 57054 155000 57060
rect 156604 57112 156656 57118
rect 156604 57054 156656 57060
rect 154028 56636 154080 56642
rect 154028 56578 154080 56584
rect 155132 5228 155184 5234
rect 155132 5170 155184 5176
rect 153936 3936 153988 3942
rect 153936 3878 153988 3884
rect 153844 3324 153896 3330
rect 152752 480 152780 3318
rect 153844 3266 153896 3272
rect 153948 480 153976 3878
rect 155144 480 155172 5170
rect 156616 4010 156644 57054
rect 156604 4004 156656 4010
rect 156604 3946 156656 3952
rect 157260 3466 157288 57122
rect 157904 57050 157932 60044
rect 158628 57928 158680 57934
rect 158628 57870 158680 57876
rect 157892 57044 157944 57050
rect 157892 56986 157944 56992
rect 158640 3466 158668 57870
rect 158916 56982 158944 60044
rect 159836 57118 159864 60044
rect 160848 57254 160876 60044
rect 161860 57322 161888 60044
rect 161848 57316 161900 57322
rect 161848 57258 161900 57264
rect 160836 57248 160888 57254
rect 160836 57190 160888 57196
rect 159824 57112 159876 57118
rect 159824 57054 159876 57060
rect 160008 57112 160060 57118
rect 160008 57054 160060 57060
rect 159916 57044 159968 57050
rect 159916 56986 159968 56992
rect 158904 56976 158956 56982
rect 158904 56918 158956 56924
rect 159928 3602 159956 56986
rect 158720 3596 158772 3602
rect 158720 3538 158772 3544
rect 159916 3596 159968 3602
rect 159916 3538 159968 3544
rect 156328 3460 156380 3466
rect 156328 3402 156380 3408
rect 157248 3460 157300 3466
rect 157248 3402 157300 3408
rect 157524 3460 157576 3466
rect 157524 3402 157576 3408
rect 158628 3460 158680 3466
rect 158628 3402 158680 3408
rect 156340 480 156368 3402
rect 157536 480 157564 3402
rect 158732 480 158760 3538
rect 160020 3482 160048 57054
rect 162780 56642 162808 60044
rect 162964 60030 163806 60058
rect 164252 60030 164818 60058
rect 160744 56636 160796 56642
rect 160744 56578 160796 56584
rect 162768 56636 162820 56642
rect 162768 56578 162820 56584
rect 160756 4010 160784 56578
rect 160744 4004 160796 4010
rect 160744 3946 160796 3952
rect 161112 4004 161164 4010
rect 161112 3946 161164 3952
rect 159928 3454 160048 3482
rect 159928 480 159956 3454
rect 161124 480 161152 3946
rect 162964 3534 162992 60030
rect 164148 56908 164200 56914
rect 164148 56850 164200 56856
rect 164160 3534 164188 56850
rect 164252 4894 164280 60030
rect 165528 56976 165580 56982
rect 165528 56918 165580 56924
rect 164884 56636 164936 56642
rect 164884 56578 164936 56584
rect 164240 4888 164292 4894
rect 164240 4830 164292 4836
rect 162952 3528 163004 3534
rect 162952 3470 163004 3476
rect 163504 3528 163556 3534
rect 163504 3470 163556 3476
rect 164148 3528 164200 3534
rect 164148 3470 164200 3476
rect 164700 3528 164752 3534
rect 164700 3470 164752 3476
rect 162308 3460 162360 3466
rect 162308 3402 162360 3408
rect 162320 480 162348 3402
rect 163516 480 163544 3470
rect 164712 480 164740 3470
rect 164896 3398 164924 56578
rect 165540 3534 165568 56918
rect 165620 55888 165672 55894
rect 165620 55830 165672 55836
rect 165632 3874 165660 55830
rect 165724 4826 165752 60044
rect 166368 60030 166750 60058
rect 167012 60030 167762 60058
rect 168484 60030 168682 60058
rect 169312 60030 169694 60058
rect 169772 60030 170706 60058
rect 166368 55894 166396 60030
rect 166356 55888 166408 55894
rect 166356 55830 166408 55836
rect 167012 5030 167040 60030
rect 168380 57316 168432 57322
rect 168380 57258 168432 57264
rect 168196 57248 168248 57254
rect 168196 57190 168248 57196
rect 167000 5024 167052 5030
rect 167000 4966 167052 4972
rect 165712 4820 165764 4826
rect 165712 4762 165764 4768
rect 165620 3868 165672 3874
rect 165620 3810 165672 3816
rect 165528 3528 165580 3534
rect 165528 3470 165580 3476
rect 165896 3528 165948 3534
rect 165896 3470 165948 3476
rect 164884 3392 164936 3398
rect 164884 3334 164936 3340
rect 165908 480 165936 3470
rect 167092 3188 167144 3194
rect 167092 3130 167144 3136
rect 167104 480 167132 3130
rect 168208 480 168236 57190
rect 168288 56840 168340 56846
rect 168288 56782 168340 56788
rect 168300 3194 168328 56782
rect 168392 3806 168420 57258
rect 168484 4962 168512 60030
rect 169312 57322 169340 60030
rect 169300 57316 169352 57322
rect 169300 57258 169352 57264
rect 169024 56704 169076 56710
rect 169024 56646 169076 56652
rect 168472 4956 168524 4962
rect 168472 4898 168524 4904
rect 169036 3942 169064 56646
rect 169772 5098 169800 60030
rect 171612 57390 171640 60044
rect 172638 60030 172744 60058
rect 171600 57384 171652 57390
rect 171600 57326 171652 57332
rect 172428 56908 172480 56914
rect 172428 56850 172480 56856
rect 171048 56772 171100 56778
rect 171048 56714 171100 56720
rect 169760 5092 169812 5098
rect 169760 5034 169812 5040
rect 169024 3936 169076 3942
rect 169024 3878 169076 3884
rect 168380 3800 168432 3806
rect 168380 3742 168432 3748
rect 169392 3596 169444 3602
rect 169392 3538 169444 3544
rect 168288 3188 168340 3194
rect 168288 3130 168340 3136
rect 169404 480 169432 3538
rect 171060 3058 171088 56714
rect 172440 3058 172468 56850
rect 172716 3330 172744 60030
rect 173636 57662 173664 60044
rect 173624 57656 173676 57662
rect 173624 57598 173676 57604
rect 174556 57458 174584 60044
rect 175384 60030 175582 60058
rect 174544 57452 174596 57458
rect 174544 57394 174596 57400
rect 175188 57452 175240 57458
rect 175188 57394 175240 57400
rect 173164 56636 173216 56642
rect 173164 56578 173216 56584
rect 173176 3942 173204 56578
rect 173164 3936 173216 3942
rect 173164 3878 173216 3884
rect 172980 3800 173032 3806
rect 172980 3742 173032 3748
rect 172704 3324 172756 3330
rect 172704 3266 172756 3272
rect 170588 3052 170640 3058
rect 170588 2994 170640 3000
rect 171048 3052 171100 3058
rect 171048 2994 171100 3000
rect 171784 3052 171836 3058
rect 171784 2994 171836 3000
rect 172428 3052 172480 3058
rect 172428 2994 172480 3000
rect 170600 480 170628 2994
rect 171796 480 171824 2994
rect 172992 480 173020 3742
rect 175200 3398 175228 57394
rect 175384 4146 175412 60030
rect 176488 57594 176516 60044
rect 176568 57656 176620 57662
rect 176568 57598 176620 57604
rect 176476 57588 176528 57594
rect 176476 57530 176528 57536
rect 175372 4140 175424 4146
rect 175372 4082 175424 4088
rect 176476 3732 176528 3738
rect 176476 3674 176528 3680
rect 174176 3392 174228 3398
rect 174176 3334 174228 3340
rect 175188 3392 175240 3398
rect 175188 3334 175240 3340
rect 175372 3392 175424 3398
rect 175372 3334 175424 3340
rect 174188 480 174216 3334
rect 175384 480 175412 3334
rect 176488 1850 176516 3674
rect 176580 3398 176608 57598
rect 177500 57526 177528 60044
rect 178052 60030 178526 60058
rect 177488 57520 177540 57526
rect 177488 57462 177540 57468
rect 177948 57452 178000 57458
rect 177948 57394 178000 57400
rect 176568 3392 176620 3398
rect 177960 3346 177988 57394
rect 178052 4078 178080 60030
rect 179328 57384 179380 57390
rect 179328 57326 179380 57332
rect 178040 4072 178092 4078
rect 178040 4014 178092 4020
rect 179340 3346 179368 57326
rect 179432 57225 179460 60044
rect 180444 57730 180472 60044
rect 180812 60030 181470 60058
rect 180432 57724 180484 57730
rect 180432 57666 180484 57672
rect 179418 57216 179474 57225
rect 179418 57151 179474 57160
rect 180812 5166 180840 60030
rect 182376 57866 182404 60044
rect 182364 57860 182416 57866
rect 182364 57802 182416 57808
rect 182088 57724 182140 57730
rect 182088 57666 182140 57672
rect 180800 5160 180852 5166
rect 180800 5102 180852 5108
rect 180156 3868 180208 3874
rect 180156 3810 180208 3816
rect 176568 3334 176620 3340
rect 177776 3318 177988 3346
rect 178972 3318 179368 3346
rect 176488 1822 176608 1850
rect 176580 480 176608 1822
rect 177776 480 177804 3318
rect 178972 480 179000 3318
rect 180168 480 180196 3810
rect 182100 3398 182128 57666
rect 183388 57594 183416 60044
rect 183572 60030 184414 60058
rect 183468 57860 183520 57866
rect 183468 57802 183520 57808
rect 183376 57588 183428 57594
rect 183376 57530 183428 57536
rect 183480 3398 183508 57802
rect 183572 3670 183600 60030
rect 185320 57798 185348 60044
rect 185308 57792 185360 57798
rect 185308 57734 185360 57740
rect 186228 57792 186280 57798
rect 186228 57734 186280 57740
rect 184848 57588 184900 57594
rect 184848 57530 184900 57536
rect 183744 4004 183796 4010
rect 183744 3946 183796 3952
rect 183560 3664 183612 3670
rect 183560 3606 183612 3612
rect 181352 3392 181404 3398
rect 181352 3334 181404 3340
rect 182088 3392 182140 3398
rect 182088 3334 182140 3340
rect 182548 3392 182600 3398
rect 182548 3334 182600 3340
rect 183468 3392 183520 3398
rect 183468 3334 183520 3340
rect 181364 480 181392 3334
rect 182560 480 182588 3334
rect 183756 480 183784 3946
rect 184860 480 184888 57530
rect 186240 3346 186268 57734
rect 186332 56574 186360 60044
rect 186424 60030 187358 60058
rect 186320 56568 186372 56574
rect 186320 56510 186372 56516
rect 186424 5234 186452 60030
rect 188264 57186 188292 60044
rect 189276 57934 189304 60044
rect 189264 57928 189316 57934
rect 189264 57870 189316 57876
rect 188252 57180 188304 57186
rect 188252 57122 188304 57128
rect 188988 57180 189040 57186
rect 188988 57122 189040 57128
rect 186412 5228 186464 5234
rect 186412 5170 186464 5176
rect 187240 3664 187292 3670
rect 187240 3606 187292 3612
rect 186056 3318 186268 3346
rect 186056 480 186084 3318
rect 187252 480 187280 3606
rect 189000 3058 189028 57122
rect 190288 57050 190316 60044
rect 190368 57928 190420 57934
rect 190368 57870 190420 57876
rect 190276 57044 190328 57050
rect 190276 56986 190328 56992
rect 190380 3126 190408 57870
rect 191208 57118 191236 60044
rect 191196 57112 191248 57118
rect 191196 57054 191248 57060
rect 192220 56642 192248 60044
rect 192208 56636 192260 56642
rect 192208 56578 192260 56584
rect 192312 55570 192340 60166
rect 194152 57322 194180 60044
rect 194140 57316 194192 57322
rect 194140 57258 194192 57264
rect 193128 57112 193180 57118
rect 193128 57054 193180 57060
rect 192128 55542 192340 55570
rect 192128 38622 192156 55542
rect 192116 38616 192168 38622
rect 192116 38558 192168 38564
rect 192024 29028 192076 29034
rect 192024 28970 192076 28976
rect 192036 22114 192064 28970
rect 192036 22086 192248 22114
rect 192220 19310 192248 22086
rect 192208 19304 192260 19310
rect 192208 19246 192260 19252
rect 192300 9716 192352 9722
rect 192300 9658 192352 9664
rect 190828 4072 190880 4078
rect 190828 4014 190880 4020
rect 189632 3120 189684 3126
rect 189632 3062 189684 3068
rect 190368 3120 190420 3126
rect 190368 3062 190420 3068
rect 188436 3052 188488 3058
rect 188436 2994 188488 3000
rect 188988 3052 189040 3058
rect 188988 2994 189040 3000
rect 188448 480 188476 2994
rect 189644 480 189672 3062
rect 190840 480 190868 4014
rect 192312 3466 192340 9658
rect 192300 3460 192352 3466
rect 192300 3402 192352 3408
rect 193140 3398 193168 57054
rect 195164 56982 195192 60044
rect 195152 56976 195204 56982
rect 195152 56918 195204 56924
rect 194508 56636 194560 56642
rect 194508 56578 194560 56584
rect 194520 4146 194548 56578
rect 195888 48340 195940 48346
rect 195888 48282 195940 48288
rect 195900 38622 195928 48282
rect 195888 38616 195940 38622
rect 195888 38558 195940 38564
rect 195888 29028 195940 29034
rect 195888 28970 195940 28976
rect 195900 19514 195928 28970
rect 195888 19508 195940 19514
rect 195888 19450 195940 19456
rect 195888 19372 195940 19378
rect 195888 19314 195940 19320
rect 195900 19281 195928 19314
rect 195886 19272 195942 19281
rect 195886 19207 195942 19216
rect 195886 9752 195942 9761
rect 195886 9687 195942 9696
rect 195900 9654 195928 9687
rect 195888 9648 195940 9654
rect 195888 9590 195940 9596
rect 193220 4140 193272 4146
rect 193220 4082 193272 4088
rect 194508 4140 194560 4146
rect 194508 4082 194560 4088
rect 192024 3392 192076 3398
rect 192024 3334 192076 3340
rect 193128 3392 193180 3398
rect 193128 3334 193180 3340
rect 192036 480 192064 3334
rect 193232 480 193260 4082
rect 196084 3602 196112 60044
rect 197096 56846 197124 60044
rect 198108 57254 198136 60044
rect 198844 60030 199042 60058
rect 199672 60030 200054 60058
rect 198096 57248 198148 57254
rect 198096 57190 198148 57196
rect 198648 57248 198700 57254
rect 198648 57190 198700 57196
rect 197268 57044 197320 57050
rect 197268 56986 197320 56992
rect 197084 56840 197136 56846
rect 197084 56782 197136 56788
rect 196162 19272 196218 19281
rect 196162 19207 196218 19216
rect 196176 9761 196204 19207
rect 196162 9752 196218 9761
rect 196162 9687 196218 9696
rect 197280 4146 197308 56986
rect 196808 4140 196860 4146
rect 196808 4082 196860 4088
rect 197268 4140 197320 4146
rect 197268 4082 197320 4088
rect 196072 3596 196124 3602
rect 196072 3538 196124 3544
rect 194416 3460 194468 3466
rect 194416 3402 194468 3408
rect 194428 480 194456 3402
rect 195612 604 195664 610
rect 195612 546 195664 552
rect 195624 480 195652 546
rect 196820 480 196848 4082
rect 198660 2990 198688 57190
rect 198844 3942 198872 60030
rect 199672 56778 199700 60030
rect 200028 57316 200080 57322
rect 200028 57258 200080 57264
rect 199660 56772 199712 56778
rect 199660 56714 199712 56720
rect 200040 4146 200068 57258
rect 201052 56914 201080 60044
rect 201512 60030 201986 60058
rect 201040 56908 201092 56914
rect 201040 56850 201092 56856
rect 201408 56908 201460 56914
rect 201408 56850 201460 56856
rect 199200 4140 199252 4146
rect 199200 4082 199252 4088
rect 200028 4140 200080 4146
rect 200028 4082 200080 4088
rect 198832 3936 198884 3942
rect 198832 3878 198884 3884
rect 198004 2984 198056 2990
rect 198004 2926 198056 2932
rect 198648 2984 198700 2990
rect 198648 2926 198700 2932
rect 198016 480 198044 2926
rect 199212 480 199240 4082
rect 201420 3398 201448 56850
rect 201512 4298 201540 60030
rect 202984 57390 203012 60044
rect 203996 57662 204024 60044
rect 204272 60030 204930 60058
rect 203984 57656 204036 57662
rect 203984 57598 204036 57604
rect 204168 57656 204220 57662
rect 204168 57598 204220 57604
rect 202972 57384 203024 57390
rect 202972 57326 203024 57332
rect 202786 57216 202842 57225
rect 202786 57151 202842 57160
rect 202696 56976 202748 56982
rect 202696 56918 202748 56924
rect 201512 4270 201724 4298
rect 201500 4140 201552 4146
rect 201500 4082 201552 4088
rect 200396 3392 200448 3398
rect 200396 3334 200448 3340
rect 201408 3392 201460 3398
rect 201408 3334 201460 3340
rect 200408 480 200436 3334
rect 201512 480 201540 4082
rect 201696 3806 201724 4270
rect 202708 4146 202736 56918
rect 202696 4140 202748 4146
rect 202696 4082 202748 4088
rect 202800 4026 202828 57151
rect 204180 13190 204208 57598
rect 203708 13184 203760 13190
rect 203708 13126 203760 13132
rect 204168 13184 204220 13190
rect 204168 13126 204220 13132
rect 202708 3998 202828 4026
rect 201684 3800 201736 3806
rect 201684 3742 201736 3748
rect 202708 480 202736 3998
rect 203720 610 203748 13126
rect 204272 3738 204300 60030
rect 205928 57458 205956 60044
rect 205916 57452 205968 57458
rect 205916 57394 205968 57400
rect 206744 57452 206796 57458
rect 206744 57394 206796 57400
rect 205548 57384 205600 57390
rect 205548 57326 205600 57332
rect 205560 4146 205588 57326
rect 206756 54210 206784 57394
rect 206940 56710 206968 60044
rect 207032 60030 207874 60058
rect 206928 56704 206980 56710
rect 206928 56646 206980 56652
rect 206756 54182 206968 54210
rect 205088 4140 205140 4146
rect 205088 4082 205140 4088
rect 205548 4140 205600 4146
rect 205548 4082 205600 4088
rect 204260 3732 204312 3738
rect 204260 3674 204312 3680
rect 203708 604 203760 610
rect 203708 546 203760 552
rect 203892 604 203944 610
rect 203892 546 203944 552
rect 203904 480 203932 546
rect 205100 480 205128 4082
rect 206940 3126 206968 54182
rect 207032 3874 207060 60030
rect 208872 57594 208900 60044
rect 209792 57730 209820 60044
rect 209884 60030 210818 60058
rect 209780 57724 209832 57730
rect 209780 57666 209832 57672
rect 208860 57588 208912 57594
rect 208860 57530 208912 57536
rect 209688 56840 209740 56846
rect 209688 56782 209740 56788
rect 208308 56704 208360 56710
rect 208308 56646 208360 56652
rect 208320 4146 208348 56646
rect 209700 4146 209728 56782
rect 207480 4140 207532 4146
rect 207480 4082 207532 4088
rect 208308 4140 208360 4146
rect 208308 4082 208360 4088
rect 208676 4140 208728 4146
rect 208676 4082 208728 4088
rect 209688 4140 209740 4146
rect 209688 4082 209740 4088
rect 207020 3868 207072 3874
rect 207020 3810 207072 3816
rect 206284 3120 206336 3126
rect 206284 3062 206336 3068
rect 206928 3120 206980 3126
rect 206928 3062 206980 3068
rect 206296 480 206324 3062
rect 207492 480 207520 4082
rect 208688 480 208716 4082
rect 209884 4010 209912 60030
rect 211068 57588 211120 57594
rect 211068 57530 211120 57536
rect 210976 56636 211028 56642
rect 210976 56578 211028 56584
rect 209872 4004 209924 4010
rect 209872 3946 209924 3952
rect 210988 2990 211016 56578
rect 209872 2984 209924 2990
rect 209872 2926 209924 2932
rect 210976 2984 211028 2990
rect 210976 2926 211028 2932
rect 209884 480 209912 2926
rect 211080 480 211108 57530
rect 211816 57526 211844 60044
rect 212736 57798 212764 60044
rect 213472 60030 213762 60058
rect 212724 57792 212776 57798
rect 212724 57734 212776 57740
rect 211804 57520 211856 57526
rect 211804 57462 211856 57468
rect 212448 56772 212500 56778
rect 212448 56714 212500 56720
rect 212460 9654 212488 56714
rect 213472 48346 213500 60030
rect 214760 57866 214788 60044
rect 215680 57934 215708 60044
rect 215668 57928 215720 57934
rect 215668 57870 215720 57876
rect 214748 57860 214800 57866
rect 214748 57802 214800 57808
rect 215208 57860 215260 57866
rect 215208 57802 215260 57808
rect 213828 57724 213880 57730
rect 213828 57666 213880 57672
rect 212632 48340 212684 48346
rect 212632 48282 212684 48288
rect 213460 48340 213512 48346
rect 213460 48282 213512 48288
rect 212644 41426 212672 48282
rect 212552 41410 212672 41426
rect 212540 41404 212672 41410
rect 212592 41398 212672 41404
rect 212724 41404 212776 41410
rect 212540 41346 212592 41352
rect 212724 41346 212776 41352
rect 212736 33810 212764 41346
rect 212552 33782 212764 33810
rect 212552 27606 212580 33782
rect 212540 27600 212592 27606
rect 212540 27542 212592 27548
rect 212632 18012 212684 18018
rect 212632 17954 212684 17960
rect 212644 12458 212672 17954
rect 212644 12430 212764 12458
rect 212448 9648 212500 9654
rect 212448 9590 212500 9596
rect 212736 3670 212764 12430
rect 212724 3664 212776 3670
rect 212724 3606 212776 3612
rect 213840 2854 213868 57666
rect 215220 4146 215248 57802
rect 216588 56636 216640 56642
rect 216588 56578 216640 56584
rect 214656 4140 214708 4146
rect 214656 4082 214708 4088
rect 215208 4140 215260 4146
rect 215208 4082 215260 4088
rect 213828 2848 213880 2854
rect 213828 2790 213880 2796
rect 212264 604 212316 610
rect 212264 546 212316 552
rect 213460 604 213512 610
rect 213460 546 213512 552
rect 212276 480 212304 546
rect 213472 480 213500 546
rect 214668 480 214696 4082
rect 216600 3534 216628 56578
rect 216692 3942 216720 60044
rect 217704 57118 217732 60044
rect 218624 57526 218652 60044
rect 219544 60030 219650 60058
rect 218612 57520 218664 57526
rect 218612 57462 218664 57468
rect 219256 57520 219308 57526
rect 219256 57462 219308 57468
rect 217692 57112 217744 57118
rect 217692 57054 217744 57060
rect 217968 57044 218020 57050
rect 217968 56986 218020 56992
rect 216680 3936 216732 3942
rect 216680 3878 216732 3884
rect 217980 3534 218008 56986
rect 218152 3596 218204 3602
rect 218152 3538 218204 3544
rect 215852 3528 215904 3534
rect 215852 3470 215904 3476
rect 216588 3528 216640 3534
rect 216588 3470 216640 3476
rect 217048 3528 217100 3534
rect 217048 3470 217100 3476
rect 217968 3528 218020 3534
rect 217968 3470 218020 3476
rect 215864 480 215892 3470
rect 217060 480 217088 3470
rect 218164 480 218192 3538
rect 219268 3482 219296 57462
rect 219348 57112 219400 57118
rect 219348 57054 219400 57060
rect 219360 3602 219388 57054
rect 219348 3596 219400 3602
rect 219348 3538 219400 3544
rect 219268 3454 219388 3482
rect 219544 3466 219572 60030
rect 220648 57186 220676 60044
rect 221568 57798 221596 60044
rect 221556 57792 221608 57798
rect 221556 57734 221608 57740
rect 222108 57792 222160 57798
rect 222108 57734 222160 57740
rect 220636 57180 220688 57186
rect 220636 57122 220688 57128
rect 220728 57180 220780 57186
rect 220728 57122 220780 57128
rect 220740 3482 220768 57122
rect 222120 3482 222148 57734
rect 222580 57254 222608 60044
rect 223592 57322 223620 60044
rect 223580 57316 223632 57322
rect 223580 57258 223632 57264
rect 222568 57248 222620 57254
rect 222568 57190 222620 57196
rect 223488 57248 223540 57254
rect 223488 57190 223540 57196
rect 223500 3534 223528 57190
rect 224512 56914 224540 60044
rect 225524 56982 225552 60044
rect 226444 57225 226472 60044
rect 227456 57662 227484 60044
rect 227444 57656 227496 57662
rect 227444 57598 227496 57604
rect 228468 57390 228496 60044
rect 229008 57656 229060 57662
rect 229008 57598 229060 57604
rect 228456 57384 228508 57390
rect 228456 57326 228508 57332
rect 228916 57316 228968 57322
rect 228916 57258 228968 57264
rect 226430 57216 226486 57225
rect 226430 57151 226486 57160
rect 225512 56976 225564 56982
rect 225512 56918 225564 56924
rect 227628 56976 227680 56982
rect 227628 56918 227680 56924
rect 224500 56908 224552 56914
rect 224500 56850 224552 56856
rect 224868 56908 224920 56914
rect 224868 56850 224920 56856
rect 219360 480 219388 3454
rect 219532 3460 219584 3466
rect 219532 3402 219584 3408
rect 220556 3454 220768 3482
rect 221752 3454 222148 3482
rect 222936 3528 222988 3534
rect 222936 3470 222988 3476
rect 223488 3528 223540 3534
rect 223488 3470 223540 3476
rect 220556 480 220584 3454
rect 221752 480 221780 3454
rect 222948 480 222976 3470
rect 224880 3058 224908 56850
rect 226248 56704 226300 56710
rect 226248 56646 226300 56652
rect 226260 3534 226288 56646
rect 227640 3534 227668 56918
rect 225328 3528 225380 3534
rect 225328 3470 225380 3476
rect 226248 3528 226300 3534
rect 226248 3470 226300 3476
rect 226524 3528 226576 3534
rect 226524 3470 226576 3476
rect 227628 3528 227680 3534
rect 227628 3470 227680 3476
rect 224132 3052 224184 3058
rect 224132 2994 224184 3000
rect 224868 3052 224920 3058
rect 224868 2994 224920 3000
rect 224144 480 224172 2994
rect 225340 480 225368 3470
rect 226536 480 226564 3470
rect 227720 3460 227772 3466
rect 227720 3402 227772 3408
rect 227732 480 227760 3402
rect 228928 480 228956 57258
rect 229020 3466 229048 57598
rect 229388 57458 229416 60044
rect 229376 57452 229428 57458
rect 229376 57394 229428 57400
rect 230400 57390 230428 60044
rect 230480 57452 230532 57458
rect 230480 57394 230532 57400
rect 230388 57384 230440 57390
rect 230388 57326 230440 57332
rect 230492 57202 230520 57394
rect 230400 57174 230520 57202
rect 230400 3482 230428 57174
rect 231412 56846 231440 60044
rect 232332 57730 232360 60044
rect 232320 57724 232372 57730
rect 232320 57666 232372 57672
rect 233148 57724 233200 57730
rect 233148 57666 233200 57672
rect 231768 57384 231820 57390
rect 231768 57326 231820 57332
rect 231400 56840 231452 56846
rect 231400 56782 231452 56788
rect 231780 3534 231808 57326
rect 233160 3534 233188 57666
rect 233344 57594 233372 60044
rect 233332 57588 233384 57594
rect 233332 57530 233384 57536
rect 234356 56778 234384 60044
rect 235276 57798 235304 60044
rect 236288 57866 236316 60044
rect 237024 60030 237314 60058
rect 236276 57860 236328 57866
rect 236276 57802 236328 57808
rect 235264 57792 235316 57798
rect 235264 57734 235316 57740
rect 234528 56840 234580 56846
rect 234528 56782 234580 56788
rect 234344 56772 234396 56778
rect 234344 56714 234396 56720
rect 234540 3534 234568 56782
rect 235908 56772 235960 56778
rect 235908 56714 235960 56720
rect 229008 3460 229060 3466
rect 229008 3402 229060 3408
rect 230124 3454 230428 3482
rect 231308 3528 231360 3534
rect 231308 3470 231360 3476
rect 231768 3528 231820 3534
rect 231768 3470 231820 3476
rect 232504 3528 232556 3534
rect 232504 3470 232556 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 233700 3528 233752 3534
rect 233700 3470 233752 3476
rect 234528 3528 234580 3534
rect 234528 3470 234580 3476
rect 230124 480 230152 3454
rect 231320 480 231348 3470
rect 232516 480 232544 3470
rect 233712 480 233740 3470
rect 235920 3330 235948 56714
rect 237024 56642 237052 60030
rect 237288 57792 237340 57798
rect 237288 57734 237340 57740
rect 237196 57588 237248 57594
rect 237196 57530 237248 57536
rect 237012 56636 237064 56642
rect 237012 56578 237064 56584
rect 234804 3324 234856 3330
rect 234804 3266 234856 3272
rect 235908 3324 235960 3330
rect 235908 3266 235960 3272
rect 234816 480 234844 3266
rect 236000 3256 236052 3262
rect 236000 3198 236052 3204
rect 236012 480 236040 3198
rect 237208 480 237236 57530
rect 237300 3262 237328 57734
rect 238220 57050 238248 60044
rect 239232 57118 239260 60044
rect 240048 57860 240100 57866
rect 240048 57802 240100 57808
rect 239220 57112 239272 57118
rect 239220 57054 239272 57060
rect 238208 57044 238260 57050
rect 238208 56986 238260 56992
rect 238668 57044 238720 57050
rect 238668 56986 238720 56992
rect 238680 3482 238708 56986
rect 240060 3534 240088 57802
rect 240244 57526 240272 60044
rect 240232 57520 240284 57526
rect 240232 57462 240284 57468
rect 241164 57186 241192 60044
rect 242176 57934 242204 60044
rect 242164 57928 242216 57934
rect 242164 57870 242216 57876
rect 241428 57520 241480 57526
rect 241428 57462 241480 57468
rect 241152 57180 241204 57186
rect 241152 57122 241204 57128
rect 241440 3534 241468 57462
rect 243096 57254 243124 60044
rect 243084 57248 243136 57254
rect 243084 57190 243136 57196
rect 242808 57112 242860 57118
rect 242808 57054 242860 57060
rect 238404 3454 238708 3482
rect 239588 3528 239640 3534
rect 239588 3470 239640 3476
rect 240048 3528 240100 3534
rect 240048 3470 240100 3476
rect 240784 3528 240836 3534
rect 240784 3470 240836 3476
rect 241428 3528 241480 3534
rect 241428 3470 241480 3476
rect 237288 3256 237340 3262
rect 237288 3198 237340 3204
rect 238404 480 238432 3454
rect 239600 480 239628 3470
rect 240796 480 240824 3470
rect 242820 3466 242848 57054
rect 244108 56914 244136 60044
rect 244188 57248 244240 57254
rect 244188 57190 244240 57196
rect 244096 56908 244148 56914
rect 244096 56850 244148 56856
rect 244200 3534 244228 57190
rect 245120 56710 245148 60044
rect 245568 57928 245620 57934
rect 245568 57870 245620 57876
rect 245476 56908 245528 56914
rect 245476 56850 245528 56856
rect 245108 56704 245160 56710
rect 245108 56646 245160 56652
rect 245488 3534 245516 56850
rect 243176 3528 243228 3534
rect 243176 3470 243228 3476
rect 244188 3528 244240 3534
rect 244188 3470 244240 3476
rect 244372 3528 244424 3534
rect 244372 3470 244424 3476
rect 245476 3528 245528 3534
rect 245476 3470 245528 3476
rect 241980 3460 242032 3466
rect 241980 3402 242032 3408
rect 242808 3460 242860 3466
rect 242808 3402 242860 3408
rect 241992 480 242020 3402
rect 243188 480 243216 3470
rect 244384 480 244412 3470
rect 245580 480 245608 57870
rect 246040 56982 246068 60044
rect 247052 57662 247080 60044
rect 247040 57656 247092 57662
rect 247040 57598 247092 57604
rect 248064 57322 248092 60044
rect 248984 57458 249012 60044
rect 248972 57452 249024 57458
rect 248972 57394 249024 57400
rect 249996 57390 250024 60044
rect 251008 57730 251036 60044
rect 250996 57724 251048 57730
rect 250996 57666 251048 57672
rect 251088 57452 251140 57458
rect 251088 57394 251140 57400
rect 249984 57384 250036 57390
rect 249984 57326 250036 57332
rect 248052 57316 248104 57322
rect 248052 57258 248104 57264
rect 248328 57316 248380 57322
rect 248328 57258 248380 57264
rect 246948 57180 247000 57186
rect 246948 57122 247000 57128
rect 246028 56976 246080 56982
rect 246028 56918 246080 56924
rect 246960 3482 246988 57122
rect 248340 3482 248368 57258
rect 249708 56976 249760 56982
rect 249708 56918 249760 56924
rect 249720 3534 249748 56918
rect 251100 3534 251128 57394
rect 251928 56846 251956 60044
rect 252468 57656 252520 57662
rect 252468 57598 252520 57604
rect 251916 56840 251968 56846
rect 251916 56782 251968 56788
rect 252480 3534 252508 57598
rect 252940 56778 252968 60044
rect 253952 57798 253980 60044
rect 253940 57792 253992 57798
rect 253940 57734 253992 57740
rect 254872 57594 254900 60044
rect 255228 57724 255280 57730
rect 255228 57666 255280 57672
rect 254860 57588 254912 57594
rect 254860 57530 254912 57536
rect 253756 57384 253808 57390
rect 253756 57326 253808 57332
rect 252928 56772 252980 56778
rect 252928 56714 252980 56720
rect 252652 3596 252704 3602
rect 252652 3538 252704 3544
rect 246776 3454 246988 3482
rect 247972 3454 248368 3482
rect 249156 3528 249208 3534
rect 249156 3470 249208 3476
rect 249708 3528 249760 3534
rect 249708 3470 249760 3476
rect 250352 3528 250404 3534
rect 250352 3470 250404 3476
rect 251088 3528 251140 3534
rect 251088 3470 251140 3476
rect 251456 3528 251508 3534
rect 251456 3470 251508 3476
rect 252468 3528 252520 3534
rect 252468 3470 252520 3476
rect 246776 480 246804 3454
rect 247972 480 248000 3454
rect 249168 480 249196 3470
rect 250364 480 250392 3470
rect 251468 480 251496 3470
rect 252664 480 252692 3538
rect 253768 3482 253796 57326
rect 253848 56840 253900 56846
rect 253848 56782 253900 56788
rect 253860 3602 253888 56782
rect 253848 3596 253900 3602
rect 253848 3538 253900 3544
rect 255240 3482 255268 57666
rect 255884 57050 255912 60044
rect 256896 57866 256924 60044
rect 256884 57860 256936 57866
rect 256884 57802 256936 57808
rect 256608 57588 256660 57594
rect 256608 57530 256660 57536
rect 255872 57044 255924 57050
rect 255872 56986 255924 56992
rect 256620 3482 256648 57530
rect 257816 57526 257844 60044
rect 257988 57792 258040 57798
rect 257988 57734 258040 57740
rect 257804 57520 257856 57526
rect 257804 57462 257856 57468
rect 258000 3534 258028 57734
rect 258828 57118 258856 60044
rect 259368 57860 259420 57866
rect 259368 57802 259420 57808
rect 258816 57112 258868 57118
rect 258816 57054 258868 57060
rect 253768 3454 253888 3482
rect 253860 480 253888 3454
rect 255056 3454 255268 3482
rect 256252 3454 256648 3482
rect 257436 3528 257488 3534
rect 257436 3470 257488 3476
rect 257988 3528 258040 3534
rect 257988 3470 258040 3476
rect 255056 480 255084 3454
rect 256252 480 256280 3454
rect 257448 480 257476 3470
rect 259380 3126 259408 57802
rect 259748 57254 259776 60044
rect 260392 60030 260774 60058
rect 259736 57248 259788 57254
rect 259736 57190 259788 57196
rect 260392 56914 260420 60030
rect 261772 57934 261800 60044
rect 261760 57928 261812 57934
rect 261760 57870 261812 57876
rect 260748 57520 260800 57526
rect 260748 57462 260800 57468
rect 260380 56908 260432 56914
rect 260380 56850 260432 56856
rect 260760 3534 260788 57462
rect 262692 57186 262720 60044
rect 263508 57928 263560 57934
rect 263508 57870 263560 57876
rect 263416 57248 263468 57254
rect 263416 57190 263468 57196
rect 262680 57180 262732 57186
rect 262680 57122 262732 57128
rect 262128 57112 262180 57118
rect 262128 57054 262180 57060
rect 259828 3528 259880 3534
rect 259828 3470 259880 3476
rect 260748 3528 260800 3534
rect 260748 3470 260800 3476
rect 258632 3120 258684 3126
rect 258632 3062 258684 3068
rect 259368 3120 259420 3126
rect 259368 3062 259420 3068
rect 258644 480 258672 3062
rect 259840 480 259868 3470
rect 262140 3262 262168 57054
rect 262220 3528 262272 3534
rect 262220 3470 262272 3476
rect 261024 3256 261076 3262
rect 261024 3198 261076 3204
rect 262128 3256 262180 3262
rect 262128 3198 262180 3204
rect 261036 480 261064 3198
rect 262232 480 262260 3470
rect 263428 480 263456 57190
rect 263520 3534 263548 57870
rect 263704 57322 263732 60044
rect 263692 57316 263744 57322
rect 263692 57258 263744 57264
rect 264716 56982 264744 60044
rect 265636 57458 265664 60044
rect 266648 57662 266676 60044
rect 267384 60030 267674 60058
rect 266636 57656 266688 57662
rect 266636 57598 266688 57604
rect 265624 57452 265676 57458
rect 265624 57394 265676 57400
rect 266268 57452 266320 57458
rect 266268 57394 266320 57400
rect 264888 57316 264940 57322
rect 264888 57258 264940 57264
rect 264704 56976 264756 56982
rect 264704 56918 264756 56924
rect 263508 3528 263560 3534
rect 264900 3482 264928 57258
rect 266280 3534 266308 57394
rect 267384 56846 267412 60030
rect 267648 57656 267700 57662
rect 267648 57598 267700 57604
rect 267372 56840 267424 56846
rect 267372 56782 267424 56788
rect 263508 3470 263560 3476
rect 264624 3454 264928 3482
rect 265808 3528 265860 3534
rect 265808 3470 265860 3476
rect 266268 3528 266320 3534
rect 266268 3470 266320 3476
rect 264624 480 264652 3454
rect 265820 480 265848 3470
rect 267660 3466 267688 57598
rect 268580 57390 268608 60044
rect 269592 57730 269620 60044
rect 269580 57724 269632 57730
rect 269580 57666 269632 57672
rect 270604 57594 270632 60044
rect 271524 57798 271552 60044
rect 272536 57866 272564 60044
rect 272524 57860 272576 57866
rect 272524 57802 272576 57808
rect 271512 57792 271564 57798
rect 271512 57734 271564 57740
rect 271696 57724 271748 57730
rect 271696 57666 271748 57672
rect 270592 57588 270644 57594
rect 270592 57530 270644 57536
rect 268568 57384 268620 57390
rect 268568 57326 268620 57332
rect 269028 57180 269080 57186
rect 269028 57122 269080 57128
rect 267004 3460 267056 3466
rect 267004 3402 267056 3408
rect 267648 3460 267700 3466
rect 267648 3402 267700 3408
rect 267016 480 267044 3402
rect 269040 3058 269068 57122
rect 270408 57044 270460 57050
rect 270408 56986 270460 56992
rect 270420 3534 270448 56986
rect 271708 3602 271736 57666
rect 273168 57588 273220 57594
rect 273168 57530 273220 57536
rect 271788 57384 271840 57390
rect 271788 57326 271840 57332
rect 270500 3596 270552 3602
rect 270500 3538 270552 3544
rect 271696 3596 271748 3602
rect 271696 3538 271748 3544
rect 269304 3528 269356 3534
rect 269304 3470 269356 3476
rect 270408 3528 270460 3534
rect 270408 3470 270460 3476
rect 268108 3052 268160 3058
rect 268108 2994 268160 3000
rect 269028 3052 269080 3058
rect 269028 2994 269080 3000
rect 268120 480 268148 2994
rect 269316 480 269344 3470
rect 270512 480 270540 3538
rect 271800 3482 271828 57326
rect 273180 3482 273208 57530
rect 273548 57526 273576 60044
rect 273536 57520 273588 57526
rect 273536 57462 273588 57468
rect 274468 57118 274496 60044
rect 275480 57934 275508 60044
rect 275468 57928 275520 57934
rect 275468 57870 275520 57876
rect 274548 57860 274600 57866
rect 274548 57802 274600 57808
rect 274456 57112 274508 57118
rect 274456 57054 274508 57060
rect 274560 3534 274588 57802
rect 275928 57792 275980 57798
rect 275928 57734 275980 57740
rect 275940 3534 275968 57734
rect 276400 57254 276428 60044
rect 277308 57520 277360 57526
rect 277308 57462 277360 57468
rect 276388 57248 276440 57254
rect 276388 57190 276440 57196
rect 277320 3534 277348 57462
rect 277412 57322 277440 60044
rect 278424 57458 278452 60044
rect 279344 57662 279372 60044
rect 280068 57928 280120 57934
rect 280068 57870 280120 57876
rect 279332 57656 279384 57662
rect 279332 57598 279384 57604
rect 278412 57452 278464 57458
rect 278412 57394 278464 57400
rect 277400 57316 277452 57322
rect 277400 57258 277452 57264
rect 278688 57316 278740 57322
rect 278688 57258 278740 57264
rect 278700 3534 278728 57258
rect 279976 57248 280028 57254
rect 279976 57190 280028 57196
rect 278872 3596 278924 3602
rect 278872 3538 278924 3544
rect 271708 3454 271828 3482
rect 272904 3454 273208 3482
rect 274088 3528 274140 3534
rect 274088 3470 274140 3476
rect 274548 3528 274600 3534
rect 274548 3470 274600 3476
rect 275284 3528 275336 3534
rect 275284 3470 275336 3476
rect 275928 3528 275980 3534
rect 275928 3470 275980 3476
rect 276480 3528 276532 3534
rect 276480 3470 276532 3476
rect 277308 3528 277360 3534
rect 277308 3470 277360 3476
rect 277676 3528 277728 3534
rect 277676 3470 277728 3476
rect 278688 3528 278740 3534
rect 278688 3470 278740 3476
rect 271708 480 271736 3454
rect 272904 480 272932 3454
rect 274100 480 274128 3470
rect 275296 480 275324 3470
rect 276492 480 276520 3470
rect 277688 480 277716 3470
rect 278884 480 278912 3538
rect 279988 3482 280016 57190
rect 280080 3602 280108 57870
rect 280356 57186 280384 60044
rect 280344 57180 280396 57186
rect 280344 57122 280396 57128
rect 281368 57050 281396 60044
rect 282288 57730 282316 60044
rect 282276 57724 282328 57730
rect 282276 57666 282328 57672
rect 281448 57656 281500 57662
rect 281448 57598 281500 57604
rect 281356 57044 281408 57050
rect 281356 56986 281408 56992
rect 280068 3596 280120 3602
rect 280068 3538 280120 3544
rect 281460 3516 281488 57598
rect 282828 57452 282880 57458
rect 282828 57394 282880 57400
rect 282840 3516 282868 57394
rect 283300 57390 283328 60044
rect 284208 57724 284260 57730
rect 284208 57666 284260 57672
rect 283288 57384 283340 57390
rect 283288 57326 283340 57332
rect 284220 3534 284248 57666
rect 284312 57594 284340 60044
rect 285232 57866 285260 60044
rect 285220 57860 285272 57866
rect 285220 57802 285272 57808
rect 286244 57798 286272 60044
rect 286232 57792 286284 57798
rect 286232 57734 286284 57740
rect 284300 57588 284352 57594
rect 284300 57530 284352 57536
rect 286968 57588 287020 57594
rect 286968 57530 287020 57536
rect 285588 57384 285640 57390
rect 285588 57326 285640 57332
rect 285600 3534 285628 57326
rect 286980 3534 287008 57530
rect 287256 57526 287284 60044
rect 287244 57520 287296 57526
rect 287244 57462 287296 57468
rect 288176 57322 288204 60044
rect 289188 57934 289216 60044
rect 289176 57928 289228 57934
rect 289176 57870 289228 57876
rect 289728 57520 289780 57526
rect 289728 57462 289780 57468
rect 288164 57316 288216 57322
rect 288164 57258 288216 57264
rect 288256 57316 288308 57322
rect 288256 57258 288308 57264
rect 287152 3596 287204 3602
rect 287152 3538 287204 3544
rect 281276 3488 281488 3516
rect 282472 3488 282868 3516
rect 283656 3528 283708 3534
rect 279988 3454 280108 3482
rect 280080 480 280108 3454
rect 281276 480 281304 3488
rect 282472 480 282500 3488
rect 283656 3470 283708 3476
rect 284208 3528 284260 3534
rect 284208 3470 284260 3476
rect 284760 3528 284812 3534
rect 284760 3470 284812 3476
rect 285588 3528 285640 3534
rect 285588 3470 285640 3476
rect 285956 3528 286008 3534
rect 285956 3470 286008 3476
rect 286968 3528 287020 3534
rect 286968 3470 287020 3476
rect 283668 480 283696 3470
rect 284772 480 284800 3470
rect 285968 480 285996 3470
rect 287164 480 287192 3538
rect 288268 3482 288296 57258
rect 288348 56976 288400 56982
rect 288348 56918 288400 56924
rect 288360 3602 288388 56918
rect 288348 3596 288400 3602
rect 288348 3538 288400 3544
rect 289740 3482 289768 57462
rect 290200 57254 290228 60044
rect 291120 57662 291148 60044
rect 291108 57656 291160 57662
rect 291108 57598 291160 57604
rect 292132 57458 292160 60044
rect 293052 57730 293080 60044
rect 293040 57724 293092 57730
rect 293040 57666 293092 57672
rect 292120 57452 292172 57458
rect 292120 57394 292172 57400
rect 292488 57452 292540 57458
rect 292488 57394 292540 57400
rect 290188 57248 290240 57254
rect 290188 57190 290240 57196
rect 291108 56636 291160 56642
rect 291108 56578 291160 56584
rect 291120 3482 291148 56578
rect 292500 3534 292528 57394
rect 294064 57390 294092 60044
rect 295076 57594 295104 60044
rect 295064 57588 295116 57594
rect 295064 57530 295116 57536
rect 294052 57384 294104 57390
rect 294052 57326 294104 57332
rect 295248 57384 295300 57390
rect 295248 57326 295300 57332
rect 293868 57248 293920 57254
rect 293868 57190 293920 57196
rect 293880 3534 293908 57190
rect 295260 3534 295288 57326
rect 295996 56982 296024 60044
rect 296628 57724 296680 57730
rect 296628 57666 296680 57672
rect 295984 56976 296036 56982
rect 295984 56918 296036 56924
rect 296640 3534 296668 57666
rect 297008 57322 297036 60044
rect 298020 57526 298048 60044
rect 298008 57520 298060 57526
rect 298008 57462 298060 57468
rect 296996 57316 297048 57322
rect 296996 57258 297048 57264
rect 298008 57316 298060 57322
rect 298008 57258 298060 57264
rect 297916 57112 297968 57118
rect 297916 57054 297968 57060
rect 297928 3602 297956 57054
rect 296720 3596 296772 3602
rect 296720 3538 296772 3544
rect 297916 3596 297968 3602
rect 297916 3538 297968 3544
rect 288268 3454 288388 3482
rect 288360 480 288388 3454
rect 289556 3454 289768 3482
rect 290752 3454 291148 3482
rect 291936 3528 291988 3534
rect 291936 3470 291988 3476
rect 292488 3528 292540 3534
rect 292488 3470 292540 3476
rect 293132 3528 293184 3534
rect 293132 3470 293184 3476
rect 293868 3528 293920 3534
rect 293868 3470 293920 3476
rect 294328 3528 294380 3534
rect 294328 3470 294380 3476
rect 295248 3528 295300 3534
rect 295248 3470 295300 3476
rect 295524 3528 295576 3534
rect 295524 3470 295576 3476
rect 296628 3528 296680 3534
rect 296628 3470 296680 3476
rect 289556 480 289584 3454
rect 290752 480 290780 3454
rect 291948 480 291976 3470
rect 293144 480 293172 3470
rect 294340 480 294368 3470
rect 295536 480 295564 3470
rect 296732 480 296760 3538
rect 298020 3482 298048 57258
rect 298940 56642 298968 60044
rect 299388 57520 299440 57526
rect 299388 57462 299440 57468
rect 298928 56636 298980 56642
rect 298928 56578 298980 56584
rect 299400 3482 299428 57462
rect 299952 57458 299980 60044
rect 299940 57452 299992 57458
rect 299940 57394 299992 57400
rect 300964 57254 300992 60044
rect 301884 57390 301912 60044
rect 302896 57730 302924 60044
rect 302884 57724 302936 57730
rect 302884 57666 302936 57672
rect 301872 57384 301924 57390
rect 301872 57326 301924 57332
rect 300952 57248 301004 57254
rect 300952 57190 301004 57196
rect 303908 57118 303936 60044
rect 304828 57322 304856 60044
rect 305840 57526 305868 60044
rect 305828 57520 305880 57526
rect 305828 57462 305880 57468
rect 306288 57520 306340 57526
rect 306288 57462 306340 57468
rect 304908 57384 304960 57390
rect 304908 57326 304960 57332
rect 304816 57316 304868 57322
rect 304816 57258 304868 57264
rect 303896 57112 303948 57118
rect 303896 57054 303948 57060
rect 302148 56772 302200 56778
rect 302148 56714 302200 56720
rect 302160 3534 302188 56714
rect 303528 56704 303580 56710
rect 303528 56646 303580 56652
rect 303540 3534 303568 56646
rect 304264 56636 304316 56642
rect 304264 56578 304316 56584
rect 297928 3454 298048 3482
rect 299124 3454 299428 3482
rect 301412 3528 301464 3534
rect 301412 3470 301464 3476
rect 302148 3528 302200 3534
rect 302148 3470 302200 3476
rect 302608 3528 302660 3534
rect 302608 3470 302660 3476
rect 303528 3528 303580 3534
rect 303528 3470 303580 3476
rect 303804 3528 303856 3534
rect 303804 3470 303856 3476
rect 297928 480 297956 3454
rect 299124 480 299152 3454
rect 300308 3324 300360 3330
rect 300308 3266 300360 3272
rect 300320 480 300348 3266
rect 301424 480 301452 3470
rect 302620 480 302648 3470
rect 303816 480 303844 3470
rect 304276 3330 304304 56578
rect 304920 3534 304948 57326
rect 306196 57316 306248 57322
rect 306196 57258 306248 57264
rect 306208 3602 306236 57258
rect 305000 3596 305052 3602
rect 305000 3538 305052 3544
rect 306196 3596 306248 3602
rect 306196 3538 306248 3544
rect 304908 3528 304960 3534
rect 304908 3470 304960 3476
rect 304264 3324 304316 3330
rect 304264 3266 304316 3272
rect 305012 480 305040 3538
rect 306300 3482 306328 57462
rect 306852 56642 306880 60044
rect 307668 56908 307720 56914
rect 307668 56850 307720 56856
rect 306840 56636 306892 56642
rect 306840 56578 306892 56584
rect 307680 3482 307708 56850
rect 307772 56778 307800 60044
rect 307760 56772 307812 56778
rect 307760 56714 307812 56720
rect 308784 56710 308812 60044
rect 309048 57588 309100 57594
rect 309048 57530 309100 57536
rect 308772 56704 308824 56710
rect 308772 56646 308824 56652
rect 309060 3534 309088 57530
rect 309704 57390 309732 60044
rect 310428 57724 310480 57730
rect 310428 57666 310480 57672
rect 309692 57384 309744 57390
rect 309692 57326 309744 57332
rect 310440 3534 310468 57666
rect 310716 57322 310744 60044
rect 311728 57526 311756 60044
rect 311808 57656 311860 57662
rect 311808 57598 311860 57604
rect 311716 57520 311768 57526
rect 311716 57462 311768 57468
rect 310704 57316 310756 57322
rect 310704 57258 310756 57264
rect 311820 3534 311848 57598
rect 312648 56914 312676 60044
rect 313660 57594 313688 60044
rect 314672 57730 314700 60044
rect 314660 57724 314712 57730
rect 314660 57666 314712 57672
rect 315592 57662 315620 60044
rect 315580 57656 315632 57662
rect 315580 57598 315632 57604
rect 313648 57588 313700 57594
rect 313648 57530 313700 57536
rect 315948 57248 316000 57254
rect 315948 57190 316000 57196
rect 312636 56908 312688 56914
rect 312636 56850 312688 56856
rect 313188 56772 313240 56778
rect 313188 56714 313240 56720
rect 313200 3534 313228 56714
rect 315304 56704 315356 56710
rect 315304 56646 315356 56652
rect 313372 4004 313424 4010
rect 313372 3946 313424 3952
rect 306208 3454 306328 3482
rect 307404 3454 307708 3482
rect 308588 3528 308640 3534
rect 308588 3470 308640 3476
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 309784 3528 309836 3534
rect 309784 3470 309836 3476
rect 310428 3528 310480 3534
rect 310428 3470 310480 3476
rect 310980 3528 311032 3534
rect 310980 3470 311032 3476
rect 311808 3528 311860 3534
rect 311808 3470 311860 3476
rect 312176 3528 312228 3534
rect 312176 3470 312228 3476
rect 313188 3528 313240 3534
rect 313188 3470 313240 3476
rect 306208 480 306236 3454
rect 307404 480 307432 3454
rect 308600 480 308628 3470
rect 309796 480 309824 3470
rect 310992 480 311020 3470
rect 312188 480 312216 3470
rect 313384 480 313412 3946
rect 315316 3534 315344 56646
rect 314568 3528 314620 3534
rect 314568 3470 314620 3476
rect 315304 3528 315356 3534
rect 315960 3482 315988 57190
rect 316604 56778 316632 60044
rect 317616 57662 317644 60044
rect 316684 57656 316736 57662
rect 316684 57598 316736 57604
rect 317604 57656 317656 57662
rect 317604 57598 317656 57604
rect 316592 56772 316644 56778
rect 316592 56714 316644 56720
rect 316696 4010 316724 57598
rect 317328 57588 317380 57594
rect 317328 57530 317380 57536
rect 316684 4004 316736 4010
rect 316684 3946 316736 3952
rect 315304 3470 315356 3476
rect 314580 480 314608 3470
rect 315776 3454 315988 3482
rect 315776 480 315804 3454
rect 317340 610 317368 57530
rect 318536 56710 318564 60044
rect 319444 57860 319496 57866
rect 319444 57802 319496 57808
rect 318524 56704 318576 56710
rect 318524 56646 318576 56652
rect 319456 3534 319484 57802
rect 319548 57254 319576 60044
rect 320560 57594 320588 60044
rect 321480 57866 321508 60044
rect 321468 57860 321520 57866
rect 321468 57802 321520 57808
rect 321468 57724 321520 57730
rect 321468 57666 321520 57672
rect 320548 57588 320600 57594
rect 320548 57530 320600 57536
rect 320088 57520 320140 57526
rect 320088 57462 320140 57468
rect 319536 57248 319588 57254
rect 319536 57190 319588 57196
rect 318064 3528 318116 3534
rect 318064 3470 318116 3476
rect 319444 3528 319496 3534
rect 319444 3470 319496 3476
rect 316960 604 317012 610
rect 316960 546 317012 552
rect 317328 604 317380 610
rect 317328 546 317380 552
rect 316972 480 317000 546
rect 318076 480 318104 3470
rect 320100 3466 320128 57462
rect 321480 3534 321508 57666
rect 322492 57526 322520 60044
rect 323504 57730 323532 60044
rect 323492 57724 323544 57730
rect 323492 57666 323544 57672
rect 322848 57656 322900 57662
rect 322848 57598 322900 57604
rect 322756 57588 322808 57594
rect 322756 57530 322808 57536
rect 322480 57520 322532 57526
rect 322480 57462 322532 57468
rect 322768 3534 322796 57530
rect 320456 3528 320508 3534
rect 320456 3470 320508 3476
rect 321468 3528 321520 3534
rect 321468 3470 321520 3476
rect 321652 3528 321704 3534
rect 321652 3470 321704 3476
rect 322756 3528 322808 3534
rect 322756 3470 322808 3476
rect 319260 3460 319312 3466
rect 319260 3402 319312 3408
rect 320088 3460 320140 3466
rect 320088 3402 320140 3408
rect 319272 480 319300 3402
rect 320468 480 320496 3470
rect 321664 480 321692 3470
rect 322860 480 322888 57598
rect 324424 57594 324452 60044
rect 325436 57662 325464 60044
rect 325424 57656 325476 57662
rect 325424 57598 325476 57604
rect 324412 57588 324464 57594
rect 324412 57530 324464 57536
rect 326356 56710 326384 60044
rect 326988 57792 327040 57798
rect 326988 57734 327040 57740
rect 324228 56704 324280 56710
rect 324228 56646 324280 56652
rect 326344 56704 326396 56710
rect 326344 56646 326396 56652
rect 324240 3482 324268 56646
rect 326344 56568 326396 56574
rect 326344 56510 326396 56516
rect 324056 3454 324268 3482
rect 324056 480 324084 3454
rect 326356 3398 326384 56510
rect 327000 3534 327028 57734
rect 327368 56642 327396 60044
rect 328380 57798 328408 60044
rect 328368 57792 328420 57798
rect 328368 57734 328420 57740
rect 329300 57662 329328 60044
rect 329944 60030 330326 60058
rect 331232 60030 331338 60058
rect 331416 60030 332258 60058
rect 332704 60030 333270 60058
rect 333992 60030 334282 60058
rect 328368 57656 328420 57662
rect 328368 57598 328420 57604
rect 329288 57656 329340 57662
rect 329288 57598 329340 57604
rect 327356 56636 327408 56642
rect 327356 56578 327408 56584
rect 328380 3534 328408 57598
rect 329944 3534 329972 60030
rect 331232 57610 331260 60030
rect 331140 57582 331260 57610
rect 326436 3528 326488 3534
rect 326436 3470 326488 3476
rect 326988 3528 327040 3534
rect 326988 3470 327040 3476
rect 327632 3528 327684 3534
rect 327632 3470 327684 3476
rect 328368 3528 328420 3534
rect 328368 3470 328420 3476
rect 328828 3528 328880 3534
rect 328828 3470 328880 3476
rect 329932 3528 329984 3534
rect 329932 3470 329984 3476
rect 325240 3392 325292 3398
rect 325240 3334 325292 3340
rect 326344 3392 326396 3398
rect 326344 3334 326396 3340
rect 325252 480 325280 3334
rect 326448 480 326476 3470
rect 327644 480 327672 3470
rect 328840 480 328868 3470
rect 331140 3330 331168 57582
rect 330024 3324 330076 3330
rect 330024 3266 330076 3272
rect 331128 3324 331180 3330
rect 331128 3266 331180 3272
rect 330036 480 330064 3266
rect 331416 2530 331444 60030
rect 332704 4146 332732 60030
rect 333992 56658 334020 60030
rect 333900 56630 334020 56658
rect 332416 4140 332468 4146
rect 332416 4082 332468 4088
rect 332692 4140 332744 4146
rect 332692 4082 332744 4088
rect 331232 2502 331444 2530
rect 331232 480 331260 2502
rect 332428 480 332456 4082
rect 333900 2854 333928 56630
rect 334360 55622 334388 60166
rect 335372 60030 336214 60058
rect 334348 55616 334400 55622
rect 334348 55558 334400 55564
rect 334164 48340 334216 48346
rect 334164 48282 334216 48288
rect 334176 41426 334204 48282
rect 333992 41398 334204 41426
rect 333992 31822 334020 41398
rect 333980 31816 334032 31822
rect 333980 31758 334032 31764
rect 334072 31680 334124 31686
rect 334072 31622 334124 31628
rect 334084 18193 334112 31622
rect 334070 18184 334126 18193
rect 334070 18119 334126 18128
rect 333978 18048 334034 18057
rect 333978 17983 334034 17992
rect 333992 17950 334020 17983
rect 333980 17944 334032 17950
rect 333980 17886 334032 17892
rect 334072 8356 334124 8362
rect 334072 8298 334124 8304
rect 334084 3330 334112 8298
rect 335372 4146 335400 60030
rect 337212 56642 337240 60044
rect 338146 60030 338252 60058
rect 339158 60030 339448 60058
rect 338224 56642 338252 60030
rect 336740 56636 336792 56642
rect 336740 56578 336792 56584
rect 337200 56636 337252 56642
rect 337200 56578 337252 56584
rect 338120 56636 338172 56642
rect 338120 56578 338172 56584
rect 338212 56636 338264 56642
rect 338212 56578 338264 56584
rect 336752 56506 336780 56578
rect 336740 56500 336792 56506
rect 336740 56442 336792 56448
rect 336740 46980 336792 46986
rect 336740 46922 336792 46928
rect 336752 37262 336780 46922
rect 338132 46918 338160 56578
rect 338120 46912 338172 46918
rect 338120 46854 338172 46860
rect 338120 37324 338172 37330
rect 338120 37266 338172 37272
rect 336740 37256 336792 37262
rect 336740 37198 336792 37204
rect 336740 27668 336792 27674
rect 336740 27610 336792 27616
rect 336752 18170 336780 27610
rect 338132 27606 338160 37266
rect 338120 27600 338172 27606
rect 338120 27542 338172 27548
rect 336752 18142 336872 18170
rect 336844 18034 336872 18142
rect 336752 18006 336872 18034
rect 336752 17950 336780 18006
rect 336740 17944 336792 17950
rect 336740 17886 336792 17892
rect 338304 9716 338356 9722
rect 338304 9658 338356 9664
rect 337108 9580 337160 9586
rect 337108 9522 337160 9528
rect 335360 4140 335412 4146
rect 335360 4082 335412 4088
rect 335912 4140 335964 4146
rect 335912 4082 335964 4088
rect 334072 3324 334124 3330
rect 334072 3266 334124 3272
rect 334716 3324 334768 3330
rect 334716 3266 334768 3272
rect 333888 2848 333940 2854
rect 333888 2790 333940 2796
rect 333612 604 333664 610
rect 333612 546 333664 552
rect 333624 480 333652 546
rect 334728 480 334756 3266
rect 335924 480 335952 4082
rect 337120 480 337148 9522
rect 338316 480 338344 9658
rect 339420 4026 339448 60030
rect 339512 60030 340170 60058
rect 340892 60030 341090 60058
rect 342102 60030 342208 60058
rect 339512 4146 339540 60030
rect 339500 4140 339552 4146
rect 339500 4082 339552 4088
rect 340696 4140 340748 4146
rect 340696 4082 340748 4088
rect 339420 3998 339540 4026
rect 339512 480 339540 3998
rect 340708 480 340736 4082
rect 340892 3534 340920 60030
rect 342180 3534 342208 60030
rect 343008 56710 343036 60044
rect 344020 57662 344048 60044
rect 344008 57656 344060 57662
rect 344008 57598 344060 57604
rect 344928 57656 344980 57662
rect 344928 57598 344980 57604
rect 342996 56704 343048 56710
rect 342996 56646 343048 56652
rect 343732 56704 343784 56710
rect 343732 56646 343784 56652
rect 340880 3528 340932 3534
rect 340880 3470 340932 3476
rect 341892 3528 341944 3534
rect 341892 3470 341944 3476
rect 342168 3528 342220 3534
rect 342168 3470 342220 3476
rect 343088 3528 343140 3534
rect 343088 3470 343140 3476
rect 343744 3482 343772 56646
rect 344940 4146 344968 57598
rect 345032 56982 345060 60044
rect 345966 60030 346256 60058
rect 345020 56976 345072 56982
rect 345020 56918 345072 56924
rect 344928 4140 344980 4146
rect 344928 4082 344980 4088
rect 345480 4140 345532 4146
rect 345480 4082 345532 4088
rect 341904 480 341932 3470
rect 343100 480 343128 3470
rect 343744 3454 344324 3482
rect 344296 480 344324 3454
rect 345492 480 345520 4082
rect 346228 3466 346256 60030
rect 346964 57662 346992 60044
rect 347976 57798 348004 60044
rect 348910 60030 349016 60058
rect 347964 57792 348016 57798
rect 347964 57734 348016 57740
rect 346952 57656 347004 57662
rect 346952 57598 347004 57604
rect 347964 57656 348016 57662
rect 347964 57598 348016 57604
rect 346308 56976 346360 56982
rect 346308 56918 346360 56924
rect 346320 3482 346348 56918
rect 346216 3460 346268 3466
rect 346320 3454 346716 3482
rect 346216 3402 346268 3408
rect 346688 480 346716 3454
rect 347872 3460 347924 3466
rect 347872 3402 347924 3408
rect 347884 480 347912 3402
rect 347976 626 348004 57598
rect 348988 3602 349016 60030
rect 349068 57792 349120 57798
rect 349068 57734 349120 57740
rect 348976 3596 349028 3602
rect 348976 3538 349028 3544
rect 349080 3534 349108 57734
rect 349908 57594 349936 60044
rect 350920 57662 350948 60044
rect 351748 60030 351854 60058
rect 352866 60030 353248 60058
rect 350908 57656 350960 57662
rect 350908 57598 350960 57604
rect 349896 57588 349948 57594
rect 349896 57530 349948 57536
rect 351748 3602 351776 60030
rect 351828 57656 351880 57662
rect 351828 57598 351880 57604
rect 351368 3596 351420 3602
rect 351368 3538 351420 3544
rect 351736 3596 351788 3602
rect 351736 3538 351788 3544
rect 349068 3528 349120 3534
rect 349068 3470 349120 3476
rect 350264 3528 350316 3534
rect 350264 3470 350316 3476
rect 347976 598 349108 626
rect 349080 480 349108 598
rect 350276 480 350304 3470
rect 351380 480 351408 3538
rect 351840 3058 351868 57598
rect 352012 57588 352064 57594
rect 352012 57530 352064 57536
rect 352024 3482 352052 57530
rect 353220 4146 353248 60030
rect 353864 57118 353892 60044
rect 354784 57254 354812 60044
rect 355810 60030 356008 60058
rect 356822 60030 357388 60058
rect 354772 57248 354824 57254
rect 354772 57190 354824 57196
rect 355876 57248 355928 57254
rect 355876 57190 355928 57196
rect 353852 57112 353904 57118
rect 353852 57054 353904 57060
rect 353208 4140 353260 4146
rect 353208 4082 353260 4088
rect 354956 3596 355008 3602
rect 354956 3538 355008 3544
rect 352024 3454 352604 3482
rect 351828 3052 351880 3058
rect 351828 2994 351880 3000
rect 352576 480 352604 3454
rect 353760 3052 353812 3058
rect 353760 2994 353812 3000
rect 353772 480 353800 2994
rect 354968 480 354996 3538
rect 355888 3194 355916 57190
rect 355980 3466 356008 60030
rect 356152 57112 356204 57118
rect 356152 57054 356204 57060
rect 356164 4282 356192 57054
rect 357360 4434 357388 60030
rect 357728 57662 357756 60044
rect 357716 57656 357768 57662
rect 357716 57598 357768 57604
rect 358636 57656 358688 57662
rect 358636 57598 358688 57604
rect 357360 4406 357480 4434
rect 356152 4276 356204 4282
rect 356152 4218 356204 4224
rect 357348 4276 357400 4282
rect 357348 4218 357400 4224
rect 356152 4140 356204 4146
rect 356152 4082 356204 4088
rect 355968 3460 356020 3466
rect 355968 3402 356020 3408
rect 355876 3188 355928 3194
rect 355876 3130 355928 3136
rect 356164 480 356192 4082
rect 357360 480 357388 4218
rect 357452 4146 357480 4406
rect 357440 4140 357492 4146
rect 357440 4082 357492 4088
rect 358648 3330 358676 57598
rect 358740 3602 358768 60044
rect 359674 60030 360148 60058
rect 360120 3874 360148 60030
rect 360672 57662 360700 60044
rect 360660 57656 360712 57662
rect 360660 57598 360712 57604
rect 361684 57594 361712 60044
rect 362618 60030 362908 60058
rect 363630 60030 364288 60058
rect 362224 57656 362276 57662
rect 362224 57598 362276 57604
rect 361672 57588 361724 57594
rect 361672 57530 361724 57536
rect 362236 4146 362264 57598
rect 362776 57588 362828 57594
rect 362776 57530 362828 57536
rect 360936 4140 360988 4146
rect 360936 4082 360988 4088
rect 362224 4140 362276 4146
rect 362224 4082 362276 4088
rect 360108 3868 360160 3874
rect 360108 3810 360160 3816
rect 358728 3596 358780 3602
rect 358728 3538 358780 3544
rect 359740 3460 359792 3466
rect 359740 3402 359792 3408
rect 358636 3324 358688 3330
rect 358636 3266 358688 3272
rect 358544 3188 358596 3194
rect 358544 3130 358596 3136
rect 358556 480 358584 3130
rect 359752 480 359780 3402
rect 360948 480 360976 4082
rect 362788 4078 362816 57530
rect 362776 4072 362828 4078
rect 362776 4014 362828 4020
rect 362880 3670 362908 60030
rect 364260 3738 364288 60030
rect 364628 57594 364656 60044
rect 365562 60030 365668 60058
rect 366574 60030 367048 60058
rect 364616 57588 364668 57594
rect 364616 57530 364668 57536
rect 364524 3868 364576 3874
rect 364524 3810 364576 3816
rect 364248 3732 364300 3738
rect 364248 3674 364300 3680
rect 362868 3664 362920 3670
rect 362868 3606 362920 3612
rect 363328 3596 363380 3602
rect 363328 3538 363380 3544
rect 362132 3324 362184 3330
rect 362132 3266 362184 3272
rect 362144 480 362172 3266
rect 363340 480 363368 3538
rect 364536 480 364564 3810
rect 365640 3330 365668 60030
rect 365720 4140 365772 4146
rect 365720 4082 365772 4088
rect 365628 3324 365680 3330
rect 365628 3266 365680 3272
rect 365732 480 365760 4082
rect 366916 4072 366968 4078
rect 366916 4014 366968 4020
rect 366928 480 366956 4014
rect 367020 3534 367048 60030
rect 367572 57662 367600 60044
rect 368492 57662 368520 60044
rect 369518 60030 369808 60058
rect 370530 60030 371188 60058
rect 367560 57656 367612 57662
rect 367560 57598 367612 57604
rect 368388 57656 368440 57662
rect 368388 57598 368440 57604
rect 368480 57656 368532 57662
rect 368480 57598 368532 57604
rect 369676 57656 369728 57662
rect 369676 57598 369728 57604
rect 368020 3664 368072 3670
rect 368020 3606 368072 3612
rect 367008 3528 367060 3534
rect 367008 3470 367060 3476
rect 368032 480 368060 3606
rect 368400 3126 368428 57598
rect 369216 3732 369268 3738
rect 369216 3674 369268 3680
rect 368388 3120 368440 3126
rect 368388 3062 368440 3068
rect 369228 480 369256 3674
rect 369688 2922 369716 57598
rect 369780 3874 369808 60030
rect 369952 57588 370004 57594
rect 369952 57530 370004 57536
rect 369768 3868 369820 3874
rect 369768 3810 369820 3816
rect 369676 2916 369728 2922
rect 369676 2858 369728 2864
rect 369964 610 369992 57530
rect 371160 3806 371188 60030
rect 371436 57798 371464 60044
rect 372462 60030 372568 60058
rect 373474 60030 373948 60058
rect 371424 57792 371476 57798
rect 371424 57734 371476 57740
rect 371148 3800 371200 3806
rect 371148 3742 371200 3748
rect 372540 3466 372568 60030
rect 373920 3602 373948 60030
rect 374380 57662 374408 60044
rect 374644 57792 374696 57798
rect 374644 57734 374696 57740
rect 374368 57656 374420 57662
rect 374368 57598 374420 57604
rect 373908 3596 373960 3602
rect 373908 3538 373960 3544
rect 372804 3528 372856 3534
rect 372804 3470 372856 3476
rect 372528 3460 372580 3466
rect 372528 3402 372580 3408
rect 371608 3324 371660 3330
rect 371608 3266 371660 3272
rect 369952 604 370004 610
rect 369952 546 370004 552
rect 370412 604 370464 610
rect 370412 546 370464 552
rect 370424 480 370452 546
rect 371620 480 371648 3266
rect 372816 480 372844 3470
rect 374656 3330 374684 57734
rect 375392 57662 375420 60044
rect 376326 60030 376708 60058
rect 377338 60030 378088 60058
rect 375288 57656 375340 57662
rect 375288 57598 375340 57604
rect 375380 57656 375432 57662
rect 375380 57598 375432 57604
rect 376576 57656 376628 57662
rect 376576 57598 376628 57604
rect 375300 3398 375328 57598
rect 376392 3868 376444 3874
rect 376392 3810 376444 3816
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374644 3324 374696 3330
rect 374644 3266 374696 3272
rect 374000 3120 374052 3126
rect 374000 3062 374052 3068
rect 374012 480 374040 3062
rect 375196 2916 375248 2922
rect 375196 2858 375248 2864
rect 375208 480 375236 2858
rect 376404 480 376432 3810
rect 376588 3262 376616 57598
rect 376680 3534 376708 60030
rect 377588 3800 377640 3806
rect 377588 3742 377640 3748
rect 376668 3528 376720 3534
rect 376668 3470 376720 3476
rect 376576 3256 376628 3262
rect 376576 3198 376628 3204
rect 377600 480 377628 3742
rect 378060 3194 378088 60030
rect 378336 57594 378364 60044
rect 379256 57662 379284 60044
rect 380282 60030 380848 60058
rect 379244 57656 379296 57662
rect 379244 57598 379296 57604
rect 380164 57656 380216 57662
rect 380164 57598 380216 57604
rect 378324 57588 378376 57594
rect 378324 57530 378376 57536
rect 379428 57588 379480 57594
rect 379428 57530 379480 57536
rect 379440 4146 379468 57530
rect 379428 4140 379480 4146
rect 379428 4082 379480 4088
rect 380176 3466 380204 57598
rect 380820 3806 380848 60030
rect 381280 57662 381308 60044
rect 381268 57656 381320 57662
rect 381268 57598 381320 57604
rect 382096 57656 382148 57662
rect 382096 57598 382148 57604
rect 380808 3800 380860 3806
rect 380808 3742 380860 3748
rect 382108 3602 382136 57598
rect 382200 3942 382228 60044
rect 383226 60030 383608 60058
rect 382188 3936 382240 3942
rect 382188 3878 382240 3884
rect 383580 3874 383608 60030
rect 384224 57390 384252 60044
rect 384212 57384 384264 57390
rect 384212 57326 384264 57332
rect 384948 57384 385000 57390
rect 384948 57326 385000 57332
rect 384960 4078 384988 57326
rect 385144 57254 385172 60044
rect 386170 60030 386276 60058
rect 387182 60030 387748 60058
rect 385132 57248 385184 57254
rect 385132 57190 385184 57196
rect 384948 4072 385000 4078
rect 384948 4014 385000 4020
rect 383568 3868 383620 3874
rect 383568 3810 383620 3816
rect 381176 3596 381228 3602
rect 381176 3538 381228 3544
rect 382096 3596 382148 3602
rect 382096 3538 382148 3544
rect 379980 3460 380032 3466
rect 379980 3402 380032 3408
rect 380164 3460 380216 3466
rect 380164 3402 380216 3408
rect 378784 3324 378836 3330
rect 378784 3266 378836 3272
rect 378048 3188 378100 3194
rect 378048 3130 378100 3136
rect 378796 480 378824 3266
rect 379992 480 380020 3402
rect 381188 480 381216 3538
rect 386248 3534 386276 60030
rect 386328 57248 386380 57254
rect 386328 57190 386380 57196
rect 386340 4010 386368 57190
rect 387064 4140 387116 4146
rect 387064 4082 387116 4088
rect 386328 4004 386380 4010
rect 386328 3946 386380 3952
rect 384672 3528 384724 3534
rect 384672 3470 384724 3476
rect 386236 3528 386288 3534
rect 386236 3470 386288 3476
rect 382372 3392 382424 3398
rect 382372 3334 382424 3340
rect 382384 480 382412 3334
rect 383568 3256 383620 3262
rect 383568 3198 383620 3204
rect 383580 480 383608 3198
rect 384684 480 384712 3470
rect 385868 3188 385920 3194
rect 385868 3130 385920 3136
rect 385880 480 385908 3130
rect 387076 480 387104 4082
rect 387720 3670 387748 60030
rect 388088 57662 388116 60044
rect 389008 60030 389114 60058
rect 390126 60030 390508 60058
rect 388076 57656 388128 57662
rect 388076 57598 388128 57604
rect 387708 3664 387760 3670
rect 387708 3606 387760 3612
rect 389008 3466 389036 60030
rect 389088 57656 389140 57662
rect 389088 57598 389140 57604
rect 389100 3738 389128 57598
rect 390480 3806 390508 60030
rect 391032 57662 391060 60044
rect 392044 57662 392072 60044
rect 392978 60030 393176 60058
rect 393990 60030 394648 60058
rect 391020 57656 391072 57662
rect 391020 57598 391072 57604
rect 391848 57656 391900 57662
rect 391848 57598 391900 57604
rect 392032 57656 392084 57662
rect 392032 57598 392084 57604
rect 391756 3936 391808 3942
rect 391756 3878 391808 3884
rect 389456 3800 389508 3806
rect 389456 3742 389508 3748
rect 390468 3800 390520 3806
rect 390468 3742 390520 3748
rect 389088 3732 389140 3738
rect 389088 3674 389140 3680
rect 388260 3460 388312 3466
rect 388260 3402 388312 3408
rect 388996 3460 389048 3466
rect 388996 3402 389048 3408
rect 388272 480 388300 3402
rect 389468 480 389496 3742
rect 390652 3596 390704 3602
rect 390652 3538 390704 3544
rect 390664 480 390692 3538
rect 391768 3210 391796 3878
rect 391860 3398 391888 57598
rect 393148 3942 393176 60030
rect 393228 57656 393280 57662
rect 393228 57598 393280 57604
rect 393136 3936 393188 3942
rect 393136 3878 393188 3884
rect 393240 3874 393268 57598
rect 394240 4072 394292 4078
rect 394240 4014 394292 4020
rect 393044 3868 393096 3874
rect 393044 3810 393096 3816
rect 393228 3868 393280 3874
rect 393228 3810 393280 3816
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391768 3182 391888 3210
rect 391860 480 391888 3182
rect 393056 480 393084 3810
rect 394252 480 394280 4014
rect 394620 3262 394648 60030
rect 394988 57662 395016 60044
rect 395922 60030 396028 60058
rect 396934 60030 397408 60058
rect 394976 57656 395028 57662
rect 394976 57598 395028 57604
rect 395896 57656 395948 57662
rect 395896 57598 395948 57604
rect 395908 4078 395936 57598
rect 395896 4072 395948 4078
rect 395896 4014 395948 4020
rect 395436 4004 395488 4010
rect 395436 3946 395488 3952
rect 394608 3256 394660 3262
rect 394608 3198 394660 3204
rect 395448 480 395476 3946
rect 396000 3602 396028 60030
rect 397380 4146 397408 60030
rect 397932 57662 397960 60044
rect 398852 57662 398880 60044
rect 399878 60030 400168 60058
rect 400890 60030 401548 60058
rect 397920 57656 397972 57662
rect 397920 57598 397972 57604
rect 398748 57656 398800 57662
rect 398748 57598 398800 57604
rect 398840 57656 398892 57662
rect 398840 57598 398892 57604
rect 400036 57656 400088 57662
rect 400036 57598 400088 57604
rect 397368 4140 397420 4146
rect 397368 4082 397420 4088
rect 397828 3664 397880 3670
rect 397828 3606 397880 3612
rect 395988 3596 396040 3602
rect 395988 3538 396040 3544
rect 396632 3528 396684 3534
rect 396632 3470 396684 3476
rect 396644 480 396672 3470
rect 397840 480 397868 3606
rect 398760 3330 398788 57598
rect 400048 4010 400076 57598
rect 400036 4004 400088 4010
rect 400036 3946 400088 3952
rect 400140 3738 400168 60030
rect 401520 3806 401548 60030
rect 401796 57662 401824 60044
rect 402822 60030 402928 60058
rect 403834 60030 404308 60058
rect 401784 57656 401836 57662
rect 401784 57598 401836 57604
rect 402796 57656 402848 57662
rect 402796 57598 402848 57604
rect 401324 3800 401376 3806
rect 401324 3742 401376 3748
rect 401508 3800 401560 3806
rect 401508 3742 401560 3748
rect 399024 3732 399076 3738
rect 399024 3674 399076 3680
rect 400128 3732 400180 3738
rect 400128 3674 400180 3680
rect 398748 3324 398800 3330
rect 398748 3266 398800 3272
rect 399036 480 399064 3674
rect 400220 3460 400272 3466
rect 400220 3402 400272 3408
rect 400232 480 400260 3402
rect 401336 480 401364 3742
rect 402808 3670 402836 57598
rect 402796 3664 402848 3670
rect 402796 3606 402848 3612
rect 402900 3534 402928 60030
rect 404280 3874 404308 60030
rect 404740 57662 404768 60044
rect 404728 57656 404780 57662
rect 404728 57598 404780 57604
rect 405648 57656 405700 57662
rect 405648 57598 405700 57604
rect 404912 3936 404964 3942
rect 404912 3878 404964 3884
rect 403716 3868 403768 3874
rect 403716 3810 403768 3816
rect 404268 3868 404320 3874
rect 404268 3810 404320 3816
rect 402888 3528 402940 3534
rect 402888 3470 402940 3476
rect 402520 3392 402572 3398
rect 402520 3334 402572 3340
rect 402532 480 402560 3334
rect 403728 480 403756 3810
rect 404924 480 404952 3878
rect 405660 3398 405688 57598
rect 405752 57118 405780 60044
rect 406778 60030 407068 60058
rect 407698 60030 408448 60058
rect 405740 57112 405792 57118
rect 405740 57054 405792 57060
rect 406936 57112 406988 57118
rect 406936 57054 406988 57060
rect 405648 3392 405700 3398
rect 405648 3334 405700 3340
rect 406948 3262 406976 57054
rect 407040 3942 407068 60030
rect 407304 4072 407356 4078
rect 407304 4014 407356 4020
rect 407028 3936 407080 3942
rect 407028 3878 407080 3884
rect 406108 3256 406160 3262
rect 406108 3198 406160 3204
rect 406936 3256 406988 3262
rect 406936 3198 406988 3204
rect 406120 480 406148 3198
rect 407316 480 407344 4014
rect 408420 3466 408448 60030
rect 408696 57662 408724 60044
rect 409630 60030 409828 60058
rect 410642 60030 411208 60058
rect 408684 57656 408736 57662
rect 408684 57598 408736 57604
rect 409696 57656 409748 57662
rect 409696 57598 409748 57604
rect 409708 4146 409736 57598
rect 409604 4140 409656 4146
rect 409604 4082 409656 4088
rect 409696 4140 409748 4146
rect 409696 4082 409748 4088
rect 409616 4026 409644 4082
rect 409616 3998 409736 4026
rect 408500 3596 408552 3602
rect 408500 3538 408552 3544
rect 408408 3460 408460 3466
rect 408408 3402 408460 3408
rect 408512 480 408540 3538
rect 409708 480 409736 3998
rect 409800 3602 409828 60030
rect 409788 3596 409840 3602
rect 409788 3538 409840 3544
rect 410892 3324 410944 3330
rect 410892 3266 410944 3272
rect 410904 480 410932 3266
rect 411180 3194 411208 60030
rect 411640 57662 411668 60044
rect 411628 57656 411680 57662
rect 411628 57598 411680 57604
rect 412456 57656 412508 57662
rect 412456 57598 412508 57604
rect 412468 4078 412496 57598
rect 412456 4072 412508 4078
rect 412456 4014 412508 4020
rect 412560 4010 412588 60044
rect 413586 60030 413968 60058
rect 412088 4004 412140 4010
rect 412088 3946 412140 3952
rect 412548 4004 412600 4010
rect 412548 3946 412600 3952
rect 411168 3188 411220 3194
rect 411168 3130 411220 3136
rect 412100 480 412128 3946
rect 413940 3738 413968 60030
rect 414584 57390 414612 60044
rect 414572 57384 414624 57390
rect 414572 57326 414624 57332
rect 415308 57384 415360 57390
rect 415308 57326 415360 57332
rect 415320 3806 415348 57326
rect 415504 57254 415532 60044
rect 416530 60030 416636 60058
rect 417542 60030 418108 60058
rect 415492 57248 415544 57254
rect 415492 57190 415544 57196
rect 414480 3800 414532 3806
rect 414480 3742 414532 3748
rect 415308 3800 415360 3806
rect 415308 3742 415360 3748
rect 413284 3732 413336 3738
rect 413284 3674 413336 3680
rect 413928 3732 413980 3738
rect 413928 3674 413980 3680
rect 413296 480 413324 3674
rect 414492 480 414520 3742
rect 416608 3670 416636 60030
rect 416688 57248 416740 57254
rect 416688 57190 416740 57196
rect 415676 3664 415728 3670
rect 415676 3606 415728 3612
rect 416596 3664 416648 3670
rect 416596 3606 416648 3612
rect 415688 480 415716 3606
rect 416700 3330 416728 57190
rect 418080 3874 418108 60030
rect 418448 57662 418476 60044
rect 419368 60030 419474 60058
rect 420486 60030 420868 60058
rect 418436 57656 418488 57662
rect 418436 57598 418488 57604
rect 417976 3868 418028 3874
rect 417976 3810 418028 3816
rect 418068 3868 418120 3874
rect 418068 3810 418120 3816
rect 416872 3528 416924 3534
rect 416872 3470 416924 3476
rect 416688 3324 416740 3330
rect 416688 3266 416740 3272
rect 416884 480 416912 3470
rect 417988 480 418016 3810
rect 419368 3534 419396 60030
rect 419448 57656 419500 57662
rect 419448 57598 419500 57604
rect 419356 3528 419408 3534
rect 419356 3470 419408 3476
rect 419460 3398 419488 57598
rect 419172 3392 419224 3398
rect 419172 3334 419224 3340
rect 419448 3392 419500 3398
rect 419448 3334 419500 3340
rect 419184 480 419212 3334
rect 420368 3256 420420 3262
rect 420368 3198 420420 3204
rect 420380 480 420408 3198
rect 420840 2990 420868 60030
rect 421392 57662 421420 60044
rect 422404 57662 422432 60044
rect 423430 60030 423628 60058
rect 424350 60030 425008 60058
rect 421380 57656 421432 57662
rect 421380 57598 421432 57604
rect 422208 57656 422260 57662
rect 422208 57598 422260 57604
rect 422392 57656 422444 57662
rect 422392 57598 422444 57604
rect 423496 57656 423548 57662
rect 423496 57598 423548 57604
rect 421564 3936 421616 3942
rect 421564 3878 421616 3884
rect 420828 2984 420880 2990
rect 420828 2926 420880 2932
rect 421576 480 421604 3878
rect 422220 3058 422248 57598
rect 423508 3942 423536 57598
rect 423496 3936 423548 3942
rect 423496 3878 423548 3884
rect 423600 3466 423628 60030
rect 423956 4140 424008 4146
rect 423956 4082 424008 4088
rect 422760 3460 422812 3466
rect 422760 3402 422812 3408
rect 423588 3460 423640 3466
rect 423588 3402 423640 3408
rect 422208 3052 422260 3058
rect 422208 2994 422260 3000
rect 422772 480 422800 3402
rect 423968 480 423996 4082
rect 424980 3262 425008 60030
rect 425348 57662 425376 60044
rect 426282 60030 426388 60058
rect 427294 60030 427768 60058
rect 425336 57656 425388 57662
rect 425336 57598 425388 57604
rect 426256 57656 426308 57662
rect 426256 57598 426308 57604
rect 425152 3596 425204 3602
rect 425152 3538 425204 3544
rect 424968 3256 425020 3262
rect 424968 3198 425020 3204
rect 425164 480 425192 3538
rect 426268 3126 426296 57598
rect 426360 3602 426388 60030
rect 427544 4072 427596 4078
rect 427544 4014 427596 4020
rect 426348 3596 426400 3602
rect 426348 3538 426400 3544
rect 426348 3188 426400 3194
rect 426348 3130 426400 3136
rect 426256 3120 426308 3126
rect 426256 3062 426308 3068
rect 426360 480 426388 3130
rect 427556 480 427584 4014
rect 427740 3194 427768 60030
rect 428292 57662 428320 60044
rect 428280 57656 428332 57662
rect 428280 57598 428332 57604
rect 429108 57656 429160 57662
rect 429108 57598 429160 57604
rect 429120 4010 429148 57598
rect 429212 57594 429240 60044
rect 430238 60030 430436 60058
rect 431250 60030 431908 60058
rect 429200 57588 429252 57594
rect 429200 57530 429252 57536
rect 430408 4146 430436 60030
rect 430488 57588 430540 57594
rect 430488 57530 430540 57536
rect 430396 4140 430448 4146
rect 430396 4082 430448 4088
rect 430500 4078 430528 57530
rect 431880 4146 431908 60030
rect 432156 57662 432184 60044
rect 433182 60030 433288 60058
rect 434194 60030 434668 60058
rect 432144 57656 432196 57662
rect 432144 57598 432196 57604
rect 433156 57656 433208 57662
rect 433156 57598 433208 57604
rect 431868 4140 431920 4146
rect 431868 4082 431920 4088
rect 430488 4072 430540 4078
rect 430488 4014 430540 4020
rect 428740 4004 428792 4010
rect 428740 3946 428792 3952
rect 429108 4004 429160 4010
rect 429108 3946 429160 3952
rect 427728 3188 427780 3194
rect 427728 3130 427780 3136
rect 428752 480 428780 3946
rect 431132 3800 431184 3806
rect 431132 3742 431184 3748
rect 429936 3732 429988 3738
rect 429936 3674 429988 3680
rect 429948 480 429976 3674
rect 431144 480 431172 3742
rect 433168 3330 433196 57598
rect 433260 3806 433288 60030
rect 434640 3874 434668 60030
rect 435100 57662 435128 60044
rect 435088 57656 435140 57662
rect 435088 57598 435140 57604
rect 436008 57656 436060 57662
rect 436008 57598 436060 57604
rect 434536 3868 434588 3874
rect 434536 3810 434588 3816
rect 434628 3868 434680 3874
rect 434628 3810 434680 3816
rect 433248 3800 433300 3806
rect 433248 3742 433300 3748
rect 434548 3754 434576 3810
rect 434548 3726 434668 3754
rect 433524 3664 433576 3670
rect 433524 3606 433576 3612
rect 432328 3324 432380 3330
rect 432328 3266 432380 3272
rect 433156 3324 433208 3330
rect 433156 3266 433208 3272
rect 432340 480 432368 3266
rect 433536 480 433564 3606
rect 434640 480 434668 3726
rect 435824 3392 435876 3398
rect 435824 3334 435876 3340
rect 435836 480 435864 3334
rect 436020 2922 436048 57598
rect 436112 57118 436140 60044
rect 437124 57254 437152 60044
rect 438058 60030 438808 60058
rect 437112 57248 437164 57254
rect 437112 57190 437164 57196
rect 436100 57112 436152 57118
rect 436100 57054 436152 57060
rect 437388 57112 437440 57118
rect 437388 57054 437440 57060
rect 437020 3528 437072 3534
rect 437020 3470 437072 3476
rect 436008 2916 436060 2922
rect 436008 2858 436060 2864
rect 437032 480 437060 3470
rect 437400 3398 437428 57054
rect 438780 3670 438808 60030
rect 439056 57662 439084 60044
rect 439044 57656 439096 57662
rect 439044 57598 439096 57604
rect 438768 3664 438820 3670
rect 438768 3606 438820 3612
rect 440068 3534 440096 60044
rect 441002 60030 441568 60058
rect 440148 57656 440200 57662
rect 440148 57598 440200 57604
rect 440056 3528 440108 3534
rect 440056 3470 440108 3476
rect 437388 3392 437440 3398
rect 437388 3334 437440 3340
rect 440160 3058 440188 57598
rect 441540 3942 441568 60030
rect 442000 57662 442028 60044
rect 442828 60030 442934 60058
rect 443946 60030 444328 60058
rect 441988 57656 442040 57662
rect 441988 57598 442040 57604
rect 440608 3936 440660 3942
rect 440608 3878 440660 3884
rect 441528 3936 441580 3942
rect 441528 3878 441580 3884
rect 439412 3052 439464 3058
rect 439412 2994 439464 3000
rect 440148 3052 440200 3058
rect 440148 2994 440200 3000
rect 438216 2984 438268 2990
rect 438216 2926 438268 2932
rect 438228 480 438256 2926
rect 439424 480 439452 2994
rect 440620 480 440648 3878
rect 442828 3466 442856 60030
rect 442908 57656 442960 57662
rect 442908 57598 442960 57604
rect 441804 3460 441856 3466
rect 441804 3402 441856 3408
rect 442816 3460 442868 3466
rect 442816 3402 442868 3408
rect 441816 480 441844 3402
rect 442920 2990 442948 57598
rect 444300 3262 444328 60030
rect 444944 57390 444972 60044
rect 444932 57384 444984 57390
rect 444932 57326 444984 57332
rect 445668 57384 445720 57390
rect 445668 57326 445720 57332
rect 445680 3806 445708 57326
rect 445864 57118 445892 60044
rect 446890 60030 447088 60058
rect 447902 60030 448468 60058
rect 445852 57112 445904 57118
rect 445852 57054 445904 57060
rect 446956 57112 447008 57118
rect 446956 57054 447008 57060
rect 445668 3800 445720 3806
rect 445668 3742 445720 3748
rect 445392 3596 445444 3602
rect 445392 3538 445444 3544
rect 443000 3256 443052 3262
rect 443000 3198 443052 3204
rect 444288 3256 444340 3262
rect 444288 3198 444340 3204
rect 442908 2984 442960 2990
rect 442908 2926 442960 2932
rect 443012 480 443040 3198
rect 444196 3120 444248 3126
rect 444196 3062 444248 3068
rect 444208 480 444236 3062
rect 445404 480 445432 3538
rect 446588 3188 446640 3194
rect 446588 3130 446640 3136
rect 446600 480 446628 3130
rect 446968 3126 446996 57054
rect 447060 3738 447088 60030
rect 447784 4004 447836 4010
rect 447784 3946 447836 3952
rect 447048 3732 447100 3738
rect 447048 3674 447100 3680
rect 446956 3120 447008 3126
rect 446956 3062 447008 3068
rect 447796 480 447824 3946
rect 448440 3126 448468 60030
rect 448808 57662 448836 60044
rect 448796 57656 448848 57662
rect 448796 57598 448848 57604
rect 449716 57656 449768 57662
rect 449716 57598 449768 57604
rect 449728 4078 449756 57598
rect 448980 4072 449032 4078
rect 448980 4014 449032 4020
rect 449716 4072 449768 4078
rect 449716 4014 449768 4020
rect 448336 3120 448388 3126
rect 448334 3088 448336 3097
rect 448428 3120 448480 3126
rect 448388 3088 448390 3097
rect 448428 3062 448480 3068
rect 448334 3023 448390 3032
rect 448992 480 449020 4014
rect 449820 4010 449848 60044
rect 450846 60030 451228 60058
rect 449808 4004 449860 4010
rect 449808 3946 449860 3952
rect 451200 3602 451228 60030
rect 451752 57662 451780 60044
rect 452764 57662 452792 60044
rect 453790 60030 453896 60058
rect 454710 60030 455368 60058
rect 451740 57656 451792 57662
rect 451740 57598 451792 57604
rect 452568 57656 452620 57662
rect 452568 57598 452620 57604
rect 452752 57656 452804 57662
rect 452752 57598 452804 57604
rect 452580 4146 452608 57598
rect 451280 4140 451332 4146
rect 451280 4082 451332 4088
rect 452568 4140 452620 4146
rect 452568 4082 452620 4088
rect 450176 3596 450228 3602
rect 450176 3538 450228 3544
rect 451188 3596 451240 3602
rect 451188 3538 451240 3544
rect 450188 480 450216 3538
rect 451186 3088 451242 3097
rect 451186 3023 451188 3032
rect 451240 3023 451242 3032
rect 451188 2994 451240 3000
rect 451292 480 451320 4082
rect 453868 3806 453896 60030
rect 453948 57656 454000 57662
rect 453948 57598 454000 57604
rect 453960 4214 453988 57598
rect 453948 4208 454000 4214
rect 453948 4150 454000 4156
rect 454868 3868 454920 3874
rect 454868 3810 454920 3816
rect 453856 3800 453908 3806
rect 453856 3742 453908 3748
rect 452476 3324 452528 3330
rect 452476 3266 452528 3272
rect 452488 480 452516 3266
rect 452580 3194 452700 3210
rect 452568 3188 452700 3194
rect 452620 3182 452700 3188
rect 452568 3130 452620 3136
rect 452672 2854 452700 3182
rect 452660 2848 452712 2854
rect 452660 2790 452712 2796
rect 453672 2848 453724 2854
rect 453672 2790 453724 2796
rect 453684 480 453712 2790
rect 454880 480 454908 3810
rect 455340 3330 455368 60030
rect 455708 57662 455736 60044
rect 456628 60030 456734 60058
rect 455696 57656 455748 57662
rect 455696 57598 455748 57604
rect 456064 3664 456116 3670
rect 456340 3664 456392 3670
rect 456116 3612 456340 3618
rect 456064 3606 456392 3612
rect 456076 3590 456380 3606
rect 456628 3369 456656 60030
rect 456708 57656 456760 57662
rect 456708 57598 456760 57604
rect 456720 3874 456748 57598
rect 457640 57390 457668 60044
rect 458652 57662 458680 60044
rect 459572 57662 459600 60044
rect 460584 57934 460612 60044
rect 461610 60030 462268 60058
rect 460572 57928 460624 57934
rect 460572 57870 460624 57876
rect 458640 57656 458692 57662
rect 458640 57598 458692 57604
rect 459468 57656 459520 57662
rect 459468 57598 459520 57604
rect 459560 57656 459612 57662
rect 459560 57598 459612 57604
rect 460848 57656 460900 57662
rect 460848 57598 460900 57604
rect 457628 57384 457680 57390
rect 457628 57326 457680 57332
rect 458272 57248 458324 57254
rect 458272 57190 458324 57196
rect 456708 3868 456760 3874
rect 456708 3810 456760 3816
rect 457260 3392 457312 3398
rect 456614 3360 456670 3369
rect 455328 3324 455380 3330
rect 457260 3334 457312 3340
rect 456614 3295 456670 3304
rect 455328 3266 455380 3272
rect 456064 2916 456116 2922
rect 456064 2858 456116 2864
rect 456076 480 456104 2858
rect 457272 480 457300 3334
rect 458284 626 458312 57190
rect 459480 3738 459508 57598
rect 459468 3732 459520 3738
rect 459468 3674 459520 3680
rect 460860 3670 460888 57598
rect 462044 3936 462096 3942
rect 462044 3878 462096 3884
rect 459652 3664 459704 3670
rect 459652 3606 459704 3612
rect 460848 3664 460900 3670
rect 460848 3606 460900 3612
rect 458284 598 458496 626
rect 458468 480 458496 598
rect 459664 480 459692 3606
rect 460756 2848 460808 2854
rect 460808 2796 460888 2802
rect 460756 2790 460888 2796
rect 460768 2774 460888 2790
rect 460860 480 460888 2774
rect 462056 480 462084 3878
rect 462240 3874 462268 60030
rect 462516 57662 462544 60044
rect 462504 57656 462556 57662
rect 462504 57598 462556 57604
rect 463528 57322 463556 60044
rect 464554 60030 465028 60058
rect 463608 57656 463660 57662
rect 463608 57598 463660 57604
rect 463516 57316 463568 57322
rect 463516 57258 463568 57264
rect 462228 3868 462280 3874
rect 462228 3810 462280 3816
rect 463620 3534 463648 57598
rect 465000 3942 465028 60030
rect 465460 57662 465488 60044
rect 466472 57730 466500 60044
rect 467498 60030 467788 60058
rect 468418 60030 469168 60058
rect 466460 57724 466512 57730
rect 466460 57666 466512 57672
rect 465448 57656 465500 57662
rect 465448 57598 465500 57604
rect 466368 57656 466420 57662
rect 466368 57598 466420 57604
rect 464988 3936 465040 3942
rect 464988 3878 465040 3884
rect 463240 3528 463292 3534
rect 463240 3470 463292 3476
rect 463608 3528 463660 3534
rect 463608 3470 463660 3476
rect 463252 480 463280 3470
rect 466380 3466 466408 57598
rect 465632 3460 465684 3466
rect 465632 3402 465684 3408
rect 466368 3460 466420 3466
rect 466368 3402 466420 3408
rect 464436 2984 464488 2990
rect 464436 2926 464488 2932
rect 464448 480 464476 2926
rect 465644 480 465672 3402
rect 466828 3256 466880 3262
rect 466828 3198 466880 3204
rect 466840 480 466868 3198
rect 467760 2990 467788 60030
rect 469140 3194 469168 60030
rect 469416 57662 469444 60044
rect 470442 60030 470548 60058
rect 471362 60030 471928 60058
rect 469404 57656 469456 57662
rect 469404 57598 469456 57604
rect 470520 3602 470548 60030
rect 471900 3806 471928 60030
rect 472360 57458 472388 60044
rect 473372 57594 473400 60044
rect 474306 60030 474688 60058
rect 473360 57588 473412 57594
rect 473360 57530 473412 57536
rect 474556 57588 474608 57594
rect 474556 57530 474608 57536
rect 472348 57452 472400 57458
rect 472348 57394 472400 57400
rect 474568 4078 474596 57530
rect 472716 4072 472768 4078
rect 472716 4014 472768 4020
rect 474556 4072 474608 4078
rect 474556 4014 474608 4020
rect 471888 3800 471940 3806
rect 471888 3742 471940 3748
rect 470324 3596 470376 3602
rect 470324 3538 470376 3544
rect 470508 3596 470560 3602
rect 470508 3538 470560 3544
rect 469128 3188 469180 3194
rect 469128 3130 469180 3136
rect 467932 3120 467984 3126
rect 467932 3062 467984 3068
rect 467748 2984 467800 2990
rect 467748 2926 467800 2932
rect 467944 480 467972 3062
rect 469128 3052 469180 3058
rect 469128 2994 469180 3000
rect 469140 480 469168 2994
rect 470336 480 470364 3538
rect 471520 3528 471572 3534
rect 471520 3470 471572 3476
rect 471532 480 471560 3470
rect 472728 480 472756 4014
rect 473912 4004 473964 4010
rect 473912 3946 473964 3952
rect 473924 480 473952 3946
rect 474660 3194 474688 60030
rect 475304 57594 475332 60044
rect 475292 57588 475344 57594
rect 475292 57530 475344 57536
rect 476224 56982 476252 60044
rect 477250 60030 477356 60058
rect 476212 56976 476264 56982
rect 476212 56918 476264 56924
rect 476304 4140 476356 4146
rect 476304 4082 476356 4088
rect 475108 3324 475160 3330
rect 475108 3266 475160 3272
rect 474648 3188 474700 3194
rect 474648 3130 474700 3136
rect 475120 480 475148 3266
rect 476316 480 476344 4082
rect 477328 4010 477356 60030
rect 478248 57526 478276 60044
rect 478236 57520 478288 57526
rect 478236 57462 478288 57468
rect 479168 57254 479196 60044
rect 480180 57866 480208 60044
rect 480168 57860 480220 57866
rect 480168 57802 480220 57808
rect 481192 57254 481220 60044
rect 482112 57798 482140 60044
rect 483124 57798 483152 60044
rect 482100 57792 482152 57798
rect 482100 57734 482152 57740
rect 482928 57792 482980 57798
rect 482928 57734 482980 57740
rect 483112 57792 483164 57798
rect 483112 57734 483164 57740
rect 479156 57248 479208 57254
rect 479156 57190 479208 57196
rect 480168 57248 480220 57254
rect 480168 57190 480220 57196
rect 481180 57248 481232 57254
rect 481180 57190 481232 57196
rect 477408 56976 477460 56982
rect 477408 56918 477460 56924
rect 477316 4004 477368 4010
rect 477316 3946 477368 3952
rect 477420 3262 477448 56918
rect 480180 3330 480208 57190
rect 482940 3398 482968 57734
rect 484136 57390 484164 60044
rect 485070 60030 485728 60058
rect 484308 57792 484360 57798
rect 484308 57734 484360 57740
rect 483112 57384 483164 57390
rect 483112 57326 483164 57332
rect 484124 57384 484176 57390
rect 484124 57326 484176 57332
rect 481088 3392 481140 3398
rect 482928 3392 482980 3398
rect 481088 3334 481140 3340
rect 482282 3360 482338 3369
rect 478696 3324 478748 3330
rect 478696 3266 478748 3272
rect 480168 3324 480220 3330
rect 480168 3266 480220 3272
rect 477408 3256 477460 3262
rect 477408 3198 477460 3204
rect 477500 2848 477552 2854
rect 477500 2790 477552 2796
rect 477512 480 477540 2790
rect 478708 480 478736 3266
rect 479892 2916 479944 2922
rect 479892 2858 479944 2864
rect 479904 480 479932 2858
rect 481100 480 481128 3334
rect 482928 3334 482980 3340
rect 482282 3295 482338 3304
rect 482296 480 482324 3295
rect 483124 626 483152 57326
rect 484320 4146 484348 57734
rect 484308 4140 484360 4146
rect 484308 4082 484360 4088
rect 485700 3806 485728 60030
rect 485964 57928 486016 57934
rect 485964 57870 486016 57876
rect 485688 3800 485740 3806
rect 485688 3742 485740 3748
rect 484584 3732 484636 3738
rect 484584 3674 484636 3680
rect 483124 598 483520 626
rect 483492 480 483520 598
rect 484596 480 484624 3674
rect 485780 3664 485832 3670
rect 485780 3606 485832 3612
rect 485792 480 485820 3606
rect 485976 610 486004 57870
rect 486068 56982 486096 60044
rect 486056 56976 486108 56982
rect 486056 56918 486108 56924
rect 487080 4826 487108 60044
rect 488014 60030 488488 60058
rect 487068 4820 487120 4826
rect 487068 4762 487120 4768
rect 488172 3868 488224 3874
rect 488172 3810 488224 3816
rect 485964 604 486016 610
rect 485964 546 486016 552
rect 486976 604 487028 610
rect 486976 546 487028 552
rect 486988 480 487016 546
rect 488184 480 488212 3810
rect 488460 3738 488488 60030
rect 489012 57798 489040 60044
rect 489184 57860 489236 57866
rect 489184 57802 489236 57808
rect 489000 57792 489052 57798
rect 489000 57734 489052 57740
rect 488448 3732 488500 3738
rect 488448 3674 488500 3680
rect 489196 2854 489224 57802
rect 489828 57792 489880 57798
rect 489828 57734 489880 57740
rect 489840 3874 489868 57734
rect 490024 57118 490052 60044
rect 490958 60030 491248 60058
rect 491970 60030 492628 60058
rect 490104 57316 490156 57322
rect 490104 57258 490156 57264
rect 490012 57112 490064 57118
rect 490012 57054 490064 57060
rect 489828 3868 489880 3874
rect 489828 3810 489880 3816
rect 490116 3346 490144 57258
rect 491220 3670 491248 60030
rect 491944 56976 491996 56982
rect 491944 56918 491996 56924
rect 491760 3936 491812 3942
rect 491760 3878 491812 3884
rect 491208 3664 491260 3670
rect 491208 3606 491260 3612
rect 490116 3318 490604 3346
rect 489368 2984 489420 2990
rect 489368 2926 489420 2932
rect 489184 2848 489236 2854
rect 489184 2790 489236 2796
rect 489380 480 489408 2926
rect 490576 480 490604 3318
rect 491772 480 491800 3878
rect 491956 2922 491984 56918
rect 492600 3942 492628 60030
rect 492876 57322 492904 60044
rect 493902 60030 494008 60058
rect 492864 57316 492916 57322
rect 492864 57258 492916 57264
rect 492588 3936 492640 3942
rect 492588 3878 492640 3884
rect 493980 3534 494008 60030
rect 494244 57724 494296 57730
rect 494244 57666 494296 57672
rect 492956 3528 493008 3534
rect 492956 3470 493008 3476
rect 493968 3528 494020 3534
rect 494256 3482 494284 57666
rect 494900 57186 494928 60044
rect 494888 57180 494940 57186
rect 494888 57122 494940 57128
rect 495820 57050 495848 60044
rect 496832 57662 496860 60044
rect 497844 57934 497872 60044
rect 497832 57928 497884 57934
rect 497832 57870 497884 57876
rect 498764 57798 498792 60044
rect 498752 57792 498804 57798
rect 498752 57734 498804 57740
rect 496912 57724 496964 57730
rect 496912 57666 496964 57672
rect 496820 57656 496872 57662
rect 496820 57598 496872 57604
rect 495808 57044 495860 57050
rect 495808 56986 495860 56992
rect 493968 3470 494020 3476
rect 491944 2916 491996 2922
rect 491944 2858 491996 2864
rect 492968 480 492996 3470
rect 494164 3454 494284 3482
rect 494164 480 494192 3454
rect 496924 3346 496952 57666
rect 499776 57662 499804 60044
rect 498108 57656 498160 57662
rect 498108 57598 498160 57604
rect 499764 57656 499816 57662
rect 499764 57598 499816 57604
rect 496924 3318 497780 3346
rect 496544 3120 496596 3126
rect 496544 3062 496596 3068
rect 495348 3052 495400 3058
rect 495348 2994 495400 3000
rect 495360 480 495388 2994
rect 496556 480 496584 3062
rect 497752 480 497780 3318
rect 498120 2990 498148 57598
rect 498936 3596 498988 3602
rect 498936 3538 498988 3544
rect 498108 2984 498160 2990
rect 498108 2926 498160 2932
rect 498948 480 498976 3538
rect 500788 3466 500816 60044
rect 501722 60030 502288 60058
rect 500868 57656 500920 57662
rect 500868 57598 500920 57604
rect 500880 3602 500908 57598
rect 501052 57452 501104 57458
rect 501052 57394 501104 57400
rect 500868 3596 500920 3602
rect 500868 3538 500920 3544
rect 500132 3460 500184 3466
rect 500132 3402 500184 3408
rect 500776 3460 500828 3466
rect 500776 3402 500828 3408
rect 500144 480 500172 3402
rect 501064 610 501092 57394
rect 502260 5234 502288 60030
rect 502720 57662 502748 60044
rect 503746 60030 504128 60058
rect 504666 60030 505048 60058
rect 502708 57656 502760 57662
rect 502708 57598 502760 57604
rect 503628 57656 503680 57662
rect 503628 57598 503680 57604
rect 502248 5228 502300 5234
rect 502248 5170 502300 5176
rect 503640 4078 503668 57598
rect 503720 57588 503772 57594
rect 503720 57530 503772 57536
rect 502432 4072 502484 4078
rect 502432 4014 502484 4020
rect 503628 4072 503680 4078
rect 503628 4014 503680 4020
rect 501052 604 501104 610
rect 501052 546 501104 552
rect 501236 604 501288 610
rect 501236 546 501288 552
rect 501248 480 501276 546
rect 502444 480 502472 4014
rect 503628 3188 503680 3194
rect 503628 3130 503680 3136
rect 503640 480 503668 3130
rect 503732 610 503760 57530
rect 504100 56710 504128 60030
rect 504088 56704 504140 56710
rect 504088 56646 504140 56652
rect 505020 5166 505048 60030
rect 505664 57662 505692 60044
rect 505652 57656 505704 57662
rect 505652 57598 505704 57604
rect 506388 57656 506440 57662
rect 506388 57598 506440 57604
rect 505008 5160 505060 5166
rect 505008 5102 505060 5108
rect 506020 3256 506072 3262
rect 506020 3198 506072 3204
rect 503720 604 503772 610
rect 503720 546 503772 552
rect 504824 604 504876 610
rect 504824 546 504876 552
rect 504836 480 504864 546
rect 506032 480 506060 3198
rect 506400 3194 506428 57598
rect 506676 57594 506704 60044
rect 506664 57588 506716 57594
rect 506664 57530 506716 57536
rect 507596 57458 507624 60044
rect 508622 60030 509188 60058
rect 507952 57520 508004 57526
rect 507952 57462 508004 57468
rect 507584 57452 507636 57458
rect 507584 57394 507636 57400
rect 507216 4004 507268 4010
rect 507216 3946 507268 3952
rect 506388 3188 506440 3194
rect 506388 3130 506440 3136
rect 507228 480 507256 3946
rect 507964 610 507992 57462
rect 509160 3126 509188 60030
rect 509528 57526 509556 60044
rect 509516 57520 509568 57526
rect 509516 57462 509568 57468
rect 509884 56704 509936 56710
rect 509884 56646 509936 56652
rect 509608 3324 509660 3330
rect 509608 3266 509660 3272
rect 509148 3120 509200 3126
rect 509148 3062 509200 3068
rect 507952 604 508004 610
rect 507952 546 508004 552
rect 508412 604 508464 610
rect 508412 546 508464 552
rect 508424 480 508452 546
rect 509620 480 509648 3266
rect 509896 3058 509924 56646
rect 510540 5098 510568 60044
rect 511566 60030 511948 60058
rect 510528 5092 510580 5098
rect 510528 5034 510580 5040
rect 511920 3058 511948 60030
rect 512472 57730 512500 60044
rect 512460 57724 512512 57730
rect 512460 57666 512512 57672
rect 513484 57662 513512 60044
rect 514510 60030 514708 60058
rect 513472 57656 513524 57662
rect 513472 57598 513524 57604
rect 514576 57656 514628 57662
rect 514576 57598 514628 57604
rect 512092 57248 512144 57254
rect 512092 57190 512144 57196
rect 509884 3052 509936 3058
rect 509884 2994 509936 3000
rect 511908 3052 511960 3058
rect 511908 2994 511960 3000
rect 510804 2848 510856 2854
rect 510804 2790 510856 2796
rect 510816 480 510844 2790
rect 512104 626 512132 57190
rect 514588 5030 514616 57598
rect 514576 5024 514628 5030
rect 514576 4966 514628 4972
rect 514680 4146 514708 60030
rect 515416 57662 515444 60044
rect 515404 57656 515456 57662
rect 515404 57598 515456 57604
rect 516428 57390 516456 60044
rect 514760 57384 514812 57390
rect 514760 57326 514812 57332
rect 516416 57384 516468 57390
rect 516416 57326 516468 57332
rect 514392 4140 514444 4146
rect 514392 4082 514444 4088
rect 514668 4140 514720 4146
rect 514668 4082 514720 4088
rect 513196 3392 513248 3398
rect 513196 3334 513248 3340
rect 512012 598 512132 626
rect 512012 480 512040 598
rect 513208 480 513236 3334
rect 514404 480 514432 4082
rect 514772 610 514800 57326
rect 516784 3800 516836 3806
rect 516784 3742 516836 3748
rect 514760 604 514812 610
rect 514760 546 514812 552
rect 515588 604 515640 610
rect 515588 546 515640 552
rect 515600 480 515628 546
rect 516796 480 516824 3742
rect 517440 3398 517468 60044
rect 518374 60030 518848 60058
rect 517428 3392 517480 3398
rect 517428 3334 517480 3340
rect 518820 3330 518848 60030
rect 519372 57866 519400 60044
rect 520384 57866 520412 60044
rect 521318 60030 521516 60058
rect 522330 60030 522988 60058
rect 519360 57860 519412 57866
rect 519360 57802 519412 57808
rect 520188 57860 520240 57866
rect 520188 57802 520240 57808
rect 520372 57860 520424 57866
rect 520372 57802 520424 57808
rect 520200 4962 520228 57802
rect 521384 5500 521436 5506
rect 521384 5442 521436 5448
rect 520188 4956 520240 4962
rect 520188 4898 520240 4904
rect 519084 4820 519136 4826
rect 519084 4762 519136 4768
rect 518808 3324 518860 3330
rect 518808 3266 518860 3272
rect 517888 2916 517940 2922
rect 517888 2858 517940 2864
rect 517900 480 517928 2858
rect 519096 480 519124 4762
rect 520280 3732 520332 3738
rect 520280 3674 520332 3680
rect 520292 480 520320 3674
rect 521396 3262 521424 5442
rect 521488 5386 521516 60030
rect 521568 57860 521620 57866
rect 521568 57802 521620 57808
rect 521580 5506 521608 57802
rect 521660 57112 521712 57118
rect 521660 57054 521712 57060
rect 521568 5500 521620 5506
rect 521568 5442 521620 5448
rect 521488 5358 521608 5386
rect 521476 3868 521528 3874
rect 521476 3810 521528 3816
rect 521384 3256 521436 3262
rect 521384 3198 521436 3204
rect 521488 480 521516 3810
rect 521580 3806 521608 5358
rect 521568 3800 521620 3806
rect 521568 3742 521620 3748
rect 521672 610 521700 57054
rect 522960 4894 522988 60030
rect 523328 56710 523356 60044
rect 523316 56704 523368 56710
rect 523316 56646 523368 56652
rect 522948 4888 523000 4894
rect 522948 4830 523000 4836
rect 524248 3738 524276 60044
rect 525260 57254 525288 60044
rect 525800 57316 525852 57322
rect 525800 57258 525852 57264
rect 525248 57248 525300 57254
rect 525248 57190 525300 57196
rect 524328 56704 524380 56710
rect 524328 56646 524380 56652
rect 524340 3874 524368 56646
rect 525064 3936 525116 3942
rect 525064 3878 525116 3884
rect 524328 3868 524380 3874
rect 524328 3810 524380 3816
rect 524236 3732 524288 3738
rect 524236 3674 524288 3680
rect 523868 3664 523920 3670
rect 523868 3606 523920 3612
rect 521660 604 521712 610
rect 521660 546 521712 552
rect 522672 604 522724 610
rect 522672 546 522724 552
rect 522684 480 522712 546
rect 523880 480 523908 3606
rect 525076 480 525104 3878
rect 525812 610 525840 57258
rect 526180 57118 526208 60044
rect 527192 57866 527220 60044
rect 527180 57860 527232 57866
rect 527180 57802 527232 57808
rect 528204 57322 528232 60044
rect 528468 57860 528520 57866
rect 528468 57802 528520 57808
rect 528192 57316 528244 57322
rect 528192 57258 528244 57264
rect 526444 57180 526496 57186
rect 526444 57122 526496 57128
rect 526168 57112 526220 57118
rect 526168 57054 526220 57060
rect 526456 4010 526484 57122
rect 526444 4004 526496 4010
rect 526444 3946 526496 3952
rect 528480 3942 528508 57802
rect 529124 57186 529152 60044
rect 529204 57928 529256 57934
rect 529204 57870 529256 57876
rect 529112 57180 529164 57186
rect 529112 57122 529164 57128
rect 528744 57044 528796 57050
rect 528744 56986 528796 56992
rect 528652 4004 528704 4010
rect 528652 3946 528704 3952
rect 528468 3936 528520 3942
rect 528468 3878 528520 3884
rect 527456 3528 527508 3534
rect 527456 3470 527508 3476
rect 525800 604 525852 610
rect 525800 546 525852 552
rect 526260 604 526312 610
rect 526260 546 526312 552
rect 526272 480 526300 546
rect 527468 480 527496 3470
rect 528664 480 528692 3946
rect 528756 3346 528784 56986
rect 529216 3602 529244 57870
rect 530136 57798 530164 60044
rect 530124 57792 530176 57798
rect 530124 57734 530176 57740
rect 531148 4826 531176 60044
rect 532082 60030 532648 60058
rect 531228 57792 531280 57798
rect 531228 57734 531280 57740
rect 531136 4820 531188 4826
rect 531136 4762 531188 4768
rect 531240 4078 531268 57734
rect 531228 4072 531280 4078
rect 531228 4014 531280 4020
rect 532620 3670 532648 60030
rect 533080 57866 533108 60044
rect 532700 57860 532752 57866
rect 532700 57802 532752 57808
rect 533068 57860 533120 57866
rect 533068 57802 533120 57808
rect 532608 3664 532660 3670
rect 532608 3606 532660 3612
rect 529204 3596 529256 3602
rect 529204 3538 529256 3544
rect 532240 3596 532292 3602
rect 532240 3538 532292 3544
rect 528756 3318 529888 3346
rect 529860 480 529888 3318
rect 531044 2984 531096 2990
rect 531044 2926 531096 2932
rect 531056 480 531084 2926
rect 532252 480 532280 3538
rect 532712 2802 532740 57802
rect 534092 57798 534120 60044
rect 534080 57792 534132 57798
rect 534080 57734 534132 57740
rect 533344 57112 533396 57118
rect 533344 57054 533396 57060
rect 533356 2990 533384 57054
rect 535012 56982 535040 60044
rect 535368 57792 535420 57798
rect 535368 57734 535420 57740
rect 535000 56976 535052 56982
rect 535000 56918 535052 56924
rect 535380 3602 535408 57734
rect 536024 56846 536052 60044
rect 537036 57866 537064 60044
rect 537024 57860 537076 57866
rect 537024 57802 537076 57808
rect 537484 57180 537536 57186
rect 537484 57122 537536 57128
rect 536012 56840 536064 56846
rect 536012 56782 536064 56788
rect 536748 56840 536800 56846
rect 536748 56782 536800 56788
rect 535368 3596 535420 3602
rect 535368 3538 535420 3544
rect 536760 3534 536788 56782
rect 536932 5228 536984 5234
rect 536932 5170 536984 5176
rect 534540 3528 534592 3534
rect 534540 3470 534592 3476
rect 536748 3528 536800 3534
rect 536748 3470 536800 3476
rect 533344 2984 533396 2990
rect 533344 2926 533396 2932
rect 532712 2774 533476 2802
rect 533448 480 533476 2774
rect 534552 480 534580 3470
rect 535736 3460 535788 3466
rect 535736 3402 535788 3408
rect 535748 480 535776 3402
rect 536944 480 536972 5170
rect 537496 2922 537524 57122
rect 537956 56642 537984 60044
rect 537944 56636 537996 56642
rect 537944 56578 537996 56584
rect 538048 22098 538076 659246
rect 538416 627881 538444 660962
rect 538496 660952 538548 660958
rect 538496 660894 538548 660900
rect 538402 627872 538458 627881
rect 538402 627807 538458 627816
rect 538508 580990 538536 660894
rect 538588 660884 538640 660890
rect 538588 660826 538640 660832
rect 538496 580984 538548 580990
rect 538496 580926 538548 580932
rect 538600 534070 538628 660826
rect 538680 660816 538732 660822
rect 538680 660758 538732 660764
rect 538588 534064 538640 534070
rect 538588 534006 538640 534012
rect 538692 487150 538720 660758
rect 538680 487144 538732 487150
rect 538680 487086 538732 487092
rect 538784 393310 538812 661710
rect 539508 660612 539560 660618
rect 539508 660554 539560 660560
rect 539230 660104 539286 660113
rect 539230 660039 539286 660048
rect 539140 660000 539192 660006
rect 539046 659968 539102 659977
rect 539140 659942 539192 659948
rect 539046 659903 539102 659912
rect 538862 659696 538918 659705
rect 538862 659631 538918 659640
rect 538772 393304 538824 393310
rect 538772 393246 538824 393252
rect 538128 57860 538180 57866
rect 538128 57802 538180 57808
rect 538036 22092 538088 22098
rect 538036 22034 538088 22040
rect 538140 3466 538168 57802
rect 538876 17950 538904 659631
rect 538954 658472 539010 658481
rect 538954 658407 539010 658416
rect 538968 88330 538996 658407
rect 538956 88324 539008 88330
rect 538956 88266 539008 88272
rect 539060 64870 539088 659903
rect 539152 158710 539180 659942
rect 539140 158704 539192 158710
rect 539140 158646 539192 158652
rect 539244 111790 539272 660039
rect 539416 658980 539468 658986
rect 539416 658922 539468 658928
rect 539324 658776 539376 658782
rect 539324 658718 539376 658724
rect 539336 252550 539364 658718
rect 539428 299470 539456 658922
rect 539520 346390 539548 660554
rect 539692 659524 539744 659530
rect 539692 659466 539744 659472
rect 539704 651370 539732 659466
rect 539784 659388 539836 659394
rect 539784 659330 539836 659336
rect 539692 651364 539744 651370
rect 539692 651306 539744 651312
rect 539600 627904 539652 627910
rect 539598 627872 539600 627881
rect 539652 627872 539654 627881
rect 539598 627807 539654 627816
rect 539796 604450 539824 659330
rect 539784 604444 539836 604450
rect 539784 604386 539836 604392
rect 539888 557530 539916 662730
rect 539968 662720 540020 662726
rect 539968 662662 540020 662668
rect 539876 557524 539928 557530
rect 539876 557466 539928 557472
rect 539980 510610 540008 662662
rect 577504 662516 577556 662522
rect 577504 662458 577556 662464
rect 540060 662040 540112 662046
rect 540060 661982 540112 661988
rect 539968 510604 540020 510610
rect 539968 510546 540020 510552
rect 540072 499526 540100 661982
rect 541716 661972 541768 661978
rect 541716 661914 541768 661920
rect 541624 661904 541676 661910
rect 541624 661846 541676 661852
rect 540888 661836 540940 661842
rect 540888 661778 540940 661784
rect 540796 661700 540848 661706
rect 540796 661642 540848 661648
rect 540612 661496 540664 661502
rect 540612 661438 540664 661444
rect 540244 661224 540296 661230
rect 540244 661166 540296 661172
rect 540152 659252 540204 659258
rect 540152 659194 540204 659200
rect 540060 499520 540112 499526
rect 540060 499462 540112 499468
rect 540164 463690 540192 659194
rect 540152 463684 540204 463690
rect 540152 463626 540204 463632
rect 539508 346384 539560 346390
rect 539508 346326 539560 346332
rect 539416 299464 539468 299470
rect 539416 299406 539468 299412
rect 539324 252544 539376 252550
rect 539324 252486 539376 252492
rect 540256 182170 540284 661166
rect 540428 660272 540480 660278
rect 540428 660214 540480 660220
rect 540336 658640 540388 658646
rect 540336 658582 540388 658588
rect 540348 229090 540376 658582
rect 540440 264926 540468 660214
rect 540520 658844 540572 658850
rect 540520 658786 540572 658792
rect 540532 276010 540560 658786
rect 540624 311846 540652 661438
rect 540704 661428 540756 661434
rect 540704 661370 540756 661376
rect 540716 322930 540744 661370
rect 540808 369850 540836 661642
rect 540900 416770 540928 661778
rect 540888 416764 540940 416770
rect 540888 416706 540940 416712
rect 541636 405686 541664 661846
rect 541728 452606 541756 661914
rect 548524 661632 548576 661638
rect 548524 661574 548576 661580
rect 541900 659592 541952 659598
rect 541900 659534 541952 659540
rect 541808 659456 541860 659462
rect 541808 659398 541860 659404
rect 541820 593366 541848 659398
rect 541912 640286 541940 659534
rect 541900 640280 541952 640286
rect 541900 640222 541952 640228
rect 541808 593360 541860 593366
rect 541808 593302 541860 593308
rect 541716 452600 541768 452606
rect 541716 452542 541768 452548
rect 541624 405680 541676 405686
rect 541624 405622 541676 405628
rect 540796 369844 540848 369850
rect 540796 369786 540848 369792
rect 548536 358766 548564 661574
rect 577516 440230 577544 662458
rect 580262 661600 580318 661609
rect 580262 661535 580318 661544
rect 580172 659116 580224 659122
rect 580172 659058 580224 659064
rect 580080 651364 580132 651370
rect 580080 651306 580132 651312
rect 580092 651137 580120 651306
rect 580078 651128 580134 651137
rect 580078 651063 580134 651072
rect 580080 640280 580132 640286
rect 580080 640222 580132 640228
rect 580092 639441 580120 640222
rect 580078 639432 580134 639441
rect 580078 639367 580134 639376
rect 580080 627904 580132 627910
rect 580080 627846 580132 627852
rect 580092 627745 580120 627846
rect 580078 627736 580134 627745
rect 580078 627671 580134 627680
rect 580080 604444 580132 604450
rect 580080 604386 580132 604392
rect 580092 604217 580120 604386
rect 580078 604208 580134 604217
rect 580078 604143 580134 604152
rect 580080 593360 580132 593366
rect 580080 593302 580132 593308
rect 580092 592521 580120 593302
rect 580078 592512 580134 592521
rect 580078 592447 580134 592456
rect 580080 580984 580132 580990
rect 580080 580926 580132 580932
rect 580092 580825 580120 580926
rect 580078 580816 580134 580825
rect 580078 580751 580134 580760
rect 580080 557524 580132 557530
rect 580080 557466 580132 557472
rect 580092 557297 580120 557466
rect 580078 557288 580134 557297
rect 580078 557223 580134 557232
rect 580184 545601 580212 659058
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580172 534064 580224 534070
rect 580172 534006 580224 534012
rect 580184 533905 580212 534006
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 579804 510604 579856 510610
rect 579804 510546 579856 510552
rect 579816 510377 579844 510546
rect 579802 510368 579858 510377
rect 579802 510303 579858 510312
rect 579988 499520 580040 499526
rect 579988 499462 580040 499468
rect 580000 498681 580028 499462
rect 579986 498672 580042 498681
rect 579986 498607 580042 498616
rect 580172 487144 580224 487150
rect 580172 487086 580224 487092
rect 580184 486849 580212 487086
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 579804 463684 579856 463690
rect 579804 463626 579856 463632
rect 579816 463457 579844 463626
rect 579802 463448 579858 463457
rect 579802 463383 579858 463392
rect 579988 452600 580040 452606
rect 579988 452542 580040 452548
rect 580000 451761 580028 452542
rect 579986 451752 580042 451761
rect 579986 451687 580042 451696
rect 577504 440224 577556 440230
rect 577504 440166 577556 440172
rect 579712 440224 579764 440230
rect 579712 440166 579764 440172
rect 579724 439929 579752 440166
rect 579710 439920 579766 439929
rect 579710 439855 579766 439864
rect 579804 416764 579856 416770
rect 579804 416706 579856 416712
rect 579816 416537 579844 416706
rect 579802 416528 579858 416537
rect 579802 416463 579858 416472
rect 579988 405680 580040 405686
rect 579988 405622 580040 405628
rect 580000 404841 580028 405622
rect 579986 404832 580042 404841
rect 579986 404767 580042 404776
rect 580172 393304 580224 393310
rect 580172 393246 580224 393252
rect 580184 393009 580212 393246
rect 580170 393000 580226 393009
rect 580170 392935 580226 392944
rect 579804 369844 579856 369850
rect 579804 369786 579856 369792
rect 579816 369617 579844 369786
rect 579802 369608 579858 369617
rect 579802 369543 579858 369552
rect 548524 358760 548576 358766
rect 548524 358702 548576 358708
rect 579988 358760 580040 358766
rect 579988 358702 580040 358708
rect 580000 357921 580028 358702
rect 579986 357912 580042 357921
rect 579986 357847 580042 357856
rect 580172 346384 580224 346390
rect 580172 346326 580224 346332
rect 580184 346089 580212 346326
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 540704 322924 540756 322930
rect 540704 322866 540756 322872
rect 579804 322924 579856 322930
rect 579804 322866 579856 322872
rect 579816 322697 579844 322866
rect 579802 322688 579858 322697
rect 579802 322623 579858 322632
rect 540612 311840 540664 311846
rect 540612 311782 540664 311788
rect 579988 311840 580040 311846
rect 579988 311782 580040 311788
rect 580000 310865 580028 311782
rect 579986 310856 580042 310865
rect 579986 310791 580042 310800
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 299169 580212 299406
rect 580170 299160 580226 299169
rect 580170 299095 580226 299104
rect 540520 276004 540572 276010
rect 540520 275946 540572 275952
rect 579804 276004 579856 276010
rect 579804 275946 579856 275952
rect 579816 275777 579844 275946
rect 579802 275768 579858 275777
rect 579802 275703 579858 275712
rect 540428 264920 540480 264926
rect 540428 264862 540480 264868
rect 579988 264920 580040 264926
rect 579988 264862 580040 264868
rect 580000 263945 580028 264862
rect 579986 263936 580042 263945
rect 579986 263871 580042 263880
rect 580172 252544 580224 252550
rect 580172 252486 580224 252492
rect 580184 252249 580212 252486
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 540336 229084 540388 229090
rect 540336 229026 540388 229032
rect 579804 229084 579856 229090
rect 579804 229026 579856 229032
rect 579816 228857 579844 229026
rect 579802 228848 579858 228857
rect 579802 228783 579858 228792
rect 540244 182164 540296 182170
rect 540244 182106 540296 182112
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 580172 158704 580224 158710
rect 580172 158646 580224 158652
rect 580184 158409 580212 158646
rect 580170 158400 580226 158409
rect 580170 158335 580226 158344
rect 539232 111784 539284 111790
rect 539232 111726 539284 111732
rect 580172 111784 580224 111790
rect 580172 111726 580224 111732
rect 580184 111489 580212 111726
rect 580170 111480 580226 111489
rect 580170 111415 580226 111424
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 539048 64864 539100 64870
rect 539048 64806 539100 64812
rect 579620 64864 579672 64870
rect 579620 64806 579672 64812
rect 579632 64569 579660 64806
rect 579618 64560 579674 64569
rect 579618 64495 579674 64504
rect 538968 57594 538996 60044
rect 541624 57792 541676 57798
rect 541624 57734 541676 57740
rect 538956 57588 539008 57594
rect 538956 57530 539008 57536
rect 538956 56976 539008 56982
rect 538956 56918 539008 56924
rect 538864 17944 538916 17950
rect 538864 17886 538916 17892
rect 538968 4078 538996 56918
rect 540244 56636 540296 56642
rect 540244 56578 540296 56584
rect 538956 4072 539008 4078
rect 538956 4014 539008 4020
rect 538036 3460 538088 3466
rect 538036 3402 538088 3408
rect 538128 3460 538180 3466
rect 538128 3402 538180 3408
rect 538048 3346 538076 3402
rect 540256 3369 540284 56578
rect 540520 5160 540572 5166
rect 540520 5102 540572 5108
rect 540242 3360 540298 3369
rect 538048 3318 538168 3346
rect 537484 2916 537536 2922
rect 537484 2858 537536 2864
rect 538140 480 538168 3318
rect 540242 3295 540298 3304
rect 539324 2848 539376 2854
rect 539324 2790 539376 2796
rect 539336 480 539364 2790
rect 540532 480 540560 5102
rect 541636 4978 541664 57734
rect 547144 57724 547196 57730
rect 547144 57666 547196 57672
rect 544384 57588 544436 57594
rect 544384 57530 544436 57536
rect 542360 57520 542412 57526
rect 542360 57462 542412 57468
rect 541636 4950 541940 4978
rect 541912 3194 541940 4950
rect 541716 3188 541768 3194
rect 541716 3130 541768 3136
rect 541900 3188 541952 3194
rect 541900 3130 541952 3136
rect 541728 480 541756 3130
rect 542372 610 542400 57462
rect 543740 57452 543792 57458
rect 543740 57394 543792 57400
rect 543752 610 543780 57394
rect 544396 2990 544424 57530
rect 545764 57180 545816 57186
rect 545764 57122 545816 57128
rect 545776 3194 545804 57122
rect 547156 3194 547184 57666
rect 549904 57656 549956 57662
rect 549904 57598 549956 57604
rect 547696 5092 547748 5098
rect 547696 5034 547748 5040
rect 545764 3188 545816 3194
rect 545764 3130 545816 3136
rect 546500 3188 546552 3194
rect 546500 3130 546552 3136
rect 547144 3188 547196 3194
rect 547144 3130 547196 3136
rect 545304 3120 545356 3126
rect 545304 3062 545356 3068
rect 544384 2984 544436 2990
rect 544384 2926 544436 2932
rect 542360 604 542412 610
rect 542360 546 542412 552
rect 542912 604 542964 610
rect 542912 546 542964 552
rect 543740 604 543792 610
rect 543740 546 543792 552
rect 544108 604 544160 610
rect 544108 546 544160 552
rect 542924 480 542952 546
rect 544120 480 544148 546
rect 545316 480 545344 3062
rect 546512 480 546540 3130
rect 547708 480 547736 5034
rect 549916 3398 549944 57598
rect 554872 57384 554924 57390
rect 554872 57326 554924 57332
rect 551192 5024 551244 5030
rect 551192 4966 551244 4972
rect 549904 3392 549956 3398
rect 549904 3334 549956 3340
rect 550088 3188 550140 3194
rect 550088 3130 550140 3136
rect 548892 3052 548944 3058
rect 548892 2994 548944 3000
rect 548904 480 548932 2994
rect 550100 480 550128 3130
rect 551204 480 551232 4966
rect 552388 4140 552440 4146
rect 552388 4082 552440 4088
rect 552400 480 552428 4082
rect 554884 3482 554912 57326
rect 566464 57316 566516 57322
rect 566464 57258 566516 57264
rect 564440 57248 564492 57254
rect 564440 57190 564492 57196
rect 558368 4956 558420 4962
rect 558368 4898 558420 4904
rect 554792 3454 554912 3482
rect 553584 3392 553636 3398
rect 553584 3334 553636 3340
rect 553596 480 553624 3334
rect 554792 480 554820 3454
rect 557172 3324 557224 3330
rect 557172 3266 557224 3272
rect 555976 3052 556028 3058
rect 555976 2994 556028 3000
rect 555988 480 556016 2994
rect 557184 480 557212 3266
rect 558380 480 558408 4898
rect 561956 4888 562008 4894
rect 561956 4830 562008 4836
rect 560760 3800 560812 3806
rect 560760 3742 560812 3748
rect 559564 3256 559616 3262
rect 559564 3198 559616 3204
rect 559576 480 559604 3198
rect 560772 480 560800 3742
rect 561968 480 561996 4830
rect 563152 4004 563204 4010
rect 563152 3946 563204 3952
rect 563164 480 563192 3946
rect 564348 3868 564400 3874
rect 564348 3810 564400 3816
rect 564360 480 564388 3810
rect 564452 3482 564480 57190
rect 566476 4146 566504 57258
rect 580276 29345 580304 661535
rect 580446 661464 580502 661473
rect 580446 661399 580502 661408
rect 580354 659152 580410 659161
rect 580354 659087 580410 659096
rect 580368 76265 580396 659087
rect 580354 76256 580410 76265
rect 580354 76191 580410 76200
rect 580460 41041 580488 661399
rect 580724 660408 580776 660414
rect 580724 660350 580776 660356
rect 580538 660240 580594 660249
rect 580538 660175 580594 660184
rect 580552 123185 580580 660175
rect 580632 659320 580684 659326
rect 580632 659262 580684 659268
rect 580644 134881 580672 659262
rect 580736 170105 580764 660350
rect 580908 660340 580960 660346
rect 580908 660282 580960 660288
rect 580816 659184 580868 659190
rect 580816 659126 580868 659132
rect 580828 205329 580856 659126
rect 580920 217025 580948 660282
rect 580906 217016 580962 217025
rect 580906 216951 580962 216960
rect 580814 205320 580870 205329
rect 580814 205255 580870 205264
rect 580722 170096 580778 170105
rect 580722 170031 580778 170040
rect 580630 134872 580686 134881
rect 580630 134807 580686 134816
rect 580538 123176 580594 123185
rect 580538 123111 580594 123120
rect 580446 41032 580502 41041
rect 580446 40967 580502 40976
rect 580262 29336 580318 29345
rect 580262 29271 580318 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 572628 4820 572680 4826
rect 572628 4762 572680 4768
rect 566464 4140 566516 4146
rect 566464 4082 566516 4088
rect 569040 4140 569092 4146
rect 569040 4082 569092 4088
rect 567844 3936 567896 3942
rect 567844 3878 567896 3884
rect 564452 3454 565584 3482
rect 565556 480 565584 3454
rect 566740 2916 566792 2922
rect 566740 2858 566792 2864
rect 566752 480 566780 2858
rect 567856 480 567884 3878
rect 569052 480 569080 4082
rect 571432 3732 571484 3738
rect 571432 3674 571484 3680
rect 570236 2848 570288 2854
rect 570236 2790 570288 2796
rect 570248 480 570276 2790
rect 571444 480 571472 3674
rect 572640 480 572668 4762
rect 577412 4072 577464 4078
rect 577412 4014 577464 4020
rect 573824 3664 573876 3670
rect 573824 3606 573876 3612
rect 573836 480 573864 3606
rect 576216 3596 576268 3602
rect 576216 3538 576268 3544
rect 575020 2984 575072 2990
rect 575020 2926 575072 2932
rect 575032 480 575060 2926
rect 576228 480 576256 3538
rect 577424 480 577452 4014
rect 578608 3528 578660 3534
rect 578608 3470 578660 3476
rect 578620 480 578648 3470
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 580998 3360 581054 3369
rect 580998 3295 581054 3304
rect 581012 480 581040 3295
rect 582196 3188 582248 3194
rect 582196 3130 582248 3136
rect 582208 480 582236 3130
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 8114 700304 8170 700360
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3974 661816 4030 661872
rect 3790 661680 3846 661736
rect 3606 661272 3662 661328
rect 3422 661000 3478 661056
rect 3146 653556 3148 653576
rect 3148 653556 3200 653576
rect 3200 653556 3202 653576
rect 3146 653520 3202 653556
rect 3146 624860 3148 624880
rect 3148 624860 3200 624880
rect 3200 624860 3202 624880
rect 3146 624824 3202 624860
rect 2778 610444 2780 610464
rect 2780 610444 2832 610464
rect 2832 610444 2834 610464
rect 2778 610408 2834 610444
rect 3146 596028 3148 596048
rect 3148 596028 3200 596048
rect 3200 596028 3202 596048
rect 3146 595992 3202 596028
rect 3146 567296 3202 567352
rect 3238 553016 3294 553072
rect 3238 538600 3294 538656
rect 3238 509904 3294 509960
rect 2778 495488 2834 495544
rect 3238 481072 3294 481128
rect 3238 452412 3240 452432
rect 3240 452412 3292 452432
rect 3292 452412 3294 452432
rect 3238 452376 3294 452412
rect 2778 437960 2834 438016
rect 3330 423680 3386 423736
rect 3330 394984 3386 395040
rect 3146 366152 3202 366208
rect 3330 337492 3332 337512
rect 3332 337492 3384 337512
rect 3384 337492 3386 337512
rect 3330 337456 3386 337492
rect 3054 308760 3110 308816
rect 3146 294344 3202 294400
rect 3330 280100 3332 280120
rect 3332 280100 3384 280120
rect 3384 280100 3386 280120
rect 3330 280064 3386 280100
rect 3330 265648 3386 265704
rect 3330 251232 3386 251288
rect 3330 236952 3386 237008
rect 3330 222536 3386 222592
rect 3330 208156 3332 208176
rect 3332 208156 3384 208176
rect 3384 208156 3386 208176
rect 3330 208120 3386 208156
rect 3330 193840 3386 193896
rect 3330 179424 3386 179480
rect 3054 165008 3110 165064
rect 3330 122032 3386 122088
rect 3330 93200 3386 93256
rect 3146 78920 3202 78976
rect 2778 64540 2780 64560
rect 2780 64540 2832 64560
rect 2832 64540 2834 64560
rect 2778 64504 2834 64540
rect 2870 21392 2926 21448
rect 3514 658960 3570 659016
rect 3698 658824 3754 658880
rect 3698 136312 3754 136368
rect 3882 323040 3938 323096
rect 4802 661136 4858 661192
rect 4066 380568 4122 380624
rect 3974 150728 4030 150784
rect 3790 107616 3846 107672
rect 9034 661952 9090 662008
rect 8942 658280 8998 658336
rect 58622 662088 58678 662144
rect 25502 659776 25558 659832
rect 69938 661544 69994 661600
rect 65706 661408 65762 661464
rect 74354 659912 74410 659968
rect 86774 660048 86830 660104
rect 61934 659640 61990 659696
rect 78586 659368 78642 659424
rect 155682 659368 155738 659424
rect 232594 660184 232650 660240
rect 356058 700304 356114 700360
rect 580170 697992 580226 698048
rect 494886 686024 494942 686080
rect 494242 685888 494298 685944
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 507766 662088 507822 662144
rect 482558 661952 482614 662008
rect 499394 661816 499450 661872
rect 511998 661680 512054 661736
rect 520462 661272 520518 661328
rect 524602 661136 524658 661192
rect 533066 661000 533122 661056
rect 503258 659776 503314 659832
rect 448518 659368 448574 659424
rect 457534 659368 457590 659424
rect 516138 659368 516194 659424
rect 5446 57160 5502 57216
rect 3606 50088 3662 50144
rect 3514 35808 3570 35864
rect 3422 7112 3478 7168
rect 55310 3612 55312 3632
rect 55312 3612 55364 3632
rect 55364 3612 55366 3632
rect 55310 3576 55366 3612
rect 63866 57160 63922 57216
rect 64694 3612 64696 3632
rect 64696 3612 64748 3632
rect 64748 3612 64750 3632
rect 64694 3576 64750 3612
rect 99102 58112 99158 58168
rect 98458 57976 98514 58032
rect 98274 29008 98330 29064
rect 98458 29008 98514 29064
rect 115294 57160 115350 57216
rect 127530 57160 127586 57216
rect 146206 57160 146262 57216
rect 179418 57160 179474 57216
rect 195886 19216 195942 19272
rect 195886 9696 195942 9752
rect 196162 19216 196218 19272
rect 196162 9696 196218 9752
rect 202786 57160 202842 57216
rect 226430 57160 226486 57216
rect 334070 18128 334126 18184
rect 333978 17992 334034 18048
rect 448334 3068 448336 3088
rect 448336 3068 448388 3088
rect 448388 3068 448390 3088
rect 448334 3032 448390 3068
rect 451186 3052 451242 3088
rect 451186 3032 451188 3052
rect 451188 3032 451240 3052
rect 451240 3032 451242 3052
rect 456614 3304 456670 3360
rect 482282 3304 482338 3360
rect 538402 627816 538458 627872
rect 539230 660048 539286 660104
rect 539046 659912 539102 659968
rect 538862 659640 538918 659696
rect 538954 658416 539010 658472
rect 539598 627852 539600 627872
rect 539600 627852 539652 627872
rect 539652 627852 539654 627872
rect 539598 627816 539654 627852
rect 580262 661544 580318 661600
rect 580078 651072 580134 651128
rect 580078 639376 580134 639432
rect 580078 627680 580134 627736
rect 580078 604152 580134 604208
rect 580078 592456 580134 592512
rect 580078 580760 580134 580816
rect 580078 557232 580134 557288
rect 580170 545536 580226 545592
rect 580170 533840 580226 533896
rect 579802 510312 579858 510368
rect 579986 498616 580042 498672
rect 580170 486784 580226 486840
rect 579802 463392 579858 463448
rect 579986 451696 580042 451752
rect 579710 439864 579766 439920
rect 579802 416472 579858 416528
rect 579986 404776 580042 404832
rect 580170 392944 580226 393000
rect 579802 369552 579858 369608
rect 579986 357856 580042 357912
rect 580170 346024 580226 346080
rect 579802 322632 579858 322688
rect 579986 310800 580042 310856
rect 580170 299104 580226 299160
rect 579802 275712 579858 275768
rect 579986 263880 580042 263936
rect 580170 252184 580226 252240
rect 579802 228792 579858 228848
rect 580170 181872 580226 181928
rect 580170 158344 580226 158400
rect 580170 111424 580226 111480
rect 580170 87896 580226 87952
rect 579618 64504 579674 64560
rect 540242 3304 540298 3360
rect 580446 661408 580502 661464
rect 580354 659096 580410 659152
rect 580354 76200 580410 76256
rect 580538 660184 580594 660240
rect 580906 216960 580962 217016
rect 580814 205264 580870 205320
rect 580722 170040 580778 170096
rect 580630 134816 580686 134872
rect 580538 123120 580594 123176
rect 580446 40976 580502 41032
rect 580262 29280 580318 29336
rect 579802 17584 579858 17640
rect 580998 3304 581054 3360
<< metal3 >>
rect 8109 700362 8175 700365
rect 356053 700362 356119 700365
rect 8109 700360 356119 700362
rect 8109 700304 8114 700360
rect 8170 700304 356058 700360
rect 356114 700304 356119 700360
rect 8109 700302 356119 700304
rect 8109 700299 8175 700302
rect 356053 700299 356119 700302
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 494881 686082 494947 686085
rect 494102 686080 494947 686082
rect 494102 686024 494886 686080
rect 494942 686024 494947 686080
rect 494102 686022 494947 686024
rect 494102 685946 494162 686022
rect 494881 686019 494947 686022
rect 494237 685946 494303 685949
rect 494102 685944 494303 685946
rect 494102 685888 494242 685944
rect 494298 685888 494303 685944
rect 494102 685886 494303 685888
rect 494237 685883 494303 685886
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect 58617 662146 58683 662149
rect 507761 662146 507827 662149
rect 58617 662144 507827 662146
rect 58617 662088 58622 662144
rect 58678 662088 507766 662144
rect 507822 662088 507827 662144
rect 58617 662086 507827 662088
rect 58617 662083 58683 662086
rect 507761 662083 507827 662086
rect 9029 662010 9095 662013
rect 482553 662010 482619 662013
rect 9029 662008 482619 662010
rect 9029 661952 9034 662008
rect 9090 661952 482558 662008
rect 482614 661952 482619 662008
rect 9029 661950 482619 661952
rect 9029 661947 9095 661950
rect 482553 661947 482619 661950
rect 3969 661874 4035 661877
rect 499389 661874 499455 661877
rect 3969 661872 499455 661874
rect 3969 661816 3974 661872
rect 4030 661816 499394 661872
rect 499450 661816 499455 661872
rect 3969 661814 499455 661816
rect 3969 661811 4035 661814
rect 499389 661811 499455 661814
rect 3785 661738 3851 661741
rect 511993 661738 512059 661741
rect 3785 661736 512059 661738
rect 3785 661680 3790 661736
rect 3846 661680 511998 661736
rect 512054 661680 512059 661736
rect 3785 661678 512059 661680
rect 3785 661675 3851 661678
rect 511993 661675 512059 661678
rect 69933 661602 69999 661605
rect 580257 661602 580323 661605
rect 69933 661600 580323 661602
rect 69933 661544 69938 661600
rect 69994 661544 580262 661600
rect 580318 661544 580323 661600
rect 69933 661542 580323 661544
rect 69933 661539 69999 661542
rect 580257 661539 580323 661542
rect 65701 661466 65767 661469
rect 580441 661466 580507 661469
rect 65701 661464 580507 661466
rect 65701 661408 65706 661464
rect 65762 661408 580446 661464
rect 580502 661408 580507 661464
rect 65701 661406 580507 661408
rect 65701 661403 65767 661406
rect 580441 661403 580507 661406
rect 3601 661330 3667 661333
rect 520457 661330 520523 661333
rect 3601 661328 520523 661330
rect 3601 661272 3606 661328
rect 3662 661272 520462 661328
rect 520518 661272 520523 661328
rect 3601 661270 520523 661272
rect 3601 661267 3667 661270
rect 520457 661267 520523 661270
rect 4797 661194 4863 661197
rect 524597 661194 524663 661197
rect 4797 661192 524663 661194
rect 4797 661136 4802 661192
rect 4858 661136 524602 661192
rect 524658 661136 524663 661192
rect 4797 661134 524663 661136
rect 4797 661131 4863 661134
rect 524597 661131 524663 661134
rect 3417 661058 3483 661061
rect 533061 661058 533127 661061
rect 3417 661056 533127 661058
rect 3417 661000 3422 661056
rect 3478 661000 533066 661056
rect 533122 661000 533127 661056
rect 3417 660998 533127 661000
rect 3417 660995 3483 660998
rect 533061 660995 533127 660998
rect 232589 660242 232655 660245
rect 580533 660242 580599 660245
rect 232589 660240 580599 660242
rect 232589 660184 232594 660240
rect 232650 660184 580538 660240
rect 580594 660184 580599 660240
rect 232589 660182 580599 660184
rect 232589 660179 232655 660182
rect 580533 660179 580599 660182
rect 86769 660106 86835 660109
rect 539225 660106 539291 660109
rect 86769 660104 539291 660106
rect 86769 660048 86774 660104
rect 86830 660048 539230 660104
rect 539286 660048 539291 660104
rect 86769 660046 539291 660048
rect 86769 660043 86835 660046
rect 539225 660043 539291 660046
rect 74349 659970 74415 659973
rect 539041 659970 539107 659973
rect 74349 659968 539107 659970
rect 74349 659912 74354 659968
rect 74410 659912 539046 659968
rect 539102 659912 539107 659968
rect 74349 659910 539107 659912
rect 74349 659907 74415 659910
rect 539041 659907 539107 659910
rect 25497 659834 25563 659837
rect 503253 659834 503319 659837
rect 25497 659832 503319 659834
rect 25497 659776 25502 659832
rect 25558 659776 503258 659832
rect 503314 659776 503319 659832
rect 25497 659774 503319 659776
rect 25497 659771 25563 659774
rect 503253 659771 503319 659774
rect 61929 659698 61995 659701
rect 538857 659698 538923 659701
rect 61929 659696 538923 659698
rect 61929 659640 61934 659696
rect 61990 659640 538862 659696
rect 538918 659640 538923 659696
rect 61929 659638 538923 659640
rect 61929 659635 61995 659638
rect 538857 659635 538923 659638
rect 78581 659426 78647 659429
rect 81198 659426 81204 659428
rect 78581 659424 81204 659426
rect 78581 659368 78586 659424
rect 78642 659368 81204 659424
rect 78581 659366 81204 659368
rect 78581 659363 78647 659366
rect 81198 659364 81204 659366
rect 81268 659364 81274 659428
rect 155677 659426 155743 659429
rect 155677 659424 155786 659426
rect 155677 659368 155682 659424
rect 155738 659368 155786 659424
rect 155677 659363 155786 659368
rect 446438 659364 446444 659428
rect 446508 659426 446514 659428
rect 448513 659426 448579 659429
rect 446508 659424 448579 659426
rect 446508 659368 448518 659424
rect 448574 659368 448579 659424
rect 446508 659366 448579 659368
rect 446508 659364 446514 659366
rect 448513 659363 448579 659366
rect 456006 659364 456012 659428
rect 456076 659426 456082 659428
rect 457529 659426 457595 659429
rect 456076 659424 457595 659426
rect 456076 659368 457534 659424
rect 457590 659368 457595 659424
rect 456076 659366 457595 659368
rect 456076 659364 456082 659366
rect 457529 659363 457595 659366
rect 512678 659364 512684 659428
rect 512748 659426 512754 659428
rect 516133 659426 516199 659429
rect 512748 659424 516199 659426
rect 512748 659368 516138 659424
rect 516194 659368 516199 659424
rect 512748 659366 516199 659368
rect 512748 659364 512754 659366
rect 516133 659363 516199 659366
rect 155726 659154 155786 659363
rect 580349 659154 580415 659157
rect 155726 659152 580415 659154
rect 155726 659096 580354 659152
rect 580410 659096 580415 659152
rect 155726 659094 580415 659096
rect 580349 659091 580415 659094
rect 3509 659018 3575 659021
rect 446438 659018 446444 659020
rect 3509 659016 446444 659018
rect 3509 658960 3514 659016
rect 3570 658960 446444 659016
rect 3509 658958 446444 658960
rect 3509 658955 3575 658958
rect 446438 658956 446444 658958
rect 446508 658956 446514 659020
rect 3693 658882 3759 658885
rect 456006 658882 456012 658884
rect 3693 658880 456012 658882
rect 3693 658824 3698 658880
rect 3754 658824 456012 658880
rect 3693 658822 456012 658824
rect 3693 658819 3759 658822
rect 456006 658820 456012 658822
rect 456076 658820 456082 658884
rect 81198 658412 81204 658476
rect 81268 658474 81274 658476
rect 538949 658474 539015 658477
rect 81268 658472 539015 658474
rect 81268 658416 538954 658472
rect 539010 658416 539015 658472
rect 81268 658414 539015 658416
rect 81268 658412 81274 658414
rect 538949 658411 539015 658414
rect 8937 658338 9003 658341
rect 512678 658338 512684 658340
rect 8937 658336 512684 658338
rect 8937 658280 8942 658336
rect 8998 658280 512684 658336
rect 8937 658278 512684 658280
rect 8937 658275 9003 658278
rect 512678 658276 512684 658278
rect 512748 658276 512754 658340
rect -960 653578 480 653668
rect 3141 653578 3207 653581
rect -960 653576 3207 653578
rect -960 653520 3146 653576
rect 3202 653520 3207 653576
rect -960 653518 3207 653520
rect -960 653428 480 653518
rect 3141 653515 3207 653518
rect 580073 651130 580139 651133
rect 583520 651130 584960 651220
rect 580073 651128 584960 651130
rect 580073 651072 580078 651128
rect 580134 651072 584960 651128
rect 580073 651070 584960 651072
rect 580073 651067 580139 651070
rect 583520 650980 584960 651070
rect 580073 639434 580139 639437
rect 583520 639434 584960 639524
rect 580073 639432 584960 639434
rect 580073 639376 580078 639432
rect 580134 639376 584960 639432
rect 580073 639374 584960 639376
rect 580073 639371 580139 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 538397 627874 538463 627877
rect 539593 627874 539659 627877
rect 538397 627872 539659 627874
rect 538397 627816 538402 627872
rect 538458 627816 539598 627872
rect 539654 627816 539659 627872
rect 538397 627814 539659 627816
rect 538397 627811 538463 627814
rect 539593 627811 539659 627814
rect 580073 627738 580139 627741
rect 583520 627738 584960 627828
rect 580073 627736 584960 627738
rect 580073 627680 580078 627736
rect 580134 627680 584960 627736
rect 580073 627678 584960 627680
rect 580073 627675 580139 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3141 624882 3207 624885
rect -960 624880 3207 624882
rect -960 624824 3146 624880
rect 3202 624824 3207 624880
rect -960 624822 3207 624824
rect -960 624732 480 624822
rect 3141 624819 3207 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 2773 610466 2839 610469
rect -960 610464 2839 610466
rect -960 610408 2778 610464
rect 2834 610408 2839 610464
rect -960 610406 2839 610408
rect -960 610316 480 610406
rect 2773 610403 2839 610406
rect 580073 604210 580139 604213
rect 583520 604210 584960 604300
rect 580073 604208 584960 604210
rect 580073 604152 580078 604208
rect 580134 604152 584960 604208
rect 580073 604150 584960 604152
rect 580073 604147 580139 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3141 596050 3207 596053
rect -960 596048 3207 596050
rect -960 595992 3146 596048
rect 3202 595992 3207 596048
rect -960 595990 3207 595992
rect -960 595900 480 595990
rect 3141 595987 3207 595990
rect 580073 592514 580139 592517
rect 583520 592514 584960 592604
rect 580073 592512 584960 592514
rect 580073 592456 580078 592512
rect 580134 592456 584960 592512
rect 580073 592454 584960 592456
rect 580073 592451 580139 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580073 580818 580139 580821
rect 583520 580818 584960 580908
rect 580073 580816 584960 580818
rect 580073 580760 580078 580816
rect 580134 580760 584960 580816
rect 580073 580758 584960 580760
rect 580073 580755 580139 580758
rect 583520 580668 584960 580758
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3141 567354 3207 567357
rect -960 567352 3207 567354
rect -960 567296 3146 567352
rect 3202 567296 3207 567352
rect -960 567294 3207 567296
rect -960 567204 480 567294
rect 3141 567291 3207 567294
rect 580073 557290 580139 557293
rect 583520 557290 584960 557380
rect 580073 557288 584960 557290
rect 580073 557232 580078 557288
rect 580134 557232 584960 557288
rect 580073 557230 584960 557232
rect 580073 557227 580139 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3233 553074 3299 553077
rect -960 553072 3299 553074
rect -960 553016 3238 553072
rect 3294 553016 3299 553072
rect -960 553014 3299 553016
rect -960 552924 480 553014
rect 3233 553011 3299 553014
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect -960 538658 480 538748
rect 3233 538658 3299 538661
rect -960 538656 3299 538658
rect -960 538600 3238 538656
rect 3294 538600 3299 538656
rect -960 538598 3299 538600
rect -960 538508 480 538598
rect 3233 538595 3299 538598
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 579797 510370 579863 510373
rect 583520 510370 584960 510460
rect 579797 510368 584960 510370
rect 579797 510312 579802 510368
rect 579858 510312 584960 510368
rect 579797 510310 584960 510312
rect 579797 510307 579863 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3233 509962 3299 509965
rect -960 509960 3299 509962
rect -960 509904 3238 509960
rect 3294 509904 3299 509960
rect -960 509902 3299 509904
rect -960 509812 480 509902
rect 3233 509899 3299 509902
rect 579981 498674 580047 498677
rect 583520 498674 584960 498764
rect 579981 498672 584960 498674
rect 579981 498616 579986 498672
rect 580042 498616 584960 498672
rect 579981 498614 584960 498616
rect 579981 498611 580047 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 2773 495546 2839 495549
rect -960 495544 2839 495546
rect -960 495488 2778 495544
rect 2834 495488 2839 495544
rect -960 495486 2839 495488
rect -960 495396 480 495486
rect 2773 495483 2839 495486
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect -960 481130 480 481220
rect 3233 481130 3299 481133
rect -960 481128 3299 481130
rect -960 481072 3238 481128
rect 3294 481072 3299 481128
rect -960 481070 3299 481072
rect -960 480980 480 481070
rect 3233 481067 3299 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 579797 463450 579863 463453
rect 583520 463450 584960 463540
rect 579797 463448 584960 463450
rect 579797 463392 579802 463448
rect 579858 463392 584960 463448
rect 579797 463390 584960 463392
rect 579797 463387 579863 463390
rect 583520 463300 584960 463390
rect -960 452434 480 452524
rect 3233 452434 3299 452437
rect -960 452432 3299 452434
rect -960 452376 3238 452432
rect 3294 452376 3299 452432
rect -960 452374 3299 452376
rect -960 452284 480 452374
rect 3233 452371 3299 452374
rect 579981 451754 580047 451757
rect 583520 451754 584960 451844
rect 579981 451752 584960 451754
rect 579981 451696 579986 451752
rect 580042 451696 584960 451752
rect 579981 451694 584960 451696
rect 579981 451691 580047 451694
rect 583520 451604 584960 451694
rect 579705 439922 579771 439925
rect 583520 439922 584960 440012
rect 579705 439920 584960 439922
rect 579705 439864 579710 439920
rect 579766 439864 584960 439920
rect 579705 439862 584960 439864
rect 579705 439859 579771 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 2773 438018 2839 438021
rect -960 438016 2839 438018
rect -960 437960 2778 438016
rect 2834 437960 2839 438016
rect -960 437958 2839 437960
rect -960 437868 480 437958
rect 2773 437955 2839 437958
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3325 423738 3391 423741
rect -960 423736 3391 423738
rect -960 423680 3330 423736
rect 3386 423680 3391 423736
rect -960 423678 3391 423680
rect -960 423588 480 423678
rect 3325 423675 3391 423678
rect 579797 416530 579863 416533
rect 583520 416530 584960 416620
rect 579797 416528 584960 416530
rect 579797 416472 579802 416528
rect 579858 416472 584960 416528
rect 579797 416470 584960 416472
rect 579797 416467 579863 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 579981 404834 580047 404837
rect 583520 404834 584960 404924
rect 579981 404832 584960 404834
rect 579981 404776 579986 404832
rect 580042 404776 584960 404832
rect 579981 404774 584960 404776
rect 579981 404771 580047 404774
rect 583520 404684 584960 404774
rect -960 395042 480 395132
rect 3325 395042 3391 395045
rect -960 395040 3391 395042
rect -960 394984 3330 395040
rect 3386 394984 3391 395040
rect -960 394982 3391 394984
rect -960 394892 480 394982
rect 3325 394979 3391 394982
rect 580165 393002 580231 393005
rect 583520 393002 584960 393092
rect 580165 393000 584960 393002
rect 580165 392944 580170 393000
rect 580226 392944 584960 393000
rect 580165 392942 584960 392944
rect 580165 392939 580231 392942
rect 583520 392852 584960 392942
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 4061 380626 4127 380629
rect -960 380624 4127 380626
rect -960 380568 4066 380624
rect 4122 380568 4127 380624
rect -960 380566 4127 380568
rect -960 380476 480 380566
rect 4061 380563 4127 380566
rect 579797 369610 579863 369613
rect 583520 369610 584960 369700
rect 579797 369608 584960 369610
rect 579797 369552 579802 369608
rect 579858 369552 584960 369608
rect 579797 369550 584960 369552
rect 579797 369547 579863 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 3141 366210 3207 366213
rect -960 366208 3207 366210
rect -960 366152 3146 366208
rect 3202 366152 3207 366208
rect -960 366150 3207 366152
rect -960 366060 480 366150
rect 3141 366147 3207 366150
rect 579981 357914 580047 357917
rect 583520 357914 584960 358004
rect 579981 357912 584960 357914
rect 579981 357856 579986 357912
rect 580042 357856 584960 357912
rect 579981 357854 584960 357856
rect 579981 357851 580047 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect -960 337514 480 337604
rect 3325 337514 3391 337517
rect -960 337512 3391 337514
rect -960 337456 3330 337512
rect 3386 337456 3391 337512
rect -960 337454 3391 337456
rect -960 337364 480 337454
rect 3325 337451 3391 337454
rect 583520 334236 584960 334476
rect -960 323098 480 323188
rect 3877 323098 3943 323101
rect -960 323096 3943 323098
rect -960 323040 3882 323096
rect 3938 323040 3943 323096
rect -960 323038 3943 323040
rect -960 322948 480 323038
rect 3877 323035 3943 323038
rect 579797 322690 579863 322693
rect 583520 322690 584960 322780
rect 579797 322688 584960 322690
rect 579797 322632 579802 322688
rect 579858 322632 584960 322688
rect 579797 322630 584960 322632
rect 579797 322627 579863 322630
rect 583520 322540 584960 322630
rect 579981 310858 580047 310861
rect 583520 310858 584960 310948
rect 579981 310856 584960 310858
rect 579981 310800 579986 310856
rect 580042 310800 584960 310856
rect 579981 310798 584960 310800
rect 579981 310795 580047 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3049 308818 3115 308821
rect -960 308816 3115 308818
rect -960 308760 3054 308816
rect 3110 308760 3115 308816
rect -960 308758 3115 308760
rect -960 308668 480 308758
rect 3049 308755 3115 308758
rect 580165 299162 580231 299165
rect 583520 299162 584960 299252
rect 580165 299160 584960 299162
rect 580165 299104 580170 299160
rect 580226 299104 584960 299160
rect 580165 299102 584960 299104
rect 580165 299099 580231 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 3141 294402 3207 294405
rect -960 294400 3207 294402
rect -960 294344 3146 294400
rect 3202 294344 3207 294400
rect -960 294342 3207 294344
rect -960 294252 480 294342
rect 3141 294339 3207 294342
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 3325 280122 3391 280125
rect -960 280120 3391 280122
rect -960 280064 3330 280120
rect 3386 280064 3391 280120
rect -960 280062 3391 280064
rect -960 279972 480 280062
rect 3325 280059 3391 280062
rect 579797 275770 579863 275773
rect 583520 275770 584960 275860
rect 579797 275768 584960 275770
rect 579797 275712 579802 275768
rect 579858 275712 584960 275768
rect 579797 275710 584960 275712
rect 579797 275707 579863 275710
rect 583520 275620 584960 275710
rect -960 265706 480 265796
rect 3325 265706 3391 265709
rect -960 265704 3391 265706
rect -960 265648 3330 265704
rect 3386 265648 3391 265704
rect -960 265646 3391 265648
rect -960 265556 480 265646
rect 3325 265643 3391 265646
rect 579981 263938 580047 263941
rect 583520 263938 584960 264028
rect 579981 263936 584960 263938
rect 579981 263880 579986 263936
rect 580042 263880 584960 263936
rect 579981 263878 584960 263880
rect 579981 263875 580047 263878
rect 583520 263788 584960 263878
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3325 251290 3391 251293
rect -960 251288 3391 251290
rect -960 251232 3330 251288
rect 3386 251232 3391 251288
rect -960 251230 3391 251232
rect -960 251140 480 251230
rect 3325 251227 3391 251230
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 3325 237010 3391 237013
rect -960 237008 3391 237010
rect -960 236952 3330 237008
rect 3386 236952 3391 237008
rect -960 236950 3391 236952
rect -960 236860 480 236950
rect 3325 236947 3391 236950
rect 579797 228850 579863 228853
rect 583520 228850 584960 228940
rect 579797 228848 584960 228850
rect 579797 228792 579802 228848
rect 579858 228792 584960 228848
rect 579797 228790 584960 228792
rect 579797 228787 579863 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 3325 222594 3391 222597
rect -960 222592 3391 222594
rect -960 222536 3330 222592
rect 3386 222536 3391 222592
rect -960 222534 3391 222536
rect -960 222444 480 222534
rect 3325 222531 3391 222534
rect 580901 217018 580967 217021
rect 583520 217018 584960 217108
rect 580901 217016 584960 217018
rect 580901 216960 580906 217016
rect 580962 216960 584960 217016
rect 580901 216958 584960 216960
rect 580901 216955 580967 216958
rect 583520 216868 584960 216958
rect -960 208178 480 208268
rect 3325 208178 3391 208181
rect -960 208176 3391 208178
rect -960 208120 3330 208176
rect 3386 208120 3391 208176
rect -960 208118 3391 208120
rect -960 208028 480 208118
rect 3325 208115 3391 208118
rect 580809 205322 580875 205325
rect 583520 205322 584960 205412
rect 580809 205320 584960 205322
rect 580809 205264 580814 205320
rect 580870 205264 584960 205320
rect 580809 205262 584960 205264
rect 580809 205259 580875 205262
rect 583520 205172 584960 205262
rect -960 193898 480 193988
rect 3325 193898 3391 193901
rect -960 193896 3391 193898
rect -960 193840 3330 193896
rect 3386 193840 3391 193896
rect -960 193838 3391 193840
rect -960 193748 480 193838
rect 3325 193835 3391 193838
rect 583520 193476 584960 193716
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3325 179482 3391 179485
rect -960 179480 3391 179482
rect -960 179424 3330 179480
rect 3386 179424 3391 179480
rect -960 179422 3391 179424
rect -960 179332 480 179422
rect 3325 179419 3391 179422
rect 580717 170098 580783 170101
rect 583520 170098 584960 170188
rect 580717 170096 584960 170098
rect 580717 170040 580722 170096
rect 580778 170040 584960 170096
rect 580717 170038 584960 170040
rect 580717 170035 580783 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 3049 165066 3115 165069
rect -960 165064 3115 165066
rect -960 165008 3054 165064
rect 3110 165008 3115 165064
rect -960 165006 3115 165008
rect -960 164916 480 165006
rect 3049 165003 3115 165006
rect 580165 158402 580231 158405
rect 583520 158402 584960 158492
rect 580165 158400 584960 158402
rect 580165 158344 580170 158400
rect 580226 158344 584960 158400
rect 580165 158342 584960 158344
rect 580165 158339 580231 158342
rect 583520 158252 584960 158342
rect -960 150786 480 150876
rect 3969 150786 4035 150789
rect -960 150784 4035 150786
rect -960 150728 3974 150784
rect 4030 150728 4035 150784
rect -960 150726 4035 150728
rect -960 150636 480 150726
rect 3969 150723 4035 150726
rect 583520 146556 584960 146796
rect -960 136370 480 136460
rect 3693 136370 3759 136373
rect -960 136368 3759 136370
rect -960 136312 3698 136368
rect 3754 136312 3759 136368
rect -960 136310 3759 136312
rect -960 136220 480 136310
rect 3693 136307 3759 136310
rect 580625 134874 580691 134877
rect 583520 134874 584960 134964
rect 580625 134872 584960 134874
rect 580625 134816 580630 134872
rect 580686 134816 584960 134872
rect 580625 134814 584960 134816
rect 580625 134811 580691 134814
rect 583520 134724 584960 134814
rect 580533 123178 580599 123181
rect 583520 123178 584960 123268
rect 580533 123176 584960 123178
rect 580533 123120 580538 123176
rect 580594 123120 584960 123176
rect 580533 123118 584960 123120
rect 580533 123115 580599 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3325 122090 3391 122093
rect -960 122088 3391 122090
rect -960 122032 3330 122088
rect 3386 122032 3391 122088
rect -960 122030 3391 122032
rect -960 121940 480 122030
rect 3325 122027 3391 122030
rect 580165 111482 580231 111485
rect 583520 111482 584960 111572
rect 580165 111480 584960 111482
rect 580165 111424 580170 111480
rect 580226 111424 584960 111480
rect 580165 111422 584960 111424
rect 580165 111419 580231 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3785 107674 3851 107677
rect -960 107672 3851 107674
rect -960 107616 3790 107672
rect 3846 107616 3851 107672
rect -960 107614 3851 107616
rect -960 107524 480 107614
rect 3785 107611 3851 107614
rect 583520 99636 584960 99876
rect -960 93258 480 93348
rect 3325 93258 3391 93261
rect -960 93256 3391 93258
rect -960 93200 3330 93256
rect 3386 93200 3391 93256
rect -960 93198 3391 93200
rect -960 93108 480 93198
rect 3325 93195 3391 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect -960 78978 480 79068
rect 3141 78978 3207 78981
rect -960 78976 3207 78978
rect -960 78920 3146 78976
rect 3202 78920 3207 78976
rect -960 78918 3207 78920
rect -960 78828 480 78918
rect 3141 78915 3207 78918
rect 580349 76258 580415 76261
rect 583520 76258 584960 76348
rect 580349 76256 584960 76258
rect 580349 76200 580354 76256
rect 580410 76200 584960 76256
rect 580349 76198 584960 76200
rect 580349 76195 580415 76198
rect 583520 76108 584960 76198
rect -960 64562 480 64652
rect 2773 64562 2839 64565
rect -960 64560 2839 64562
rect -960 64504 2778 64560
rect 2834 64504 2839 64560
rect -960 64502 2839 64504
rect -960 64412 480 64502
rect 2773 64499 2839 64502
rect 579613 64562 579679 64565
rect 583520 64562 584960 64652
rect 579613 64560 584960 64562
rect 579613 64504 579618 64560
rect 579674 64504 584960 64560
rect 579613 64502 584960 64504
rect 579613 64499 579679 64502
rect 583520 64412 584960 64502
rect 99097 58170 99163 58173
rect 98318 58168 99163 58170
rect 98318 58112 99102 58168
rect 99158 58112 99163 58168
rect 98318 58110 99163 58112
rect 98318 58034 98378 58110
rect 99097 58107 99163 58110
rect 98453 58034 98519 58037
rect 98318 58032 98519 58034
rect 98318 57976 98458 58032
rect 98514 57976 98519 58032
rect 98318 57974 98519 57976
rect 98453 57971 98519 57974
rect 5441 57218 5507 57221
rect 63861 57218 63927 57221
rect 5441 57216 63927 57218
rect 5441 57160 5446 57216
rect 5502 57160 63866 57216
rect 63922 57160 63927 57216
rect 5441 57158 63927 57160
rect 5441 57155 5507 57158
rect 63861 57155 63927 57158
rect 115289 57218 115355 57221
rect 127525 57218 127591 57221
rect 115289 57216 127591 57218
rect 115289 57160 115294 57216
rect 115350 57160 127530 57216
rect 127586 57160 127591 57216
rect 115289 57158 127591 57160
rect 115289 57155 115355 57158
rect 127525 57155 127591 57158
rect 146201 57218 146267 57221
rect 179413 57218 179479 57221
rect 146201 57216 179479 57218
rect 146201 57160 146206 57216
rect 146262 57160 179418 57216
rect 179474 57160 179479 57216
rect 146201 57158 179479 57160
rect 146201 57155 146267 57158
rect 179413 57155 179479 57158
rect 202781 57218 202847 57221
rect 226425 57218 226491 57221
rect 202781 57216 226491 57218
rect 202781 57160 202786 57216
rect 202842 57160 226430 57216
rect 226486 57160 226491 57216
rect 202781 57158 226491 57160
rect 202781 57155 202847 57158
rect 226425 57155 226491 57158
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3601 50146 3667 50149
rect -960 50144 3667 50146
rect -960 50088 3606 50144
rect 3662 50088 3667 50144
rect -960 50086 3667 50088
rect -960 49996 480 50086
rect 3601 50083 3667 50086
rect 580441 41034 580507 41037
rect 583520 41034 584960 41124
rect 580441 41032 584960 41034
rect 580441 40976 580446 41032
rect 580502 40976 584960 41032
rect 580441 40974 584960 40976
rect 580441 40971 580507 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 3509 35866 3575 35869
rect -960 35864 3575 35866
rect -960 35808 3514 35864
rect 3570 35808 3575 35864
rect -960 35806 3575 35808
rect -960 35716 480 35806
rect 3509 35803 3575 35806
rect 580257 29338 580323 29341
rect 583520 29338 584960 29428
rect 580257 29336 584960 29338
rect 580257 29280 580262 29336
rect 580318 29280 584960 29336
rect 580257 29278 584960 29280
rect 580257 29275 580323 29278
rect 583520 29188 584960 29278
rect 98269 29066 98335 29069
rect 98453 29066 98519 29069
rect 98269 29064 98519 29066
rect 98269 29008 98274 29064
rect 98330 29008 98458 29064
rect 98514 29008 98519 29064
rect 98269 29006 98519 29008
rect 98269 29003 98335 29006
rect 98453 29003 98519 29006
rect -960 21450 480 21540
rect 2865 21450 2931 21453
rect -960 21448 2931 21450
rect -960 21392 2870 21448
rect 2926 21392 2931 21448
rect -960 21390 2931 21392
rect -960 21300 480 21390
rect 2865 21387 2931 21390
rect 195881 19274 195947 19277
rect 196157 19274 196223 19277
rect 195881 19272 196223 19274
rect 195881 19216 195886 19272
rect 195942 19216 196162 19272
rect 196218 19216 196223 19272
rect 195881 19214 196223 19216
rect 195881 19211 195947 19214
rect 196157 19211 196223 19214
rect 334065 18186 334131 18189
rect 333838 18184 334131 18186
rect 333838 18128 334070 18184
rect 334126 18128 334131 18184
rect 333838 18126 334131 18128
rect 333838 18050 333898 18126
rect 334065 18123 334131 18126
rect 333973 18050 334039 18053
rect 333838 18048 334039 18050
rect 333838 17992 333978 18048
rect 334034 17992 334039 18048
rect 333838 17990 334039 17992
rect 333973 17987 334039 17990
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect 195881 9754 195947 9757
rect 196157 9754 196223 9757
rect 195881 9752 196223 9754
rect 195881 9696 195886 9752
rect 195942 9696 196162 9752
rect 196218 9696 196223 9752
rect 195881 9694 196223 9696
rect 195881 9691 195947 9694
rect 196157 9691 196223 9694
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
rect 55305 3634 55371 3637
rect 64689 3634 64755 3637
rect 55305 3632 64755 3634
rect 55305 3576 55310 3632
rect 55366 3576 64694 3632
rect 64750 3576 64755 3632
rect 55305 3574 64755 3576
rect 55305 3571 55371 3574
rect 64689 3571 64755 3574
rect 456609 3362 456675 3365
rect 482277 3362 482343 3365
rect 456609 3360 482343 3362
rect 456609 3304 456614 3360
rect 456670 3304 482282 3360
rect 482338 3304 482343 3360
rect 456609 3302 482343 3304
rect 456609 3299 456675 3302
rect 482277 3299 482343 3302
rect 540237 3362 540303 3365
rect 580993 3362 581059 3365
rect 540237 3360 581059 3362
rect 540237 3304 540242 3360
rect 540298 3304 580998 3360
rect 581054 3304 581059 3360
rect 540237 3302 581059 3304
rect 540237 3299 540303 3302
rect 580993 3299 581059 3302
rect 448329 3090 448395 3093
rect 451181 3090 451247 3093
rect 448329 3088 451247 3090
rect 448329 3032 448334 3088
rect 448390 3032 451186 3088
rect 451242 3032 451247 3088
rect 448329 3030 451247 3032
rect 448329 3027 448395 3030
rect 451181 3027 451247 3030
<< via3 >>
rect 81204 659364 81268 659428
rect 446444 659364 446508 659428
rect 456012 659364 456076 659428
rect 512684 659364 512748 659428
rect 446444 658956 446508 659020
rect 456012 658820 456076 658884
rect 81204 658412 81268 658476
rect 512684 658276 512748 658340
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 672054 59004 707102
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 81203 659428 81269 659429
rect 81203 659364 81204 659428
rect 81268 659364 81269 659428
rect 81203 659363 81269 659364
rect 81206 658477 81266 659363
rect 81203 658476 81269 658477
rect 81203 658412 81204 658476
rect 81268 658412 81269 658476
rect 81203 658411 81269 658412
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 672054 131004 707102
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 387654 242604 423098
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 446443 659428 446509 659429
rect 446443 659364 446444 659428
rect 446508 659364 446509 659428
rect 446443 659363 446509 659364
rect 446446 659021 446506 659363
rect 446443 659020 446509 659021
rect 446443 658956 446444 659020
rect 446508 658956 446509 659020
rect 446443 658955 446509 658956
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 456011 659428 456077 659429
rect 456011 659364 456012 659428
rect 456076 659364 456077 659428
rect 456011 659363 456077 659364
rect 456014 658885 456074 659363
rect 456011 658884 456077 658885
rect 456011 658820 456012 658884
rect 456076 658820 456077 658884
rect 456011 658819 456077 658820
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 512683 659428 512749 659429
rect 512683 659364 512684 659428
rect 512748 659364 512749 659428
rect 512683 659363 512749 659364
rect 512686 658341 512746 659363
rect 512683 658340 512749 658341
rect 512683 658276 512684 658340
rect 512748 658276 512749 658340
rect 512683 658275 512749 658276
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use user_proj_example  mprj
timestamp 1607720773
transform 1 0 60000 0 1 60000
box 0 0 479012 600000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
