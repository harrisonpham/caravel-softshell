VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2901.310 3429.395 2901.590 3429.765 ;
        RECT 2901.380 88.245 2901.520 3429.395 ;
        RECT 2901.310 87.875 2901.590 88.245 ;
      LAYER via2 ;
        RECT 2901.310 3429.440 2901.590 3429.720 ;
        RECT 2901.310 87.920 2901.590 88.200 ;
      LAYER met3 ;
        RECT 2901.285 3429.730 2901.615 3429.745 ;
        RECT 2866.000 3429.430 2901.615 3429.730 ;
        RECT 2901.285 3429.415 2901.615 3429.430 ;
        RECT 2901.285 88.210 2901.615 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2901.285 87.910 2924.800 88.210 ;
        RECT 2901.285 87.895 2901.615 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2899.450 2435.660 2899.770 2435.720 ;
        RECT 2866.000 2435.520 2899.770 2435.660 ;
        RECT 2899.450 2435.460 2899.770 2435.520 ;
      LAYER via ;
        RECT 2899.480 2435.460 2899.740 2435.720 ;
      LAYER met2 ;
        RECT 2899.480 2435.430 2899.740 2435.750 ;
        RECT 2899.540 2434.245 2899.680 2435.430 ;
        RECT 2899.470 2433.875 2899.750 2434.245 ;
      LAYER via2 ;
        RECT 2899.470 2433.920 2899.750 2434.200 ;
      LAYER met3 ;
        RECT 2899.445 2434.210 2899.775 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2899.445 2433.910 2924.800 2434.210 ;
        RECT 2899.445 2433.895 2899.775 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2898.530 2670.260 2898.850 2670.320 ;
        RECT 2866.000 2670.120 2898.850 2670.260 ;
        RECT 2898.530 2670.060 2898.850 2670.120 ;
      LAYER via ;
        RECT 2898.560 2670.060 2898.820 2670.320 ;
      LAYER met2 ;
        RECT 2898.560 2670.030 2898.820 2670.350 ;
        RECT 2898.620 2669.525 2898.760 2670.030 ;
        RECT 2898.550 2669.155 2898.830 2669.525 ;
      LAYER via2 ;
        RECT 2898.550 2669.200 2898.830 2669.480 ;
      LAYER met3 ;
        RECT 2898.525 2669.490 2898.855 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2898.525 2669.190 2924.800 2669.490 ;
        RECT 2898.525 2669.175 2898.855 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2898.530 2904.860 2898.850 2904.920 ;
        RECT 2866.000 2904.720 2898.850 2904.860 ;
        RECT 2898.530 2904.660 2898.850 2904.720 ;
      LAYER via ;
        RECT 2898.560 2904.660 2898.820 2904.920 ;
      LAYER met2 ;
        RECT 2898.560 2904.630 2898.820 2904.950 ;
        RECT 2898.620 2904.125 2898.760 2904.630 ;
        RECT 2898.550 2903.755 2898.830 2904.125 ;
      LAYER via2 ;
        RECT 2898.550 2903.800 2898.830 2904.080 ;
      LAYER met3 ;
        RECT 2898.525 2904.090 2898.855 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2898.525 2903.790 2924.800 2904.090 ;
        RECT 2898.525 2903.775 2898.855 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2898.530 3139.460 2898.850 3139.520 ;
        RECT 2866.000 3139.320 2898.850 3139.460 ;
        RECT 2898.530 3139.260 2898.850 3139.320 ;
      LAYER via ;
        RECT 2898.560 3139.260 2898.820 3139.520 ;
      LAYER met2 ;
        RECT 2898.560 3139.230 2898.820 3139.550 ;
        RECT 2898.620 3138.725 2898.760 3139.230 ;
        RECT 2898.550 3138.355 2898.830 3138.725 ;
      LAYER via2 ;
        RECT 2898.550 3138.400 2898.830 3138.680 ;
      LAYER met3 ;
        RECT 2898.525 3138.690 2898.855 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2898.525 3138.390 2924.800 3138.690 ;
        RECT 2898.525 3138.375 2898.855 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2898.530 3374.060 2898.850 3374.120 ;
        RECT 2866.000 3373.920 2898.850 3374.060 ;
        RECT 2898.530 3373.860 2898.850 3373.920 ;
      LAYER via ;
        RECT 2898.560 3373.860 2898.820 3374.120 ;
      LAYER met2 ;
        RECT 2898.560 3373.830 2898.820 3374.150 ;
        RECT 2898.620 3373.325 2898.760 3373.830 ;
        RECT 2898.550 3372.955 2898.830 3373.325 ;
      LAYER via2 ;
        RECT 2898.550 3373.000 2898.830 3373.280 ;
      LAYER met3 ;
        RECT 2898.525 3373.290 2898.855 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2898.525 3372.990 2924.800 3373.290 ;
        RECT 2898.525 3372.975 2898.855 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3517.370 2798.480 3517.600 ;
        RECT 2798.340 3517.230 2798.940 3517.370 ;
        RECT 2798.800 3466.000 2798.940 3517.230 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3466.000 2474.640 3517.230 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3517.370 2149.420 3517.600 ;
        RECT 2149.280 3517.230 2149.880 3517.370 ;
        RECT 2149.740 3466.000 2149.880 3517.230 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3517.370 1825.120 3517.600 ;
        RECT 1824.980 3517.230 1825.580 3517.370 ;
        RECT 1825.440 3466.000 1825.580 3517.230 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3517.370 1500.820 3517.600 ;
        RECT 1500.680 3517.230 1501.280 3517.370 ;
        RECT 1501.140 3466.000 1501.280 3517.230 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2900.830 324.260 2901.150 324.320 ;
        RECT 2866.000 324.120 2901.150 324.260 ;
        RECT 2900.830 324.060 2901.150 324.120 ;
      LAYER via ;
        RECT 2900.860 324.060 2901.120 324.320 ;
      LAYER met2 ;
        RECT 2900.860 324.030 2901.120 324.350 ;
        RECT 2900.920 322.845 2901.060 324.030 ;
        RECT 2900.850 322.475 2901.130 322.845 ;
      LAYER via2 ;
        RECT 2900.850 322.520 2901.130 322.800 ;
      LAYER met3 ;
        RECT 2900.825 322.810 2901.155 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2900.825 322.510 2924.800 322.810 ;
        RECT 2900.825 322.495 2901.155 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 3466.000 1179.740 3498.270 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3498.500 851.850 3498.560 ;
        RECT 855.210 3498.500 855.530 3498.560 ;
        RECT 851.530 3498.360 855.530 3498.500 ;
        RECT 851.530 3498.300 851.850 3498.360 ;
        RECT 855.210 3498.300 855.530 3498.360 ;
      LAYER via ;
        RECT 851.560 3498.300 851.820 3498.560 ;
        RECT 855.240 3498.300 855.500 3498.560 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3498.590 851.760 3517.600 ;
        RECT 851.560 3498.270 851.820 3498.590 ;
        RECT 855.240 3498.270 855.500 3498.590 ;
        RECT 855.300 3466.000 855.440 3498.270 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.910 3498.500 531.230 3498.560 ;
        RECT 527.230 3498.360 531.230 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.910 3498.300 531.230 3498.360 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.940 3498.300 531.200 3498.560 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.940 3498.270 531.200 3498.590 ;
        RECT 531.000 3466.000 531.140 3498.270 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3502.240 202.790 3502.300 ;
        RECT 1718.170 3502.240 1718.490 3502.300 ;
        RECT 202.470 3502.100 1718.490 3502.240 ;
        RECT 202.470 3502.040 202.790 3502.100 ;
        RECT 1718.170 3502.040 1718.490 3502.100 ;
      LAYER via ;
        RECT 202.500 3502.040 202.760 3502.300 ;
        RECT 1718.200 3502.040 1718.460 3502.300 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3502.330 202.700 3517.600 ;
        RECT 202.500 3502.010 202.760 3502.330 ;
        RECT 1718.200 3502.010 1718.460 3502.330 ;
        RECT 1718.260 3466.000 1718.400 3502.010 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 27.670 3428.120 27.990 3428.180 ;
        RECT 27.670 3427.980 54.000 3428.120 ;
        RECT 27.670 3427.920 27.990 3427.980 ;
        RECT 13.870 3411.460 14.190 3411.520 ;
        RECT 27.670 3411.460 27.990 3411.520 ;
        RECT 13.870 3411.320 27.990 3411.460 ;
        RECT 13.870 3411.260 14.190 3411.320 ;
        RECT 27.670 3411.260 27.990 3411.320 ;
      LAYER via ;
        RECT 27.700 3427.920 27.960 3428.180 ;
        RECT 13.900 3411.260 14.160 3411.520 ;
        RECT 27.700 3411.260 27.960 3411.520 ;
      LAYER met2 ;
        RECT 27.700 3427.890 27.960 3428.210 ;
        RECT 27.760 3411.550 27.900 3427.890 ;
        RECT 13.900 3411.405 14.160 3411.550 ;
        RECT 13.890 3411.035 14.170 3411.405 ;
        RECT 27.700 3411.230 27.960 3411.550 ;
      LAYER via2 ;
        RECT 13.890 3411.080 14.170 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 13.865 3411.370 14.195 3411.385 ;
        RECT -4.800 3411.070 14.195 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 13.865 3411.055 14.195 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 33.650 3427.100 33.970 3427.160 ;
        RECT 33.650 3426.960 54.000 3427.100 ;
        RECT 33.650 3426.900 33.970 3426.960 ;
        RECT 13.870 3124.500 14.190 3124.560 ;
        RECT 33.650 3124.500 33.970 3124.560 ;
        RECT 13.870 3124.360 33.970 3124.500 ;
        RECT 13.870 3124.300 14.190 3124.360 ;
        RECT 33.650 3124.300 33.970 3124.360 ;
      LAYER via ;
        RECT 33.680 3426.900 33.940 3427.160 ;
        RECT 13.900 3124.300 14.160 3124.560 ;
        RECT 33.680 3124.300 33.940 3124.560 ;
      LAYER met2 ;
        RECT 33.680 3426.870 33.940 3427.190 ;
        RECT 33.740 3124.590 33.880 3426.870 ;
        RECT 13.900 3124.445 14.160 3124.590 ;
        RECT 13.890 3124.075 14.170 3124.445 ;
        RECT 33.680 3124.270 33.940 3124.590 ;
      LAYER via2 ;
        RECT 13.890 3124.120 14.170 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 13.865 3124.410 14.195 3124.425 ;
        RECT -4.800 3124.110 14.195 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 13.865 3124.095 14.195 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 33.190 3426.080 33.510 3426.140 ;
        RECT 33.190 3425.940 54.000 3426.080 ;
        RECT 33.190 3425.880 33.510 3425.940 ;
        RECT 13.870 2836.860 14.190 2836.920 ;
        RECT 33.190 2836.860 33.510 2836.920 ;
        RECT 13.870 2836.720 33.510 2836.860 ;
        RECT 13.870 2836.660 14.190 2836.720 ;
        RECT 33.190 2836.660 33.510 2836.720 ;
      LAYER via ;
        RECT 33.220 3425.880 33.480 3426.140 ;
        RECT 13.900 2836.660 14.160 2836.920 ;
        RECT 33.220 2836.660 33.480 2836.920 ;
      LAYER met2 ;
        RECT 33.220 3425.850 33.480 3426.170 ;
        RECT 33.280 2836.950 33.420 3425.850 ;
        RECT 13.900 2836.805 14.160 2836.950 ;
        RECT 13.890 2836.435 14.170 2836.805 ;
        RECT 33.220 2836.630 33.480 2836.950 ;
      LAYER via2 ;
        RECT 13.890 2836.480 14.170 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 13.865 2836.770 14.195 2836.785 ;
        RECT -4.800 2836.470 14.195 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 13.865 2836.455 14.195 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.730 3425.060 33.050 3425.120 ;
        RECT 32.730 3424.920 54.000 3425.060 ;
        RECT 32.730 3424.860 33.050 3424.920 ;
        RECT 13.870 2549.900 14.190 2549.960 ;
        RECT 32.730 2549.900 33.050 2549.960 ;
        RECT 13.870 2549.760 33.050 2549.900 ;
        RECT 13.870 2549.700 14.190 2549.760 ;
        RECT 32.730 2549.700 33.050 2549.760 ;
      LAYER via ;
        RECT 32.760 3424.860 33.020 3425.120 ;
        RECT 13.900 2549.700 14.160 2549.960 ;
        RECT 32.760 2549.700 33.020 2549.960 ;
      LAYER met2 ;
        RECT 32.760 3424.830 33.020 3425.150 ;
        RECT 32.820 2549.990 32.960 3424.830 ;
        RECT 13.900 2549.845 14.160 2549.990 ;
        RECT 13.890 2549.475 14.170 2549.845 ;
        RECT 32.760 2549.670 33.020 2549.990 ;
      LAYER via2 ;
        RECT 13.890 2549.520 14.170 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 13.865 2549.810 14.195 2549.825 ;
        RECT -4.800 2549.510 14.195 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 13.865 2549.495 14.195 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.270 3424.040 32.590 3424.100 ;
        RECT 32.270 3423.900 54.000 3424.040 ;
        RECT 32.270 3423.840 32.590 3423.900 ;
        RECT 14.330 2262.260 14.650 2262.320 ;
        RECT 32.270 2262.260 32.590 2262.320 ;
        RECT 14.330 2262.120 32.590 2262.260 ;
        RECT 14.330 2262.060 14.650 2262.120 ;
        RECT 32.270 2262.060 32.590 2262.120 ;
      LAYER via ;
        RECT 32.300 3423.840 32.560 3424.100 ;
        RECT 14.360 2262.060 14.620 2262.320 ;
        RECT 32.300 2262.060 32.560 2262.320 ;
      LAYER met2 ;
        RECT 32.300 3423.810 32.560 3424.130 ;
        RECT 32.360 2262.350 32.500 3423.810 ;
        RECT 14.360 2262.205 14.620 2262.350 ;
        RECT 14.350 2261.835 14.630 2262.205 ;
        RECT 32.300 2262.030 32.560 2262.350 ;
      LAYER via2 ;
        RECT 14.350 2261.880 14.630 2262.160 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 14.325 2262.170 14.655 2262.185 ;
        RECT -4.800 2261.870 14.655 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 14.325 2261.855 14.655 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 31.810 3423.700 32.130 3423.760 ;
        RECT 31.810 3423.560 54.000 3423.700 ;
        RECT 31.810 3423.500 32.130 3423.560 ;
        RECT 14.330 1975.300 14.650 1975.360 ;
        RECT 31.810 1975.300 32.130 1975.360 ;
        RECT 14.330 1975.160 32.130 1975.300 ;
        RECT 14.330 1975.100 14.650 1975.160 ;
        RECT 31.810 1975.100 32.130 1975.160 ;
      LAYER via ;
        RECT 31.840 3423.500 32.100 3423.760 ;
        RECT 14.360 1975.100 14.620 1975.360 ;
        RECT 31.840 1975.100 32.100 1975.360 ;
      LAYER met2 ;
        RECT 31.840 3423.470 32.100 3423.790 ;
        RECT 31.900 1975.390 32.040 3423.470 ;
        RECT 14.360 1975.245 14.620 1975.390 ;
        RECT 14.350 1974.875 14.630 1975.245 ;
        RECT 31.840 1975.070 32.100 1975.390 ;
      LAYER via2 ;
        RECT 14.350 1974.920 14.630 1975.200 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 14.325 1975.210 14.655 1975.225 ;
        RECT -4.800 1974.910 14.655 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 14.325 1974.895 14.655 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2900.830 558.860 2901.150 558.920 ;
        RECT 2866.000 558.720 2901.150 558.860 ;
        RECT 2900.830 558.660 2901.150 558.720 ;
      LAYER via ;
        RECT 2900.860 558.660 2901.120 558.920 ;
      LAYER met2 ;
        RECT 2900.860 558.630 2901.120 558.950 ;
        RECT 2900.920 557.445 2901.060 558.630 ;
        RECT 2900.850 557.075 2901.130 557.445 ;
      LAYER via2 ;
        RECT 2900.850 557.120 2901.130 557.400 ;
      LAYER met3 ;
        RECT 2900.825 557.410 2901.155 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2900.825 557.110 2924.800 557.410 ;
        RECT 2900.825 557.095 2901.155 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 31.350 3422.680 31.670 3422.740 ;
        RECT 31.350 3422.540 54.000 3422.680 ;
        RECT 31.350 3422.480 31.670 3422.540 ;
        RECT 14.790 1688.000 15.110 1688.060 ;
        RECT 31.350 1688.000 31.670 1688.060 ;
        RECT 14.790 1687.860 31.670 1688.000 ;
        RECT 14.790 1687.800 15.110 1687.860 ;
        RECT 31.350 1687.800 31.670 1687.860 ;
      LAYER via ;
        RECT 31.380 3422.480 31.640 3422.740 ;
        RECT 14.820 1687.800 15.080 1688.060 ;
        RECT 31.380 1687.800 31.640 1688.060 ;
      LAYER met2 ;
        RECT 31.380 3422.450 31.640 3422.770 ;
        RECT 31.440 1688.090 31.580 3422.450 ;
        RECT 14.820 1687.770 15.080 1688.090 ;
        RECT 31.380 1687.770 31.640 1688.090 ;
        RECT 14.880 1687.605 15.020 1687.770 ;
        RECT 14.810 1687.235 15.090 1687.605 ;
      LAYER via2 ;
        RECT 14.810 1687.280 15.090 1687.560 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 14.785 1687.570 15.115 1687.585 ;
        RECT -4.800 1687.270 15.115 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 14.785 1687.255 15.115 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.250 1476.520 15.570 1476.580 ;
        RECT 15.250 1476.380 54.000 1476.520 ;
        RECT 15.250 1476.320 15.570 1476.380 ;
      LAYER via ;
        RECT 15.280 1476.320 15.540 1476.580 ;
      LAYER met2 ;
        RECT 15.280 1476.290 15.540 1476.610 ;
        RECT 15.340 1472.045 15.480 1476.290 ;
        RECT 15.270 1471.675 15.550 1472.045 ;
      LAYER via2 ;
        RECT 15.270 1471.720 15.550 1472.000 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 15.245 1472.010 15.575 1472.025 ;
        RECT -4.800 1471.710 15.575 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 15.245 1471.695 15.575 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 1256.540 16.030 1256.600 ;
        RECT 30.890 1256.540 31.210 1256.600 ;
        RECT 15.710 1256.400 31.210 1256.540 ;
        RECT 15.710 1256.340 16.030 1256.400 ;
        RECT 30.890 1256.340 31.210 1256.400 ;
      LAYER via ;
        RECT 15.740 1256.340 16.000 1256.600 ;
        RECT 30.920 1256.340 31.180 1256.600 ;
      LAYER met2 ;
        RECT 30.910 3425.315 31.190 3425.685 ;
        RECT 30.980 1256.630 31.120 3425.315 ;
        RECT 15.740 1256.485 16.000 1256.630 ;
        RECT 15.730 1256.115 16.010 1256.485 ;
        RECT 30.920 1256.310 31.180 1256.630 ;
      LAYER via2 ;
        RECT 30.910 3425.360 31.190 3425.640 ;
        RECT 15.730 1256.160 16.010 1256.440 ;
      LAYER met3 ;
        RECT 30.885 3425.650 31.215 3425.665 ;
        RECT 30.885 3425.350 54.000 3425.650 ;
        RECT 30.885 3425.335 31.215 3425.350 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 15.705 1256.450 16.035 1256.465 ;
        RECT -4.800 1256.150 16.035 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 15.705 1256.135 16.035 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.450 3416.560 24.770 3416.620 ;
        RECT 24.450 3416.420 54.000 3416.560 ;
        RECT 24.450 3416.360 24.770 3416.420 ;
        RECT 13.870 1040.980 14.190 1041.040 ;
        RECT 24.450 1040.980 24.770 1041.040 ;
        RECT 13.870 1040.840 24.770 1040.980 ;
        RECT 13.870 1040.780 14.190 1040.840 ;
        RECT 24.450 1040.780 24.770 1040.840 ;
      LAYER via ;
        RECT 24.480 3416.360 24.740 3416.620 ;
        RECT 13.900 1040.780 14.160 1041.040 ;
        RECT 24.480 1040.780 24.740 1041.040 ;
      LAYER met2 ;
        RECT 24.480 3416.330 24.740 3416.650 ;
        RECT 24.540 1041.070 24.680 3416.330 ;
        RECT 13.900 1040.925 14.160 1041.070 ;
        RECT 13.890 1040.555 14.170 1040.925 ;
        RECT 24.480 1040.750 24.740 1041.070 ;
      LAYER via2 ;
        RECT 13.890 1040.600 14.170 1040.880 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 13.865 1040.890 14.195 1040.905 ;
        RECT -4.800 1040.590 14.195 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 13.865 1040.575 14.195 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 827.800 16.030 827.860 ;
        RECT 15.710 827.660 54.000 827.800 ;
        RECT 15.710 827.600 16.030 827.660 ;
      LAYER via ;
        RECT 15.740 827.600 16.000 827.860 ;
      LAYER met2 ;
        RECT 15.740 827.570 16.000 827.890 ;
        RECT 15.800 825.365 15.940 827.570 ;
        RECT 15.730 824.995 16.010 825.365 ;
      LAYER via2 ;
        RECT 15.730 825.040 16.010 825.320 ;
      LAYER met3 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 15.705 825.330 16.035 825.345 ;
        RECT -4.800 825.030 16.035 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 15.705 825.015 16.035 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 613.940 16.950 614.000 ;
        RECT 16.630 613.800 54.000 613.940 ;
        RECT 16.630 613.740 16.950 613.800 ;
      LAYER via ;
        RECT 16.660 613.740 16.920 614.000 ;
      LAYER met2 ;
        RECT 16.660 613.710 16.920 614.030 ;
        RECT 16.720 610.485 16.860 613.710 ;
        RECT 16.650 610.115 16.930 610.485 ;
      LAYER via2 ;
        RECT 16.650 610.160 16.930 610.440 ;
      LAYER met3 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 16.625 610.450 16.955 610.465 ;
        RECT -4.800 610.150 16.955 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 16.625 610.135 16.955 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 400.080 16.950 400.140 ;
        RECT 16.630 399.940 54.000 400.080 ;
        RECT 16.630 399.880 16.950 399.940 ;
      LAYER via ;
        RECT 16.660 399.880 16.920 400.140 ;
      LAYER met2 ;
        RECT 16.660 399.850 16.920 400.170 ;
        RECT 16.720 394.925 16.860 399.850 ;
        RECT 16.650 394.555 16.930 394.925 ;
      LAYER via2 ;
        RECT 16.650 394.600 16.930 394.880 ;
      LAYER met3 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 16.625 394.890 16.955 394.905 ;
        RECT -4.800 394.590 16.955 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 16.625 394.575 16.955 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 3430.755 17.850 3431.125 ;
        RECT 17.640 179.365 17.780 3430.755 ;
        RECT 17.570 178.995 17.850 179.365 ;
      LAYER via2 ;
        RECT 17.570 3430.800 17.850 3431.080 ;
        RECT 17.570 179.040 17.850 179.320 ;
      LAYER met3 ;
        RECT 17.545 3431.090 17.875 3431.105 ;
        RECT 17.545 3430.790 54.000 3431.090 ;
        RECT 17.545 3430.775 17.875 3430.790 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.545 179.330 17.875 179.345 ;
        RECT -4.800 179.030 17.875 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.545 179.015 17.875 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2900.830 793.460 2901.150 793.520 ;
        RECT 2866.000 793.320 2901.150 793.460 ;
        RECT 2900.830 793.260 2901.150 793.320 ;
      LAYER via ;
        RECT 2900.860 793.260 2901.120 793.520 ;
      LAYER met2 ;
        RECT 2900.860 793.230 2901.120 793.550 ;
        RECT 2900.920 792.045 2901.060 793.230 ;
        RECT 2900.850 791.675 2901.130 792.045 ;
      LAYER via2 ;
        RECT 2900.850 791.720 2901.130 792.000 ;
      LAYER met3 ;
        RECT 2900.825 792.010 2901.155 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2900.825 791.710 2924.800 792.010 ;
        RECT 2900.825 791.695 2901.155 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2887.950 3429.480 2888.270 3429.540 ;
        RECT 2866.000 3429.340 2888.270 3429.480 ;
        RECT 2887.950 3429.280 2888.270 3429.340 ;
        RECT 2887.950 1028.060 2888.270 1028.120 ;
        RECT 2903.590 1028.060 2903.910 1028.120 ;
        RECT 2887.950 1027.920 2903.910 1028.060 ;
        RECT 2887.950 1027.860 2888.270 1027.920 ;
        RECT 2903.590 1027.860 2903.910 1027.920 ;
      LAYER via ;
        RECT 2887.980 3429.280 2888.240 3429.540 ;
        RECT 2887.980 1027.860 2888.240 1028.120 ;
        RECT 2903.620 1027.860 2903.880 1028.120 ;
      LAYER met2 ;
        RECT 2887.980 3429.250 2888.240 3429.570 ;
        RECT 2888.040 1028.150 2888.180 3429.250 ;
        RECT 2887.980 1027.830 2888.240 1028.150 ;
        RECT 2903.620 1027.830 2903.880 1028.150 ;
        RECT 2903.680 1026.645 2903.820 1027.830 ;
        RECT 2903.610 1026.275 2903.890 1026.645 ;
      LAYER via2 ;
        RECT 2903.610 1026.320 2903.890 1026.600 ;
      LAYER met3 ;
        RECT 2903.585 1026.610 2903.915 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2903.585 1026.310 2924.800 1026.610 ;
        RECT 2903.585 1026.295 2903.915 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2888.410 3430.160 2888.730 3430.220 ;
        RECT 2866.000 3430.020 2888.730 3430.160 ;
        RECT 2888.410 3429.960 2888.730 3430.020 ;
        RECT 2888.410 1262.660 2888.730 1262.720 ;
        RECT 2899.910 1262.660 2900.230 1262.720 ;
        RECT 2888.410 1262.520 2900.230 1262.660 ;
        RECT 2888.410 1262.460 2888.730 1262.520 ;
        RECT 2899.910 1262.460 2900.230 1262.520 ;
      LAYER via ;
        RECT 2888.440 3429.960 2888.700 3430.220 ;
        RECT 2888.440 1262.460 2888.700 1262.720 ;
        RECT 2899.940 1262.460 2900.200 1262.720 ;
      LAYER met2 ;
        RECT 2888.440 3429.930 2888.700 3430.250 ;
        RECT 2888.500 1262.750 2888.640 3429.930 ;
        RECT 2888.440 1262.430 2888.700 1262.750 ;
        RECT 2899.940 1262.430 2900.200 1262.750 ;
        RECT 2900.000 1261.245 2900.140 1262.430 ;
        RECT 2899.930 1260.875 2900.210 1261.245 ;
      LAYER via2 ;
        RECT 2899.930 1260.920 2900.210 1261.200 ;
      LAYER met3 ;
        RECT 2899.905 1261.210 2900.235 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2899.905 1260.910 2924.800 1261.210 ;
        RECT 2899.905 1260.895 2900.235 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2900.830 1497.260 2901.150 1497.320 ;
        RECT 2866.000 1497.120 2901.150 1497.260 ;
        RECT 2900.830 1497.060 2901.150 1497.120 ;
      LAYER via ;
        RECT 2900.860 1497.060 2901.120 1497.320 ;
      LAYER met2 ;
        RECT 2900.860 1497.030 2901.120 1497.350 ;
        RECT 2900.920 1495.845 2901.060 1497.030 ;
        RECT 2900.850 1495.475 2901.130 1495.845 ;
      LAYER via2 ;
        RECT 2900.850 1495.520 2901.130 1495.800 ;
      LAYER met3 ;
        RECT 2900.825 1495.810 2901.155 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2900.825 1495.510 2924.800 1495.810 ;
        RECT 2900.825 1495.495 2901.155 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2888.870 3431.180 2889.190 3431.240 ;
        RECT 2866.000 3431.040 2889.190 3431.180 ;
        RECT 2888.870 3430.980 2889.190 3431.040 ;
        RECT 2888.870 1731.860 2889.190 1731.920 ;
        RECT 2899.450 1731.860 2899.770 1731.920 ;
        RECT 2888.870 1731.720 2899.770 1731.860 ;
        RECT 2888.870 1731.660 2889.190 1731.720 ;
        RECT 2899.450 1731.660 2899.770 1731.720 ;
      LAYER via ;
        RECT 2888.900 3430.980 2889.160 3431.240 ;
        RECT 2888.900 1731.660 2889.160 1731.920 ;
        RECT 2899.480 1731.660 2899.740 1731.920 ;
      LAYER met2 ;
        RECT 2888.900 3430.950 2889.160 3431.270 ;
        RECT 2888.960 1731.950 2889.100 3430.950 ;
        RECT 2888.900 1731.630 2889.160 1731.950 ;
        RECT 2899.480 1731.630 2899.740 1731.950 ;
        RECT 2899.540 1730.445 2899.680 1731.630 ;
        RECT 2899.470 1730.075 2899.750 1730.445 ;
      LAYER via2 ;
        RECT 2899.470 1730.120 2899.750 1730.400 ;
      LAYER met3 ;
        RECT 2899.445 1730.410 2899.775 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2899.445 1730.110 2924.800 1730.410 ;
        RECT 2899.445 1730.095 2899.775 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2899.910 1966.460 2900.230 1966.520 ;
        RECT 2866.000 1966.320 2900.230 1966.460 ;
        RECT 2899.910 1966.260 2900.230 1966.320 ;
      LAYER via ;
        RECT 2899.940 1966.260 2900.200 1966.520 ;
      LAYER met2 ;
        RECT 2899.940 1966.230 2900.200 1966.550 ;
        RECT 2900.000 1965.045 2900.140 1966.230 ;
        RECT 2899.930 1964.675 2900.210 1965.045 ;
      LAYER via2 ;
        RECT 2899.930 1964.720 2900.210 1965.000 ;
      LAYER met3 ;
        RECT 2899.905 1965.010 2900.235 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2899.905 1964.710 2924.800 1965.010 ;
        RECT 2899.905 1964.695 2900.235 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2889.330 3423.360 2889.650 3423.420 ;
        RECT 2866.000 3423.220 2889.650 3423.360 ;
        RECT 2889.330 3423.160 2889.650 3423.220 ;
        RECT 2889.330 2201.060 2889.650 2201.120 ;
        RECT 2899.450 2201.060 2899.770 2201.120 ;
        RECT 2889.330 2200.920 2899.770 2201.060 ;
        RECT 2889.330 2200.860 2889.650 2200.920 ;
        RECT 2899.450 2200.860 2899.770 2200.920 ;
      LAYER via ;
        RECT 2889.360 3423.160 2889.620 3423.420 ;
        RECT 2889.360 2200.860 2889.620 2201.120 ;
        RECT 2899.480 2200.860 2899.740 2201.120 ;
      LAYER met2 ;
        RECT 2889.360 3423.130 2889.620 3423.450 ;
        RECT 2889.420 2201.150 2889.560 3423.130 ;
        RECT 2889.360 2200.830 2889.620 2201.150 ;
        RECT 2899.480 2200.830 2899.740 2201.150 ;
        RECT 2899.540 2199.645 2899.680 2200.830 ;
        RECT 2899.470 2199.275 2899.750 2199.645 ;
      LAYER via2 ;
        RECT 2899.470 2199.320 2899.750 2199.600 ;
      LAYER met3 ;
        RECT 2899.445 2199.610 2899.775 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2899.445 2199.310 2924.800 2199.610 ;
        RECT 2899.445 2199.295 2899.775 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2887.490 206.960 2887.810 207.020 ;
        RECT 2902.670 206.960 2902.990 207.020 ;
        RECT 2887.490 206.820 2902.990 206.960 ;
        RECT 2887.490 206.760 2887.810 206.820 ;
        RECT 2902.670 206.760 2902.990 206.820 ;
      LAYER via ;
        RECT 2887.520 206.760 2887.780 207.020 ;
        RECT 2902.700 206.760 2902.960 207.020 ;
      LAYER met2 ;
        RECT 2887.510 3430.075 2887.790 3430.445 ;
        RECT 2887.580 207.050 2887.720 3430.075 ;
        RECT 2887.520 206.730 2887.780 207.050 ;
        RECT 2902.700 206.730 2902.960 207.050 ;
        RECT 2902.760 205.205 2902.900 206.730 ;
        RECT 2902.690 204.835 2902.970 205.205 ;
      LAYER via2 ;
        RECT 2887.510 3430.120 2887.790 3430.400 ;
        RECT 2902.690 204.880 2902.970 205.160 ;
      LAYER met3 ;
        RECT 2887.485 3430.410 2887.815 3430.425 ;
        RECT 2866.000 3430.110 2887.815 3430.410 ;
        RECT 2887.485 3430.095 2887.815 3430.110 ;
        RECT 2902.665 205.170 2902.995 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2902.665 204.870 2924.800 205.170 ;
        RECT 2902.665 204.855 2902.995 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2898.990 3424.380 2899.310 3424.440 ;
        RECT 2866.000 3424.240 2899.310 3424.380 ;
        RECT 2898.990 3424.180 2899.310 3424.240 ;
      LAYER via ;
        RECT 2899.020 3424.180 2899.280 3424.440 ;
      LAYER met2 ;
        RECT 2899.020 3424.150 2899.280 3424.470 ;
        RECT 2899.080 2551.885 2899.220 3424.150 ;
        RECT 2899.010 2551.515 2899.290 2551.885 ;
      LAYER via2 ;
        RECT 2899.010 2551.560 2899.290 2551.840 ;
      LAYER met3 ;
        RECT 2898.985 2551.850 2899.315 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2898.985 2551.550 2924.800 2551.850 ;
        RECT 2898.985 2551.535 2899.315 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2889.790 3425.740 2890.110 3425.800 ;
        RECT 2866.000 3425.600 2890.110 3425.740 ;
        RECT 2889.790 3425.540 2890.110 3425.600 ;
        RECT 2889.790 2786.880 2890.110 2786.940 ;
        RECT 2898.070 2786.880 2898.390 2786.940 ;
        RECT 2889.790 2786.740 2898.390 2786.880 ;
        RECT 2889.790 2786.680 2890.110 2786.740 ;
        RECT 2898.070 2786.680 2898.390 2786.740 ;
      LAYER via ;
        RECT 2889.820 3425.540 2890.080 3425.800 ;
        RECT 2889.820 2786.680 2890.080 2786.940 ;
        RECT 2898.100 2786.680 2898.360 2786.940 ;
      LAYER met2 ;
        RECT 2889.820 3425.510 2890.080 3425.830 ;
        RECT 2889.880 2786.970 2890.020 3425.510 ;
        RECT 2889.820 2786.650 2890.080 2786.970 ;
        RECT 2898.100 2786.650 2898.360 2786.970 ;
        RECT 2898.160 2786.485 2898.300 2786.650 ;
        RECT 2898.090 2786.115 2898.370 2786.485 ;
      LAYER via2 ;
        RECT 2898.090 2786.160 2898.370 2786.440 ;
      LAYER met3 ;
        RECT 2898.065 2786.450 2898.395 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2898.065 2786.150 2924.800 2786.450 ;
        RECT 2898.065 2786.135 2898.395 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2890.250 3426.420 2890.570 3426.480 ;
        RECT 2866.000 3426.280 2890.570 3426.420 ;
        RECT 2890.250 3426.220 2890.570 3426.280 ;
        RECT 2890.250 3022.160 2890.570 3022.220 ;
        RECT 2898.070 3022.160 2898.390 3022.220 ;
        RECT 2890.250 3022.020 2898.390 3022.160 ;
        RECT 2890.250 3021.960 2890.570 3022.020 ;
        RECT 2898.070 3021.960 2898.390 3022.020 ;
      LAYER via ;
        RECT 2890.280 3426.220 2890.540 3426.480 ;
        RECT 2890.280 3021.960 2890.540 3022.220 ;
        RECT 2898.100 3021.960 2898.360 3022.220 ;
      LAYER met2 ;
        RECT 2890.280 3426.190 2890.540 3426.510 ;
        RECT 2890.340 3022.250 2890.480 3426.190 ;
        RECT 2890.280 3021.930 2890.540 3022.250 ;
        RECT 2898.100 3021.930 2898.360 3022.250 ;
        RECT 2898.160 3021.085 2898.300 3021.930 ;
        RECT 2898.090 3020.715 2898.370 3021.085 ;
      LAYER via2 ;
        RECT 2898.090 3020.760 2898.370 3021.040 ;
      LAYER met3 ;
        RECT 2898.065 3021.050 2898.395 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2898.065 3020.750 2924.800 3021.050 ;
        RECT 2898.065 3020.735 2898.395 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2890.710 3427.440 2891.030 3427.500 ;
        RECT 2866.000 3427.300 2891.030 3427.440 ;
        RECT 2890.710 3427.240 2891.030 3427.300 ;
        RECT 2890.710 3256.760 2891.030 3256.820 ;
        RECT 2898.070 3256.760 2898.390 3256.820 ;
        RECT 2890.710 3256.620 2898.390 3256.760 ;
        RECT 2890.710 3256.560 2891.030 3256.620 ;
        RECT 2898.070 3256.560 2898.390 3256.620 ;
      LAYER via ;
        RECT 2890.740 3427.240 2891.000 3427.500 ;
        RECT 2890.740 3256.560 2891.000 3256.820 ;
        RECT 2898.100 3256.560 2898.360 3256.820 ;
      LAYER met2 ;
        RECT 2890.740 3427.210 2891.000 3427.530 ;
        RECT 2890.800 3256.850 2890.940 3427.210 ;
        RECT 2890.740 3256.530 2891.000 3256.850 ;
        RECT 2898.100 3256.530 2898.360 3256.850 ;
        RECT 2898.160 3255.685 2898.300 3256.530 ;
        RECT 2898.090 3255.315 2898.370 3255.685 ;
      LAYER via2 ;
        RECT 2898.090 3255.360 2898.370 3255.640 ;
      LAYER met3 ;
        RECT 2898.065 3255.650 2898.395 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2898.065 3255.350 2924.800 3255.650 ;
        RECT 2898.065 3255.335 2898.395 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1151.910 3484.900 1152.230 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 1151.910 3484.760 2901.150 3484.900 ;
        RECT 1151.910 3484.700 1152.230 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 1151.940 3484.700 1152.200 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 1151.940 3484.670 1152.200 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 1152.000 3466.000 1152.140 3484.670 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1220.910 3502.920 1221.230 3502.980 ;
        RECT 2635.870 3502.920 2636.190 3502.980 ;
        RECT 1220.910 3502.780 2636.190 3502.920 ;
        RECT 1220.910 3502.720 1221.230 3502.780 ;
        RECT 2635.870 3502.720 2636.190 3502.780 ;
      LAYER via ;
        RECT 1220.940 3502.720 1221.200 3502.980 ;
        RECT 2635.900 3502.720 2636.160 3502.980 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3503.010 2636.100 3517.600 ;
        RECT 1220.940 3502.690 1221.200 3503.010 ;
        RECT 2635.900 3502.690 2636.160 3503.010 ;
        RECT 1221.000 3466.000 1221.140 3502.690 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.010 3504.280 1283.330 3504.340 ;
        RECT 2311.570 3504.280 2311.890 3504.340 ;
        RECT 1283.010 3504.140 2311.890 3504.280 ;
        RECT 1283.010 3504.080 1283.330 3504.140 ;
        RECT 2311.570 3504.080 2311.890 3504.140 ;
      LAYER via ;
        RECT 1283.040 3504.080 1283.300 3504.340 ;
        RECT 2311.600 3504.080 2311.860 3504.340 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3504.370 2311.800 3517.600 ;
        RECT 1283.040 3504.050 1283.300 3504.370 ;
        RECT 2311.600 3504.050 2311.860 3504.370 ;
        RECT 1283.100 3466.000 1283.240 3504.050 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.010 3500.880 1352.330 3500.940 ;
        RECT 1987.270 3500.880 1987.590 3500.940 ;
        RECT 1352.010 3500.740 1987.590 3500.880 ;
        RECT 1352.010 3500.680 1352.330 3500.740 ;
        RECT 1987.270 3500.680 1987.590 3500.740 ;
      LAYER via ;
        RECT 1352.040 3500.680 1352.300 3500.940 ;
        RECT 1987.300 3500.680 1987.560 3500.940 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3500.970 1987.500 3517.600 ;
        RECT 1352.040 3500.650 1352.300 3500.970 ;
        RECT 1987.300 3500.650 1987.560 3500.970 ;
        RECT 1352.100 3466.000 1352.240 3500.650 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1421.010 3499.520 1421.330 3499.580 ;
        RECT 1662.510 3499.520 1662.830 3499.580 ;
        RECT 1421.010 3499.380 1662.830 3499.520 ;
        RECT 1421.010 3499.320 1421.330 3499.380 ;
        RECT 1662.510 3499.320 1662.830 3499.380 ;
      LAYER via ;
        RECT 1421.040 3499.320 1421.300 3499.580 ;
        RECT 1662.540 3499.320 1662.800 3499.580 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3499.610 1662.740 3517.600 ;
        RECT 1421.040 3499.290 1421.300 3499.610 ;
        RECT 1662.540 3499.290 1662.800 3499.610 ;
        RECT 1421.100 3466.000 1421.240 3499.290 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3499.180 1338.530 3499.240 ;
        RECT 1476.670 3499.180 1476.990 3499.240 ;
        RECT 1338.210 3499.040 1476.990 3499.180 ;
        RECT 1338.210 3498.980 1338.530 3499.040 ;
        RECT 1476.670 3498.980 1476.990 3499.040 ;
      LAYER via ;
        RECT 1338.240 3498.980 1338.500 3499.240 ;
        RECT 1476.700 3498.980 1476.960 3499.240 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3499.270 1338.440 3517.600 ;
        RECT 1338.240 3498.950 1338.500 3499.270 ;
        RECT 1476.700 3498.950 1476.960 3499.270 ;
        RECT 1476.760 3466.000 1476.900 3498.950 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2902.230 3430.075 2902.510 3430.445 ;
        RECT 2902.300 439.805 2902.440 3430.075 ;
        RECT 2902.230 439.435 2902.510 439.805 ;
      LAYER via2 ;
        RECT 2902.230 3430.120 2902.510 3430.400 ;
        RECT 2902.230 439.480 2902.510 439.760 ;
      LAYER met3 ;
        RECT 2866.000 3431.470 2893.090 3431.770 ;
        RECT 2892.790 3430.410 2893.090 3431.470 ;
        RECT 2902.205 3430.410 2902.535 3430.425 ;
        RECT 2892.790 3430.110 2902.535 3430.410 ;
        RECT 2902.205 3430.095 2902.535 3430.110 ;
        RECT 2902.205 439.770 2902.535 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2902.205 439.470 2924.800 439.770 ;
        RECT 2902.205 439.455 2902.535 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3500.540 1014.230 3500.600 ;
        RECT 1545.670 3500.540 1545.990 3500.600 ;
        RECT 1013.910 3500.400 1545.990 3500.540 ;
        RECT 1013.910 3500.340 1014.230 3500.400 ;
        RECT 1545.670 3500.340 1545.990 3500.400 ;
      LAYER via ;
        RECT 1013.940 3500.340 1014.200 3500.600 ;
        RECT 1545.700 3500.340 1545.960 3500.600 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3500.630 1014.140 3517.600 ;
        RECT 1013.940 3500.310 1014.200 3500.630 ;
        RECT 1545.700 3500.310 1545.960 3500.630 ;
        RECT 1545.760 3466.000 1545.900 3500.310 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3504.620 689.470 3504.680 ;
        RECT 1607.770 3504.620 1608.090 3504.680 ;
        RECT 689.150 3504.480 1608.090 3504.620 ;
        RECT 689.150 3504.420 689.470 3504.480 ;
        RECT 1607.770 3504.420 1608.090 3504.480 ;
      LAYER via ;
        RECT 689.180 3504.420 689.440 3504.680 ;
        RECT 1607.800 3504.420 1608.060 3504.680 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3504.710 689.380 3517.600 ;
        RECT 689.180 3504.390 689.440 3504.710 ;
        RECT 1607.800 3504.390 1608.060 3504.710 ;
        RECT 1607.860 3466.000 1608.000 3504.390 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 3503.260 365.170 3503.320 ;
        RECT 1676.770 3503.260 1677.090 3503.320 ;
        RECT 364.850 3503.120 1677.090 3503.260 ;
        RECT 364.850 3503.060 365.170 3503.120 ;
        RECT 1676.770 3503.060 1677.090 3503.120 ;
      LAYER via ;
        RECT 364.880 3503.060 365.140 3503.320 ;
        RECT 1676.800 3503.060 1677.060 3503.320 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3503.350 365.080 3517.600 ;
        RECT 364.880 3503.030 365.140 3503.350 ;
        RECT 1676.800 3503.030 1677.060 3503.350 ;
        RECT 1676.860 3466.000 1677.000 3503.030 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.550 3501.560 40.870 3501.620 ;
        RECT 1738.870 3501.560 1739.190 3501.620 ;
        RECT 40.550 3501.420 1739.190 3501.560 ;
        RECT 40.550 3501.360 40.870 3501.420 ;
        RECT 1738.870 3501.360 1739.190 3501.420 ;
      LAYER via ;
        RECT 40.580 3501.360 40.840 3501.620 ;
        RECT 1738.900 3501.360 1739.160 3501.620 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.650 40.780 3517.600 ;
        RECT 40.580 3501.330 40.840 3501.650 ;
        RECT 1738.900 3501.330 1739.160 3501.650 ;
        RECT 1738.960 3466.000 1739.100 3501.330 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 3270.360 14.190 3270.420 ;
        RECT 13.870 3270.220 54.000 3270.360 ;
        RECT 13.870 3270.160 14.190 3270.220 ;
      LAYER via ;
        RECT 13.900 3270.160 14.160 3270.420 ;
      LAYER met2 ;
        RECT 13.900 3270.130 14.160 3270.450 ;
        RECT 13.960 3267.925 14.100 3270.130 ;
        RECT 13.890 3267.555 14.170 3267.925 ;
      LAYER via2 ;
        RECT 13.890 3267.600 14.170 3267.880 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 13.865 3267.890 14.195 3267.905 ;
        RECT -4.800 3267.590 14.195 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 13.865 3267.575 14.195 3267.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 2980.680 14.190 2980.740 ;
        RECT 13.870 2980.540 54.000 2980.680 ;
        RECT 13.870 2980.480 14.190 2980.540 ;
      LAYER via ;
        RECT 13.900 2980.480 14.160 2980.740 ;
      LAYER met2 ;
        RECT 13.900 2980.450 14.160 2980.770 ;
        RECT 13.960 2980.285 14.100 2980.450 ;
        RECT 13.890 2979.915 14.170 2980.285 ;
      LAYER via2 ;
        RECT 13.890 2979.960 14.170 2980.240 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 13.865 2980.250 14.195 2980.265 ;
        RECT -4.800 2979.950 14.195 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 13.865 2979.935 14.195 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 2697.800 14.190 2697.860 ;
        RECT 13.870 2697.660 54.000 2697.800 ;
        RECT 13.870 2697.600 14.190 2697.660 ;
      LAYER via ;
        RECT 13.900 2697.600 14.160 2697.860 ;
      LAYER met2 ;
        RECT 13.900 2697.570 14.160 2697.890 ;
        RECT 13.960 2693.325 14.100 2697.570 ;
        RECT 13.890 2692.955 14.170 2693.325 ;
      LAYER via2 ;
        RECT 13.890 2693.000 14.170 2693.280 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 13.865 2693.290 14.195 2693.305 ;
        RECT -4.800 2692.990 14.195 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 13.865 2692.975 14.195 2692.990 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 2408.120 14.650 2408.180 ;
        RECT 14.330 2407.980 54.000 2408.120 ;
        RECT 14.330 2407.920 14.650 2407.980 ;
      LAYER via ;
        RECT 14.360 2407.920 14.620 2408.180 ;
      LAYER met2 ;
        RECT 14.360 2407.890 14.620 2408.210 ;
        RECT 14.420 2405.685 14.560 2407.890 ;
        RECT 14.350 2405.315 14.630 2405.685 ;
      LAYER via2 ;
        RECT 14.350 2405.360 14.630 2405.640 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 14.325 2405.650 14.655 2405.665 ;
        RECT -4.800 2405.350 14.655 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 14.325 2405.335 14.655 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 2125.240 14.650 2125.300 ;
        RECT 14.330 2125.100 54.000 2125.240 ;
        RECT 14.330 2125.040 14.650 2125.100 ;
      LAYER via ;
        RECT 14.360 2125.040 14.620 2125.300 ;
      LAYER met2 ;
        RECT 14.360 2125.010 14.620 2125.330 ;
        RECT 14.420 2118.725 14.560 2125.010 ;
        RECT 14.350 2118.355 14.630 2118.725 ;
      LAYER via2 ;
        RECT 14.350 2118.400 14.630 2118.680 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 14.325 2118.690 14.655 2118.705 ;
        RECT -4.800 2118.390 14.655 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 14.325 2118.375 14.655 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 1835.220 15.110 1835.280 ;
        RECT 14.790 1835.080 54.000 1835.220 ;
        RECT 14.790 1835.020 15.110 1835.080 ;
      LAYER via ;
        RECT 14.820 1835.020 15.080 1835.280 ;
      LAYER met2 ;
        RECT 14.820 1834.990 15.080 1835.310 ;
        RECT 14.880 1831.085 15.020 1834.990 ;
        RECT 14.810 1830.715 15.090 1831.085 ;
      LAYER via2 ;
        RECT 14.810 1830.760 15.090 1831.040 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 14.785 1831.050 15.115 1831.065 ;
        RECT -4.800 1830.750 15.115 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 14.785 1830.735 15.115 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2904.070 3432.115 2904.350 3432.485 ;
        RECT 2904.140 674.405 2904.280 3432.115 ;
        RECT 2904.070 674.035 2904.350 674.405 ;
      LAYER via2 ;
        RECT 2904.070 3432.160 2904.350 3432.440 ;
        RECT 2904.070 674.080 2904.350 674.360 ;
      LAYER met3 ;
        RECT 2904.045 3432.450 2904.375 3432.465 ;
        RECT 2866.000 3432.150 2904.375 3432.450 ;
        RECT 2904.045 3432.135 2904.375 3432.150 ;
        RECT 2904.045 674.370 2904.375 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2904.045 674.070 2924.800 674.370 ;
        RECT 2904.045 674.055 2904.375 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3431.520 15.570 3431.580 ;
        RECT 15.250 3431.380 54.000 3431.520 ;
        RECT 15.250 3431.320 15.570 3431.380 ;
      LAYER via ;
        RECT 15.280 3431.320 15.540 3431.580 ;
      LAYER met2 ;
        RECT 15.280 3431.290 15.540 3431.610 ;
        RECT 15.340 1544.125 15.480 3431.290 ;
        RECT 15.270 1543.755 15.550 1544.125 ;
      LAYER via2 ;
        RECT 15.270 1543.800 15.550 1544.080 ;
      LAYER met3 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 15.245 1544.090 15.575 1544.105 ;
        RECT -4.800 1543.790 15.575 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 15.245 1543.775 15.575 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 3430.840 16.490 3430.900 ;
        RECT 16.170 3430.700 54.000 3430.840 ;
        RECT 16.170 3430.640 16.490 3430.700 ;
      LAYER via ;
        RECT 16.200 3430.640 16.460 3430.900 ;
      LAYER met2 ;
        RECT 16.200 3430.610 16.460 3430.930 ;
        RECT 16.260 1328.565 16.400 3430.610 ;
        RECT 16.190 1328.195 16.470 1328.565 ;
      LAYER via2 ;
        RECT 16.190 1328.240 16.470 1328.520 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 16.165 1328.530 16.495 1328.545 ;
        RECT -4.800 1328.230 16.495 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 16.165 1328.215 16.495 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 1117.820 16.950 1117.880 ;
        RECT 16.630 1117.680 54.000 1117.820 ;
        RECT 16.630 1117.620 16.950 1117.680 ;
      LAYER via ;
        RECT 16.660 1117.620 16.920 1117.880 ;
      LAYER met2 ;
        RECT 16.660 1117.590 16.920 1117.910 ;
        RECT 16.720 1113.005 16.860 1117.590 ;
        RECT 16.650 1112.635 16.930 1113.005 ;
      LAYER via2 ;
        RECT 16.650 1112.680 16.930 1112.960 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 16.625 1112.970 16.955 1112.985 ;
        RECT -4.800 1112.670 16.955 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 16.625 1112.655 16.955 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 897.500 14.190 897.560 ;
        RECT 23.990 897.500 24.310 897.560 ;
        RECT 13.870 897.360 24.310 897.500 ;
        RECT 13.870 897.300 14.190 897.360 ;
        RECT 23.990 897.300 24.310 897.360 ;
      LAYER via ;
        RECT 13.900 897.300 14.160 897.560 ;
        RECT 24.020 897.300 24.280 897.560 ;
      LAYER met2 ;
        RECT 24.010 3435.515 24.290 3435.885 ;
        RECT 24.080 897.590 24.220 3435.515 ;
        RECT 13.900 897.445 14.160 897.590 ;
        RECT 13.890 897.075 14.170 897.445 ;
        RECT 24.020 897.270 24.280 897.590 ;
      LAYER via2 ;
        RECT 24.010 3435.560 24.290 3435.840 ;
        RECT 13.890 897.120 14.170 897.400 ;
      LAYER met3 ;
        RECT 23.985 3435.850 24.315 3435.865 ;
        RECT 23.985 3435.550 54.000 3435.850 ;
        RECT 23.985 3435.535 24.315 3435.550 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 13.865 897.410 14.195 897.425 ;
        RECT -4.800 897.110 14.195 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 13.865 897.095 14.195 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 682.960 16.950 683.020 ;
        RECT 16.630 682.820 54.000 682.960 ;
        RECT 16.630 682.760 16.950 682.820 ;
      LAYER via ;
        RECT 16.660 682.760 16.920 683.020 ;
      LAYER met2 ;
        RECT 16.660 682.730 16.920 683.050 ;
        RECT 16.720 681.885 16.860 682.730 ;
        RECT 16.650 681.515 16.930 681.885 ;
      LAYER via2 ;
        RECT 16.650 681.560 16.930 681.840 ;
      LAYER met3 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 16.625 681.850 16.955 681.865 ;
        RECT -4.800 681.550 16.955 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 16.625 681.535 16.955 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.490 3434.155 18.770 3434.525 ;
        RECT 18.560 466.325 18.700 3434.155 ;
        RECT 18.490 465.955 18.770 466.325 ;
      LAYER via2 ;
        RECT 18.490 3434.200 18.770 3434.480 ;
        RECT 18.490 466.000 18.770 466.280 ;
      LAYER met3 ;
        RECT 18.465 3434.490 18.795 3434.505 ;
        RECT 18.465 3434.190 54.000 3434.490 ;
        RECT 18.465 3434.175 18.795 3434.190 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 18.465 466.290 18.795 466.305 ;
        RECT -4.800 465.990 18.795 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 18.465 465.975 18.795 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.030 3417.155 18.310 3417.525 ;
        RECT 18.100 250.765 18.240 3417.155 ;
        RECT 18.030 250.395 18.310 250.765 ;
      LAYER via2 ;
        RECT 18.030 3417.200 18.310 3417.480 ;
        RECT 18.030 250.440 18.310 250.720 ;
      LAYER met3 ;
        RECT 18.005 3417.490 18.335 3417.505 ;
        RECT 18.005 3417.190 54.000 3417.490 ;
        RECT 18.005 3417.175 18.335 3417.190 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 18.005 250.730 18.335 250.745 ;
        RECT -4.800 250.430 18.335 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 18.005 250.415 18.335 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.110 3418.515 17.390 3418.885 ;
        RECT 34.130 3418.515 34.410 3418.885 ;
        RECT 17.180 35.885 17.320 3418.515 ;
        RECT 34.200 3416.165 34.340 3418.515 ;
        RECT 34.130 3415.795 34.410 3416.165 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 17.110 3418.560 17.390 3418.840 ;
        RECT 34.130 3418.560 34.410 3418.840 ;
        RECT 34.130 3415.840 34.410 3416.120 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 17.085 3418.850 17.415 3418.865 ;
        RECT 34.105 3418.850 34.435 3418.865 ;
        RECT 17.085 3418.550 34.435 3418.850 ;
        RECT 17.085 3418.535 17.415 3418.550 ;
        RECT 34.105 3418.535 34.435 3418.550 ;
        RECT 34.105 3416.130 34.435 3416.145 ;
        RECT 34.105 3415.830 54.000 3416.130 ;
        RECT 34.105 3415.815 34.435 3415.830 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2900.390 3434.835 2900.670 3435.205 ;
        RECT 2900.460 909.685 2900.600 3434.835 ;
        RECT 2900.390 909.315 2900.670 909.685 ;
      LAYER via2 ;
        RECT 2900.390 3434.880 2900.670 3435.160 ;
        RECT 2900.390 909.360 2900.670 909.640 ;
      LAYER met3 ;
        RECT 2900.365 3435.170 2900.695 3435.185 ;
        RECT 2866.000 3434.870 2900.695 3435.170 ;
        RECT 2900.365 3434.855 2900.695 3434.870 ;
        RECT 2900.365 909.650 2900.695 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.365 909.350 2924.800 909.650 ;
        RECT 2900.365 909.335 2900.695 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2903.590 3416.220 2903.910 3416.280 ;
        RECT 2866.000 3416.080 2903.910 3416.220 ;
        RECT 2903.590 3416.020 2903.910 3416.080 ;
      LAYER via ;
        RECT 2903.620 3416.020 2903.880 3416.280 ;
      LAYER met2 ;
        RECT 2903.620 3415.990 2903.880 3416.310 ;
        RECT 2903.680 1144.285 2903.820 3415.990 ;
        RECT 2903.610 1143.915 2903.890 1144.285 ;
      LAYER via2 ;
        RECT 2903.610 1143.960 2903.890 1144.240 ;
      LAYER met3 ;
        RECT 2903.585 1144.250 2903.915 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2903.585 1143.950 2924.800 1144.250 ;
        RECT 2903.585 1143.935 2903.915 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2904.510 3421.660 2904.830 3421.720 ;
        RECT 2866.000 3421.520 2904.830 3421.660 ;
        RECT 2904.510 3421.460 2904.830 3421.520 ;
      LAYER via ;
        RECT 2904.540 3421.460 2904.800 3421.720 ;
      LAYER met2 ;
        RECT 2904.540 3421.430 2904.800 3421.750 ;
        RECT 2904.600 1378.885 2904.740 3421.430 ;
        RECT 2904.530 1378.515 2904.810 1378.885 ;
      LAYER via2 ;
        RECT 2904.530 1378.560 2904.810 1378.840 ;
      LAYER met3 ;
        RECT 2904.505 1378.850 2904.835 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2904.505 1378.550 2924.800 1378.850 ;
        RECT 2904.505 1378.535 2904.835 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 3419.280 2901.150 3419.340 ;
        RECT 2866.000 3419.140 2901.150 3419.280 ;
        RECT 2900.830 3419.080 2901.150 3419.140 ;
      LAYER via ;
        RECT 2900.860 3419.080 2901.120 3419.340 ;
      LAYER met2 ;
        RECT 2900.860 3419.050 2901.120 3419.370 ;
        RECT 2900.920 1613.485 2901.060 3419.050 ;
        RECT 2900.850 1613.115 2901.130 1613.485 ;
      LAYER via2 ;
        RECT 2900.850 1613.160 2901.130 1613.440 ;
      LAYER met3 ;
        RECT 2900.825 1613.450 2901.155 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.825 1613.150 2924.800 1613.450 ;
        RECT 2900.825 1613.135 2901.155 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2899.910 1849.160 2900.230 1849.220 ;
        RECT 2866.000 1849.020 2900.230 1849.160 ;
        RECT 2899.910 1848.960 2900.230 1849.020 ;
      LAYER via ;
        RECT 2899.940 1848.960 2900.200 1849.220 ;
      LAYER met2 ;
        RECT 2899.940 1848.930 2900.200 1849.250 ;
        RECT 2900.000 1848.085 2900.140 1848.930 ;
        RECT 2899.930 1847.715 2900.210 1848.085 ;
      LAYER via2 ;
        RECT 2899.930 1847.760 2900.210 1848.040 ;
      LAYER met3 ;
        RECT 2899.905 1848.050 2900.235 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2899.905 1847.750 2924.800 1848.050 ;
        RECT 2899.905 1847.735 2900.235 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2899.910 3426.080 2900.230 3426.140 ;
        RECT 2866.000 3425.940 2900.230 3426.080 ;
        RECT 2899.910 3425.880 2900.230 3425.940 ;
      LAYER via ;
        RECT 2899.940 3425.880 2900.200 3426.140 ;
      LAYER met2 ;
        RECT 2899.940 3425.850 2900.200 3426.170 ;
        RECT 2900.000 2082.685 2900.140 3425.850 ;
        RECT 2899.930 2082.315 2900.210 2082.685 ;
      LAYER via2 ;
        RECT 2899.930 2082.360 2900.210 2082.640 ;
      LAYER met3 ;
        RECT 2899.905 2082.650 2900.235 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2899.905 2082.350 2924.800 2082.650 ;
        RECT 2899.905 2082.335 2900.235 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2899.450 2318.360 2899.770 2318.420 ;
        RECT 2866.000 2318.220 2899.770 2318.360 ;
        RECT 2899.450 2318.160 2899.770 2318.220 ;
      LAYER via ;
        RECT 2899.480 2318.160 2899.740 2318.420 ;
      LAYER met2 ;
        RECT 2899.480 2318.130 2899.740 2318.450 ;
        RECT 2899.540 2317.285 2899.680 2318.130 ;
        RECT 2899.470 2316.915 2899.750 2317.285 ;
      LAYER via2 ;
        RECT 2899.470 2316.960 2899.750 2317.240 ;
      LAYER met3 ;
        RECT 2899.445 2317.250 2899.775 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2899.445 2316.950 2924.800 2317.250 ;
        RECT 2899.445 2316.935 2899.775 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2899.450 151.540 2899.770 151.600 ;
        RECT 2866.000 151.400 2899.770 151.540 ;
        RECT 2899.450 151.340 2899.770 151.400 ;
      LAYER via ;
        RECT 2899.480 151.340 2899.740 151.600 ;
      LAYER met2 ;
        RECT 2899.480 151.310 2899.740 151.630 ;
        RECT 2899.540 146.725 2899.680 151.310 ;
        RECT 2899.470 146.355 2899.750 146.725 ;
      LAYER via2 ;
        RECT 2899.470 146.400 2899.750 146.680 ;
      LAYER met3 ;
        RECT 2899.445 146.690 2899.775 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2899.445 146.390 2924.800 146.690 ;
        RECT 2899.445 146.375 2899.775 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2899.450 3418.260 2899.770 3418.320 ;
        RECT 2866.000 3418.120 2899.770 3418.260 ;
        RECT 2899.450 3418.060 2899.770 3418.120 ;
      LAYER via ;
        RECT 2899.480 3418.060 2899.740 3418.320 ;
      LAYER met2 ;
        RECT 2899.480 3418.030 2899.740 3418.350 ;
        RECT 2899.540 2493.405 2899.680 3418.030 ;
        RECT 2899.470 2493.035 2899.750 2493.405 ;
      LAYER via2 ;
        RECT 2899.470 2493.080 2899.750 2493.360 ;
      LAYER met3 ;
        RECT 2899.445 2493.370 2899.775 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2899.445 2493.070 2924.800 2493.370 ;
        RECT 2899.445 2493.055 2899.775 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2898.530 2732.140 2898.850 2732.200 ;
        RECT 2866.000 2732.000 2898.850 2732.140 ;
        RECT 2898.530 2731.940 2898.850 2732.000 ;
      LAYER via ;
        RECT 2898.560 2731.940 2898.820 2732.200 ;
      LAYER met2 ;
        RECT 2898.560 2731.910 2898.820 2732.230 ;
        RECT 2898.620 2728.005 2898.760 2731.910 ;
        RECT 2898.550 2727.635 2898.830 2728.005 ;
      LAYER via2 ;
        RECT 2898.550 2727.680 2898.830 2727.960 ;
      LAYER met3 ;
        RECT 2898.525 2727.970 2898.855 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2898.525 2727.670 2924.800 2727.970 ;
        RECT 2898.525 2727.655 2898.855 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2898.530 2966.740 2898.850 2966.800 ;
        RECT 2866.000 2966.600 2898.850 2966.740 ;
        RECT 2898.530 2966.540 2898.850 2966.600 ;
      LAYER via ;
        RECT 2898.560 2966.540 2898.820 2966.800 ;
      LAYER met2 ;
        RECT 2898.560 2966.510 2898.820 2966.830 ;
        RECT 2898.620 2962.605 2898.760 2966.510 ;
        RECT 2898.550 2962.235 2898.830 2962.605 ;
      LAYER via2 ;
        RECT 2898.550 2962.280 2898.830 2962.560 ;
      LAYER met3 ;
        RECT 2898.525 2962.570 2898.855 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2898.525 2962.270 2924.800 2962.570 ;
        RECT 2898.525 2962.255 2898.855 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2898.530 3201.340 2898.850 3201.400 ;
        RECT 2866.000 3201.200 2898.850 3201.340 ;
        RECT 2898.530 3201.140 2898.850 3201.200 ;
      LAYER via ;
        RECT 2898.560 3201.140 2898.820 3201.400 ;
      LAYER met2 ;
        RECT 2898.560 3201.110 2898.820 3201.430 ;
        RECT 2898.620 3197.205 2898.760 3201.110 ;
        RECT 2898.550 3196.835 2898.830 3197.205 ;
      LAYER via2 ;
        RECT 2898.550 3196.880 2898.830 3197.160 ;
      LAYER met3 ;
        RECT 2898.525 3197.170 2898.855 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2898.525 3196.870 2924.800 3197.170 ;
        RECT 2898.525 3196.855 2898.855 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 3434.920 2901.150 3434.980 ;
        RECT 2866.000 3434.780 2901.150 3434.920 ;
        RECT 2900.830 3434.720 2901.150 3434.780 ;
      LAYER via ;
        RECT 2900.860 3434.720 2901.120 3434.980 ;
      LAYER met2 ;
        RECT 2900.860 3434.690 2901.120 3435.010 ;
        RECT 2900.920 3431.805 2901.060 3434.690 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1241.610 3502.580 1241.930 3502.640 ;
        RECT 2717.290 3502.580 2717.610 3502.640 ;
        RECT 1241.610 3502.440 2717.610 3502.580 ;
        RECT 1241.610 3502.380 1241.930 3502.440 ;
        RECT 2717.290 3502.380 2717.610 3502.440 ;
      LAYER via ;
        RECT 1241.640 3502.380 1241.900 3502.640 ;
        RECT 2717.320 3502.380 2717.580 3502.640 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3502.670 2717.520 3517.600 ;
        RECT 1241.640 3502.350 1241.900 3502.670 ;
        RECT 2717.320 3502.350 2717.580 3502.670 ;
        RECT 1241.700 3466.000 1241.840 3502.350 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1310.610 3503.940 1310.930 3504.000 ;
        RECT 2392.530 3503.940 2392.850 3504.000 ;
        RECT 1310.610 3503.800 2392.850 3503.940 ;
        RECT 1310.610 3503.740 1310.930 3503.800 ;
        RECT 2392.530 3503.740 2392.850 3503.800 ;
      LAYER via ;
        RECT 1310.640 3503.740 1310.900 3504.000 ;
        RECT 2392.560 3503.740 2392.820 3504.000 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3504.030 2392.760 3517.600 ;
        RECT 1310.640 3503.710 1310.900 3504.030 ;
        RECT 2392.560 3503.710 2392.820 3504.030 ;
        RECT 1310.700 3466.000 1310.840 3503.710 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1372.710 3501.220 1373.030 3501.280 ;
        RECT 2068.230 3501.220 2068.550 3501.280 ;
        RECT 1372.710 3501.080 2068.550 3501.220 ;
        RECT 1372.710 3501.020 1373.030 3501.080 ;
        RECT 2068.230 3501.020 2068.550 3501.080 ;
      LAYER via ;
        RECT 1372.740 3501.020 1373.000 3501.280 ;
        RECT 2068.260 3501.020 2068.520 3501.280 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3501.310 2068.460 3517.600 ;
        RECT 1372.740 3500.990 1373.000 3501.310 ;
        RECT 2068.260 3500.990 2068.520 3501.310 ;
        RECT 1372.800 3466.000 1372.940 3500.990 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1441.710 3499.860 1442.030 3499.920 ;
        RECT 1743.930 3499.860 1744.250 3499.920 ;
        RECT 1441.710 3499.720 1744.250 3499.860 ;
        RECT 1441.710 3499.660 1442.030 3499.720 ;
        RECT 1743.930 3499.660 1744.250 3499.720 ;
      LAYER via ;
        RECT 1441.740 3499.660 1442.000 3499.920 ;
        RECT 1743.960 3499.660 1744.220 3499.920 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3499.950 1744.160 3517.600 ;
        RECT 1441.740 3499.630 1442.000 3499.950 ;
        RECT 1743.960 3499.630 1744.220 3499.950 ;
        RECT 1441.800 3466.000 1441.940 3499.630 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.170 3498.840 1419.490 3498.900 ;
        RECT 1497.370 3498.840 1497.690 3498.900 ;
        RECT 1419.170 3498.700 1497.690 3498.840 ;
        RECT 1419.170 3498.640 1419.490 3498.700 ;
        RECT 1497.370 3498.640 1497.690 3498.700 ;
      LAYER via ;
        RECT 1419.200 3498.640 1419.460 3498.900 ;
        RECT 1497.400 3498.640 1497.660 3498.900 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3498.930 1419.400 3517.600 ;
        RECT 1419.200 3498.610 1419.460 3498.930 ;
        RECT 1497.400 3498.610 1497.660 3498.930 ;
        RECT 1497.460 3466.000 1497.600 3498.610 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2901.770 3427.355 2902.050 3427.725 ;
        RECT 2901.840 381.325 2901.980 3427.355 ;
        RECT 2901.770 380.955 2902.050 381.325 ;
      LAYER via2 ;
        RECT 2901.770 3427.400 2902.050 3427.680 ;
        RECT 2901.770 381.000 2902.050 381.280 ;
      LAYER met3 ;
        RECT 2901.745 3427.690 2902.075 3427.705 ;
        RECT 2866.000 3427.390 2902.075 3427.690 ;
        RECT 2901.745 3427.375 2902.075 3427.390 ;
        RECT 2901.745 381.290 2902.075 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2901.745 380.990 2924.800 381.290 ;
        RECT 2901.745 380.975 2902.075 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1094.870 3500.200 1095.190 3500.260 ;
        RECT 1566.370 3500.200 1566.690 3500.260 ;
        RECT 1094.870 3500.060 1566.690 3500.200 ;
        RECT 1094.870 3500.000 1095.190 3500.060 ;
        RECT 1566.370 3500.000 1566.690 3500.060 ;
      LAYER via ;
        RECT 1094.900 3500.000 1095.160 3500.260 ;
        RECT 1566.400 3500.000 1566.660 3500.260 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3500.290 1095.100 3517.600 ;
        RECT 1094.900 3499.970 1095.160 3500.290 ;
        RECT 1566.400 3499.970 1566.660 3500.290 ;
        RECT 1566.460 3466.000 1566.600 3499.970 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 770.570 3504.960 770.890 3505.020 ;
        RECT 1628.470 3504.960 1628.790 3505.020 ;
        RECT 770.570 3504.820 1628.790 3504.960 ;
        RECT 770.570 3504.760 770.890 3504.820 ;
        RECT 1628.470 3504.760 1628.790 3504.820 ;
      LAYER via ;
        RECT 770.600 3504.760 770.860 3505.020 ;
        RECT 1628.500 3504.760 1628.760 3505.020 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3505.050 770.800 3517.600 ;
        RECT 770.600 3504.730 770.860 3505.050 ;
        RECT 1628.500 3504.730 1628.760 3505.050 ;
        RECT 1628.560 3466.000 1628.700 3504.730 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3503.600 446.130 3503.660 ;
        RECT 1697.470 3503.600 1697.790 3503.660 ;
        RECT 445.810 3503.460 1697.790 3503.600 ;
        RECT 445.810 3503.400 446.130 3503.460 ;
        RECT 1697.470 3503.400 1697.790 3503.460 ;
      LAYER via ;
        RECT 445.840 3503.400 446.100 3503.660 ;
        RECT 1697.500 3503.400 1697.760 3503.660 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3503.690 446.040 3517.600 ;
        RECT 445.840 3503.370 446.100 3503.690 ;
        RECT 1697.500 3503.370 1697.760 3503.690 ;
        RECT 1697.560 3466.000 1697.700 3503.370 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3501.900 121.830 3501.960 ;
        RECT 1759.570 3501.900 1759.890 3501.960 ;
        RECT 121.510 3501.760 1759.890 3501.900 ;
        RECT 121.510 3501.700 121.830 3501.760 ;
        RECT 1759.570 3501.700 1759.890 3501.760 ;
      LAYER via ;
        RECT 121.540 3501.700 121.800 3501.960 ;
        RECT 1759.600 3501.700 1759.860 3501.960 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3501.990 121.740 3517.600 ;
        RECT 121.540 3501.670 121.800 3501.990 ;
        RECT 1759.600 3501.670 1759.860 3501.990 ;
        RECT 1759.660 3466.000 1759.800 3501.670 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 3346.520 14.190 3346.580 ;
        RECT 13.870 3346.380 54.000 3346.520 ;
        RECT 13.870 3346.320 14.190 3346.380 ;
      LAYER via ;
        RECT 13.900 3346.320 14.160 3346.580 ;
      LAYER met2 ;
        RECT 13.900 3346.290 14.160 3346.610 ;
        RECT 13.960 3340.005 14.100 3346.290 ;
        RECT 13.890 3339.635 14.170 3340.005 ;
      LAYER via2 ;
        RECT 13.890 3339.680 14.170 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 13.865 3339.970 14.195 3339.985 ;
        RECT -4.800 3339.670 14.195 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 13.865 3339.655 14.195 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 25.370 3419.280 25.690 3419.340 ;
        RECT 25.370 3419.140 54.000 3419.280 ;
        RECT 25.370 3419.080 25.690 3419.140 ;
        RECT 13.870 3052.420 14.190 3052.480 ;
        RECT 25.370 3052.420 25.690 3052.480 ;
        RECT 13.870 3052.280 25.690 3052.420 ;
        RECT 13.870 3052.220 14.190 3052.280 ;
        RECT 25.370 3052.220 25.690 3052.280 ;
      LAYER via ;
        RECT 25.400 3419.080 25.660 3419.340 ;
        RECT 13.900 3052.220 14.160 3052.480 ;
        RECT 25.400 3052.220 25.660 3052.480 ;
      LAYER met2 ;
        RECT 25.400 3419.050 25.660 3419.370 ;
        RECT 25.460 3052.510 25.600 3419.050 ;
        RECT 13.900 3052.365 14.160 3052.510 ;
        RECT 13.890 3051.995 14.170 3052.365 ;
        RECT 25.400 3052.190 25.660 3052.510 ;
      LAYER via2 ;
        RECT 13.890 3052.040 14.170 3052.320 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 13.865 3052.330 14.195 3052.345 ;
        RECT -4.800 3052.030 14.195 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 13.865 3052.015 14.195 3052.030 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 2766.820 14.190 2766.880 ;
        RECT 13.870 2766.680 54.000 2766.820 ;
        RECT 13.870 2766.620 14.190 2766.680 ;
      LAYER via ;
        RECT 13.900 2766.620 14.160 2766.880 ;
      LAYER met2 ;
        RECT 13.900 2766.590 14.160 2766.910 ;
        RECT 13.960 2765.405 14.100 2766.590 ;
        RECT 13.890 2765.035 14.170 2765.405 ;
      LAYER via2 ;
        RECT 13.890 2765.080 14.170 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 13.865 2765.370 14.195 2765.385 ;
        RECT -4.800 2765.070 14.195 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 13.865 2765.055 14.195 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 3433.560 14.650 3433.620 ;
        RECT 14.330 3433.420 54.000 3433.560 ;
        RECT 14.330 3433.360 14.650 3433.420 ;
      LAYER via ;
        RECT 14.360 3433.360 14.620 3433.620 ;
      LAYER met2 ;
        RECT 14.360 3433.330 14.620 3433.650 ;
        RECT 14.420 2477.765 14.560 3433.330 ;
        RECT 14.350 2477.395 14.630 2477.765 ;
      LAYER via2 ;
        RECT 14.350 2477.440 14.630 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 14.325 2477.730 14.655 2477.745 ;
        RECT -4.800 2477.430 14.655 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 14.325 2477.415 14.655 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 24.910 3432.880 25.230 3432.940 ;
        RECT 24.910 3432.740 54.000 3432.880 ;
        RECT 24.910 3432.680 25.230 3432.740 ;
        RECT 13.870 2193.580 14.190 2193.640 ;
        RECT 24.910 2193.580 25.230 2193.640 ;
        RECT 13.870 2193.440 25.230 2193.580 ;
        RECT 13.870 2193.380 14.190 2193.440 ;
        RECT 24.910 2193.380 25.230 2193.440 ;
      LAYER via ;
        RECT 24.940 3432.680 25.200 3432.940 ;
        RECT 13.900 2193.380 14.160 2193.640 ;
        RECT 24.940 2193.380 25.200 2193.640 ;
      LAYER met2 ;
        RECT 24.940 3432.650 25.200 3432.970 ;
        RECT 25.000 2193.670 25.140 3432.650 ;
        RECT 13.900 2193.350 14.160 2193.670 ;
        RECT 24.940 2193.350 25.200 2193.670 ;
        RECT 13.960 2190.125 14.100 2193.350 ;
        RECT 13.890 2189.755 14.170 2190.125 ;
      LAYER via2 ;
        RECT 13.890 2189.800 14.170 2190.080 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 13.865 2190.090 14.195 2190.105 ;
        RECT -4.800 2189.790 14.195 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 13.865 2189.775 14.195 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 3417.580 15.110 3417.640 ;
        RECT 14.790 3417.440 54.000 3417.580 ;
        RECT 14.790 3417.380 15.110 3417.440 ;
      LAYER via ;
        RECT 14.820 3417.380 15.080 3417.640 ;
      LAYER met2 ;
        RECT 14.820 3417.350 15.080 3417.670 ;
        RECT 14.880 1903.165 15.020 3417.350 ;
        RECT 14.810 1902.795 15.090 1903.165 ;
      LAYER via2 ;
        RECT 14.810 1902.840 15.090 1903.120 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 14.785 1903.130 15.115 1903.145 ;
        RECT -4.800 1902.830 15.115 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 14.785 1902.815 15.115 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2903.150 3433.475 2903.430 3433.845 ;
        RECT 2903.220 615.925 2903.360 3433.475 ;
        RECT 2903.150 615.555 2903.430 615.925 ;
      LAYER via2 ;
        RECT 2903.150 3433.520 2903.430 3433.800 ;
        RECT 2903.150 615.600 2903.430 615.880 ;
      LAYER met3 ;
        RECT 2903.125 3433.810 2903.455 3433.825 ;
        RECT 2866.000 3433.510 2903.455 3433.810 ;
        RECT 2903.125 3433.495 2903.455 3433.510 ;
        RECT 2903.125 615.890 2903.455 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2903.125 615.590 2924.800 615.890 ;
        RECT 2903.125 615.575 2903.455 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 37.790 3431.860 38.110 3431.920 ;
        RECT 37.790 3431.720 54.000 3431.860 ;
        RECT 37.790 3431.660 38.110 3431.720 ;
        RECT 14.790 1615.580 15.110 1615.640 ;
        RECT 37.790 1615.580 38.110 1615.640 ;
        RECT 14.790 1615.440 38.110 1615.580 ;
        RECT 14.790 1615.380 15.110 1615.440 ;
        RECT 37.790 1615.380 38.110 1615.440 ;
      LAYER via ;
        RECT 37.820 3431.660 38.080 3431.920 ;
        RECT 14.820 1615.380 15.080 1615.640 ;
        RECT 37.820 1615.380 38.080 1615.640 ;
      LAYER met2 ;
        RECT 37.820 3431.630 38.080 3431.950 ;
        RECT 37.880 1615.670 38.020 3431.630 ;
        RECT 14.820 1615.525 15.080 1615.670 ;
        RECT 14.810 1615.155 15.090 1615.525 ;
        RECT 37.820 1615.350 38.080 1615.670 ;
      LAYER via2 ;
        RECT 14.810 1615.200 15.090 1615.480 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 14.785 1615.490 15.115 1615.505 ;
        RECT -4.800 1615.190 15.115 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 14.785 1615.175 15.115 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 3416.900 16.030 3416.960 ;
        RECT 15.710 3416.760 54.000 3416.900 ;
        RECT 15.710 3416.700 16.030 3416.760 ;
      LAYER via ;
        RECT 15.740 3416.700 16.000 3416.960 ;
      LAYER met2 ;
        RECT 15.740 3416.670 16.000 3416.990 ;
        RECT 15.800 1400.645 15.940 3416.670 ;
        RECT 15.730 1400.275 16.010 1400.645 ;
      LAYER via2 ;
        RECT 15.730 1400.320 16.010 1400.600 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 15.705 1400.610 16.035 1400.625 ;
        RECT -4.800 1400.310 16.035 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 15.705 1400.295 16.035 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 3430.500 16.950 3430.560 ;
        RECT 16.630 3430.360 54.000 3430.500 ;
        RECT 16.630 3430.300 16.950 3430.360 ;
      LAYER via ;
        RECT 16.660 3430.300 16.920 3430.560 ;
      LAYER met2 ;
        RECT 16.660 3430.270 16.920 3430.590 ;
        RECT 16.720 1185.085 16.860 3430.270 ;
        RECT 16.650 1184.715 16.930 1185.085 ;
      LAYER via2 ;
        RECT 16.650 1184.760 16.930 1185.040 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 16.625 1185.050 16.955 1185.065 ;
        RECT -4.800 1184.750 16.955 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 16.625 1184.735 16.955 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 3429.820 20.630 3429.880 ;
        RECT 20.310 3429.680 54.000 3429.820 ;
        RECT 20.310 3429.620 20.630 3429.680 ;
      LAYER via ;
        RECT 20.340 3429.620 20.600 3429.880 ;
      LAYER met2 ;
        RECT 20.340 3429.590 20.600 3429.910 ;
        RECT 20.400 969.525 20.540 3429.590 ;
        RECT 20.330 969.155 20.610 969.525 ;
      LAYER via2 ;
        RECT 20.330 969.200 20.610 969.480 ;
      LAYER met3 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 20.305 969.490 20.635 969.505 ;
        RECT -4.800 969.190 20.635 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 20.305 969.175 20.635 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.870 3417.835 20.150 3418.205 ;
        RECT 19.940 753.965 20.080 3417.835 ;
        RECT 19.870 753.595 20.150 753.965 ;
      LAYER via2 ;
        RECT 19.870 3417.880 20.150 3418.160 ;
        RECT 19.870 753.640 20.150 753.920 ;
      LAYER met3 ;
        RECT 19.845 3418.170 20.175 3418.185 ;
        RECT 19.845 3417.870 54.000 3418.170 ;
        RECT 19.845 3417.855 20.175 3417.870 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 19.845 753.930 20.175 753.945 ;
        RECT -4.800 753.630 20.175 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 19.845 753.615 20.175 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.410 3432.795 19.690 3433.165 ;
        RECT 19.480 538.405 19.620 3432.795 ;
        RECT 19.410 538.035 19.690 538.405 ;
      LAYER via2 ;
        RECT 19.410 3432.840 19.690 3433.120 ;
        RECT 19.410 538.080 19.690 538.360 ;
      LAYER met3 ;
        RECT 19.385 3433.130 19.715 3433.145 ;
        RECT 19.385 3432.830 54.000 3433.130 ;
        RECT 19.385 3432.815 19.715 3432.830 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 19.385 538.370 19.715 538.385 ;
        RECT -4.800 538.070 19.715 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 19.385 538.055 19.715 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.950 3416.475 19.230 3416.845 ;
        RECT 19.020 322.845 19.160 3416.475 ;
        RECT 18.950 322.475 19.230 322.845 ;
      LAYER via2 ;
        RECT 18.950 3416.520 19.230 3416.800 ;
        RECT 18.950 322.520 19.230 322.800 ;
      LAYER met3 ;
        RECT 18.925 3416.810 19.255 3416.825 ;
        RECT 18.925 3416.510 54.000 3416.810 ;
        RECT 18.925 3416.495 19.255 3416.510 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 18.925 322.810 19.255 322.825 ;
        RECT -4.800 322.510 19.255 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 18.925 322.495 19.255 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 110.400 17.870 110.460 ;
        RECT 17.550 110.260 54.000 110.400 ;
        RECT 17.550 110.200 17.870 110.260 ;
      LAYER via ;
        RECT 17.580 110.200 17.840 110.460 ;
      LAYER met2 ;
        RECT 17.580 110.170 17.840 110.490 ;
        RECT 17.640 107.285 17.780 110.170 ;
        RECT 17.570 106.915 17.850 107.285 ;
      LAYER via2 ;
        RECT 17.570 106.960 17.850 107.240 ;
      LAYER met3 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 17.545 107.250 17.875 107.265 ;
        RECT -4.800 106.950 17.875 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 17.545 106.935 17.875 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2902.670 3415.880 2902.990 3415.940 ;
        RECT 2866.000 3415.740 2902.990 3415.880 ;
        RECT 2902.670 3415.680 2902.990 3415.740 ;
      LAYER via ;
        RECT 2902.700 3415.680 2902.960 3415.940 ;
      LAYER met2 ;
        RECT 2902.700 3415.650 2902.960 3415.970 ;
        RECT 2902.760 850.525 2902.900 3415.650 ;
        RECT 2902.690 850.155 2902.970 850.525 ;
      LAYER via2 ;
        RECT 2902.690 850.200 2902.970 850.480 ;
      LAYER met3 ;
        RECT 2902.665 850.490 2902.995 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2902.665 850.190 2924.800 850.490 ;
        RECT 2902.665 850.175 2902.995 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 2866.000 1089.800 2901.150 1089.940 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 1324.540 2901.150 1324.600 ;
        RECT 2866.000 1324.400 2901.150 1324.540 ;
        RECT 2900.830 1324.340 2901.150 1324.400 ;
      LAYER via ;
        RECT 2900.860 1324.340 2901.120 1324.600 ;
      LAYER met2 ;
        RECT 2900.860 1324.310 2901.120 1324.630 ;
        RECT 2900.920 1319.725 2901.060 1324.310 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 1559.140 2901.150 1559.200 ;
        RECT 2866.000 1559.000 2901.150 1559.140 ;
        RECT 2900.830 1558.940 2901.150 1559.000 ;
      LAYER via ;
        RECT 2900.860 1558.940 2901.120 1559.200 ;
      LAYER met2 ;
        RECT 2900.860 1558.910 2901.120 1559.230 ;
        RECT 2900.920 1554.325 2901.060 1558.910 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
      LAYER via2 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
      LAYER met3 ;
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2899.910 1793.740 2900.230 1793.800 ;
        RECT 2866.000 1793.600 2900.230 1793.740 ;
        RECT 2899.910 1793.540 2900.230 1793.600 ;
      LAYER via ;
        RECT 2899.940 1793.540 2900.200 1793.800 ;
      LAYER met2 ;
        RECT 2899.940 1793.510 2900.200 1793.830 ;
        RECT 2900.000 1789.605 2900.140 1793.510 ;
        RECT 2899.930 1789.235 2900.210 1789.605 ;
      LAYER via2 ;
        RECT 2899.930 1789.280 2900.210 1789.560 ;
      LAYER met3 ;
        RECT 2899.905 1789.570 2900.235 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2899.905 1789.270 2924.800 1789.570 ;
        RECT 2899.905 1789.255 2900.235 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2899.910 2028.340 2900.230 2028.400 ;
        RECT 2866.000 2028.200 2900.230 2028.340 ;
        RECT 2899.910 2028.140 2900.230 2028.200 ;
      LAYER via ;
        RECT 2899.940 2028.140 2900.200 2028.400 ;
      LAYER met2 ;
        RECT 2899.940 2028.110 2900.200 2028.430 ;
        RECT 2900.000 2024.205 2900.140 2028.110 ;
        RECT 2899.930 2023.835 2900.210 2024.205 ;
      LAYER via2 ;
        RECT 2899.930 2023.880 2900.210 2024.160 ;
      LAYER met3 ;
        RECT 2899.905 2024.170 2900.235 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2899.905 2023.870 2924.800 2024.170 ;
        RECT 2899.905 2023.855 2900.235 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2899.450 2262.940 2899.770 2263.000 ;
        RECT 2866.000 2262.800 2899.770 2262.940 ;
        RECT 2899.450 2262.740 2899.770 2262.800 ;
      LAYER via ;
        RECT 2899.480 2262.740 2899.740 2263.000 ;
      LAYER met2 ;
        RECT 2899.480 2262.710 2899.740 2263.030 ;
        RECT 2899.540 2258.805 2899.680 2262.710 ;
        RECT 2899.470 2258.435 2899.750 2258.805 ;
      LAYER via2 ;
        RECT 2899.470 2258.480 2899.750 2258.760 ;
      LAYER met3 ;
        RECT 2899.445 2258.770 2899.775 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2899.445 2258.470 2924.800 2258.770 ;
        RECT 2899.445 2258.455 2899.775 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 633.030 18.260 633.350 18.320 ;
        RECT 738.370 18.260 738.690 18.320 ;
        RECT 633.030 18.120 738.690 18.260 ;
        RECT 633.030 18.060 633.350 18.120 ;
        RECT 738.370 18.060 738.690 18.120 ;
      LAYER via ;
        RECT 633.060 18.060 633.320 18.320 ;
        RECT 738.400 18.060 738.660 18.320 ;
      LAYER met2 ;
        RECT 738.460 18.350 738.600 54.000 ;
        RECT 633.060 18.030 633.320 18.350 ;
        RECT 738.400 18.030 738.660 18.350 ;
        RECT 633.120 2.400 633.260 18.030 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2415.160 3.130 2415.300 54.000 ;
        RECT 2415.160 2.990 2417.600 3.130 ;
        RECT 2417.460 2.400 2417.600 2.990 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2429.330 2.960 2429.650 3.020 ;
        RECT 2434.850 2.960 2435.170 3.020 ;
        RECT 2429.330 2.820 2435.170 2.960 ;
        RECT 2429.330 2.760 2429.650 2.820 ;
        RECT 2434.850 2.760 2435.170 2.820 ;
      LAYER via ;
        RECT 2429.360 2.760 2429.620 3.020 ;
        RECT 2434.880 2.760 2435.140 3.020 ;
      LAYER met2 ;
        RECT 2429.420 3.050 2429.560 54.000 ;
        RECT 2429.360 2.730 2429.620 3.050 ;
        RECT 2434.880 2.730 2435.140 3.050 ;
        RECT 2434.940 2.400 2435.080 2.730 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2449.570 2.960 2449.890 3.020 ;
        RECT 2452.790 2.960 2453.110 3.020 ;
        RECT 2449.570 2.820 2453.110 2.960 ;
        RECT 2449.570 2.760 2449.890 2.820 ;
        RECT 2452.790 2.760 2453.110 2.820 ;
      LAYER via ;
        RECT 2449.600 2.760 2449.860 3.020 ;
        RECT 2452.820 2.760 2453.080 3.020 ;
      LAYER met2 ;
        RECT 2449.660 3.050 2449.800 54.000 ;
        RECT 2449.600 2.730 2449.860 3.050 ;
        RECT 2452.820 2.730 2453.080 3.050 ;
        RECT 2452.880 2.400 2453.020 2.730 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2471.280 3.130 2471.420 54.000 ;
        RECT 2470.820 2.990 2471.420 3.130 ;
        RECT 2470.820 2.400 2470.960 2.990 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2484.070 2.960 2484.390 3.020 ;
        RECT 2488.670 2.960 2488.990 3.020 ;
        RECT 2484.070 2.820 2488.990 2.960 ;
        RECT 2484.070 2.760 2484.390 2.820 ;
        RECT 2488.670 2.760 2488.990 2.820 ;
      LAYER via ;
        RECT 2484.100 2.760 2484.360 3.020 ;
        RECT 2488.700 2.760 2488.960 3.020 ;
      LAYER met2 ;
        RECT 2484.160 3.050 2484.300 54.000 ;
        RECT 2484.100 2.730 2484.360 3.050 ;
        RECT 2488.700 2.730 2488.960 3.050 ;
        RECT 2488.760 2.400 2488.900 2.730 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2352.510 25.060 2352.830 25.120 ;
        RECT 2506.150 25.060 2506.470 25.120 ;
        RECT 2352.510 24.920 2506.470 25.060 ;
        RECT 2352.510 24.860 2352.830 24.920 ;
        RECT 2506.150 24.860 2506.470 24.920 ;
      LAYER via ;
        RECT 2352.540 24.860 2352.800 25.120 ;
        RECT 2506.180 24.860 2506.440 25.120 ;
      LAYER met2 ;
        RECT 2352.600 25.150 2352.740 54.000 ;
        RECT 2352.540 24.830 2352.800 25.150 ;
        RECT 2506.180 24.830 2506.440 25.150 ;
        RECT 2506.240 2.400 2506.380 24.830 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2366.310 26.420 2366.630 26.480 ;
        RECT 2524.090 26.420 2524.410 26.480 ;
        RECT 2366.310 26.280 2524.410 26.420 ;
        RECT 2366.310 26.220 2366.630 26.280 ;
        RECT 2524.090 26.220 2524.410 26.280 ;
      LAYER via ;
        RECT 2366.340 26.220 2366.600 26.480 ;
        RECT 2524.120 26.220 2524.380 26.480 ;
      LAYER met2 ;
        RECT 2366.400 26.510 2366.540 54.000 ;
        RECT 2366.340 26.190 2366.600 26.510 ;
        RECT 2524.120 26.190 2524.380 26.510 ;
        RECT 2524.180 2.400 2524.320 26.190 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2380.110 25.740 2380.430 25.800 ;
        RECT 2542.030 25.740 2542.350 25.800 ;
        RECT 2380.110 25.600 2542.350 25.740 ;
        RECT 2380.110 25.540 2380.430 25.600 ;
        RECT 2542.030 25.540 2542.350 25.600 ;
      LAYER via ;
        RECT 2380.140 25.540 2380.400 25.800 ;
        RECT 2542.060 25.540 2542.320 25.800 ;
      LAYER met2 ;
        RECT 2380.200 25.830 2380.340 54.000 ;
        RECT 2380.140 25.510 2380.400 25.830 ;
        RECT 2542.060 25.510 2542.320 25.830 ;
        RECT 2542.120 2.400 2542.260 25.510 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2393.910 26.080 2394.230 26.140 ;
        RECT 2559.970 26.080 2560.290 26.140 ;
        RECT 2393.910 25.940 2560.290 26.080 ;
        RECT 2393.910 25.880 2394.230 25.940 ;
        RECT 2559.970 25.880 2560.290 25.940 ;
      LAYER via ;
        RECT 2393.940 25.880 2394.200 26.140 ;
        RECT 2560.000 25.880 2560.260 26.140 ;
      LAYER met2 ;
        RECT 2394.000 26.170 2394.140 54.000 ;
        RECT 2393.940 25.850 2394.200 26.170 ;
        RECT 2560.000 25.850 2560.260 26.170 ;
        RECT 2560.060 2.400 2560.200 25.850 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2414.150 26.760 2414.470 26.820 ;
        RECT 2577.910 26.760 2578.230 26.820 ;
        RECT 2414.150 26.620 2578.230 26.760 ;
        RECT 2414.150 26.560 2414.470 26.620 ;
        RECT 2577.910 26.560 2578.230 26.620 ;
      LAYER via ;
        RECT 2414.180 26.560 2414.440 26.820 ;
        RECT 2577.940 26.560 2578.200 26.820 ;
      LAYER met2 ;
        RECT 2414.240 26.850 2414.380 54.000 ;
        RECT 2414.180 26.530 2414.440 26.850 ;
        RECT 2577.940 26.530 2578.200 26.850 ;
        RECT 2578.000 2.400 2578.140 26.530 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 811.510 17.580 811.830 17.640 ;
        RECT 813.810 17.580 814.130 17.640 ;
        RECT 811.510 17.440 814.130 17.580 ;
        RECT 811.510 17.380 811.830 17.440 ;
        RECT 813.810 17.380 814.130 17.440 ;
      LAYER via ;
        RECT 811.540 17.380 811.800 17.640 ;
        RECT 813.840 17.380 814.100 17.640 ;
      LAYER met2 ;
        RECT 813.900 17.670 814.040 54.000 ;
        RECT 811.540 17.350 811.800 17.670 ;
        RECT 813.840 17.350 814.100 17.670 ;
        RECT 811.600 2.400 811.740 17.350 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2428.410 24.720 2428.730 24.780 ;
        RECT 2595.390 24.720 2595.710 24.780 ;
        RECT 2428.410 24.580 2595.710 24.720 ;
        RECT 2428.410 24.520 2428.730 24.580 ;
        RECT 2595.390 24.520 2595.710 24.580 ;
      LAYER via ;
        RECT 2428.440 24.520 2428.700 24.780 ;
        RECT 2595.420 24.520 2595.680 24.780 ;
      LAYER met2 ;
        RECT 2428.500 24.810 2428.640 54.000 ;
        RECT 2428.440 24.490 2428.700 24.810 ;
        RECT 2595.420 24.490 2595.680 24.810 ;
        RECT 2595.480 2.400 2595.620 24.490 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2442.210 24.380 2442.530 24.440 ;
        RECT 2613.330 24.380 2613.650 24.440 ;
        RECT 2442.210 24.240 2613.650 24.380 ;
        RECT 2442.210 24.180 2442.530 24.240 ;
        RECT 2613.330 24.180 2613.650 24.240 ;
      LAYER via ;
        RECT 2442.240 24.180 2442.500 24.440 ;
        RECT 2613.360 24.180 2613.620 24.440 ;
      LAYER met2 ;
        RECT 2442.300 24.470 2442.440 54.000 ;
        RECT 2442.240 24.150 2442.500 24.470 ;
        RECT 2613.360 24.150 2613.620 24.470 ;
        RECT 2613.420 2.400 2613.560 24.150 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2628.970 2.960 2629.290 3.020 ;
        RECT 2631.270 2.960 2631.590 3.020 ;
        RECT 2628.970 2.820 2631.590 2.960 ;
        RECT 2628.970 2.760 2629.290 2.820 ;
        RECT 2631.270 2.760 2631.590 2.820 ;
      LAYER via ;
        RECT 2629.000 2.760 2629.260 3.020 ;
        RECT 2631.300 2.760 2631.560 3.020 ;
      LAYER met2 ;
        RECT 2629.060 3.050 2629.200 54.000 ;
        RECT 2629.000 2.730 2629.260 3.050 ;
        RECT 2631.300 2.730 2631.560 3.050 ;
        RECT 2631.360 2.400 2631.500 2.730 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2476.250 24.040 2476.570 24.100 ;
        RECT 2649.210 24.040 2649.530 24.100 ;
        RECT 2476.250 23.900 2649.530 24.040 ;
        RECT 2476.250 23.840 2476.570 23.900 ;
        RECT 2649.210 23.840 2649.530 23.900 ;
      LAYER via ;
        RECT 2476.280 23.840 2476.540 24.100 ;
        RECT 2649.240 23.840 2649.500 24.100 ;
      LAYER met2 ;
        RECT 2476.340 24.130 2476.480 54.000 ;
        RECT 2476.280 23.810 2476.540 24.130 ;
        RECT 2649.240 23.810 2649.500 24.130 ;
        RECT 2649.300 2.400 2649.440 23.810 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2507.990 27.440 2508.310 27.500 ;
        RECT 2667.150 27.440 2667.470 27.500 ;
        RECT 2507.990 27.300 2667.470 27.440 ;
        RECT 2507.990 27.240 2508.310 27.300 ;
        RECT 2667.150 27.240 2667.470 27.300 ;
      LAYER via ;
        RECT 2508.020 27.240 2508.280 27.500 ;
        RECT 2667.180 27.240 2667.440 27.500 ;
      LAYER met2 ;
        RECT 2508.080 27.530 2508.220 54.000 ;
        RECT 2508.020 27.210 2508.280 27.530 ;
        RECT 2667.180 27.210 2667.440 27.530 ;
        RECT 2667.240 2.400 2667.380 27.210 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2504.310 25.400 2504.630 25.460 ;
        RECT 2684.630 25.400 2684.950 25.460 ;
        RECT 2504.310 25.260 2684.950 25.400 ;
        RECT 2504.310 25.200 2504.630 25.260 ;
        RECT 2684.630 25.200 2684.950 25.260 ;
      LAYER via ;
        RECT 2504.340 25.200 2504.600 25.460 ;
        RECT 2684.660 25.200 2684.920 25.460 ;
      LAYER met2 ;
        RECT 2504.400 25.490 2504.540 54.000 ;
        RECT 2504.340 25.170 2504.600 25.490 ;
        RECT 2684.660 25.170 2684.920 25.490 ;
        RECT 2684.720 2.400 2684.860 25.170 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2528.690 26.420 2529.010 26.480 ;
        RECT 2702.570 26.420 2702.890 26.480 ;
        RECT 2528.690 26.280 2702.890 26.420 ;
        RECT 2528.690 26.220 2529.010 26.280 ;
        RECT 2702.570 26.220 2702.890 26.280 ;
      LAYER via ;
        RECT 2528.720 26.220 2528.980 26.480 ;
        RECT 2702.600 26.220 2702.860 26.480 ;
      LAYER met2 ;
        RECT 2528.780 26.510 2528.920 54.000 ;
        RECT 2528.720 26.190 2528.980 26.510 ;
        RECT 2702.600 26.190 2702.860 26.510 ;
        RECT 2702.660 2.400 2702.800 26.190 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2535.590 25.060 2535.910 25.120 ;
        RECT 2720.510 25.060 2720.830 25.120 ;
        RECT 2535.590 24.920 2720.830 25.060 ;
        RECT 2535.590 24.860 2535.910 24.920 ;
        RECT 2720.510 24.860 2720.830 24.920 ;
      LAYER via ;
        RECT 2535.620 24.860 2535.880 25.120 ;
        RECT 2720.540 24.860 2720.800 25.120 ;
      LAYER met2 ;
        RECT 2535.680 25.150 2535.820 54.000 ;
        RECT 2535.620 24.830 2535.880 25.150 ;
        RECT 2720.540 24.830 2720.800 25.150 ;
        RECT 2720.600 2.400 2720.740 24.830 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2556.290 25.740 2556.610 25.800 ;
        RECT 2738.450 25.740 2738.770 25.800 ;
        RECT 2556.290 25.600 2738.770 25.740 ;
        RECT 2556.290 25.540 2556.610 25.600 ;
        RECT 2738.450 25.540 2738.770 25.600 ;
      LAYER via ;
        RECT 2556.320 25.540 2556.580 25.800 ;
        RECT 2738.480 25.540 2738.740 25.800 ;
      LAYER met2 ;
        RECT 2556.380 25.830 2556.520 54.000 ;
        RECT 2556.320 25.510 2556.580 25.830 ;
        RECT 2738.480 25.510 2738.740 25.830 ;
        RECT 2738.540 2.400 2738.680 25.510 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2576.990 26.080 2577.310 26.140 ;
        RECT 2755.930 26.080 2756.250 26.140 ;
        RECT 2576.990 25.940 2756.250 26.080 ;
        RECT 2576.990 25.880 2577.310 25.940 ;
        RECT 2755.930 25.880 2756.250 25.940 ;
      LAYER via ;
        RECT 2577.020 25.880 2577.280 26.140 ;
        RECT 2755.960 25.880 2756.220 26.140 ;
      LAYER met2 ;
        RECT 2577.080 26.170 2577.220 54.000 ;
        RECT 2577.020 25.850 2577.280 26.170 ;
        RECT 2755.960 25.850 2756.220 26.170 ;
        RECT 2756.020 2.400 2756.160 25.850 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 829.450 17.580 829.770 17.640 ;
        RECT 834.510 17.580 834.830 17.640 ;
        RECT 829.450 17.440 834.830 17.580 ;
        RECT 829.450 17.380 829.770 17.440 ;
        RECT 834.510 17.380 834.830 17.440 ;
      LAYER via ;
        RECT 829.480 17.380 829.740 17.640 ;
        RECT 834.540 17.380 834.800 17.640 ;
      LAYER met2 ;
        RECT 834.600 17.670 834.740 54.000 ;
        RECT 829.480 17.350 829.740 17.670 ;
        RECT 834.540 17.350 834.800 17.670 ;
        RECT 829.540 2.400 829.680 17.350 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2611.490 26.760 2611.810 26.820 ;
        RECT 2773.870 26.760 2774.190 26.820 ;
        RECT 2611.490 26.620 2774.190 26.760 ;
        RECT 2611.490 26.560 2611.810 26.620 ;
        RECT 2773.870 26.560 2774.190 26.620 ;
      LAYER via ;
        RECT 2611.520 26.560 2611.780 26.820 ;
        RECT 2773.900 26.560 2774.160 26.820 ;
      LAYER met2 ;
        RECT 2611.580 26.850 2611.720 54.000 ;
        RECT 2611.520 26.530 2611.780 26.850 ;
        RECT 2773.900 26.530 2774.160 26.850 ;
        RECT 2773.960 2.400 2774.100 26.530 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2593.550 31.180 2593.870 31.240 ;
        RECT 2791.810 31.180 2792.130 31.240 ;
        RECT 2593.550 31.040 2792.130 31.180 ;
        RECT 2593.550 30.980 2593.870 31.040 ;
        RECT 2791.810 30.980 2792.130 31.040 ;
      LAYER via ;
        RECT 2593.580 30.980 2593.840 31.240 ;
        RECT 2791.840 30.980 2792.100 31.240 ;
      LAYER met2 ;
        RECT 2593.640 31.270 2593.780 54.000 ;
        RECT 2593.580 30.950 2593.840 31.270 ;
        RECT 2791.840 30.950 2792.100 31.270 ;
        RECT 2791.900 2.400 2792.040 30.950 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2614.250 24.380 2614.570 24.440 ;
        RECT 2809.750 24.380 2810.070 24.440 ;
        RECT 2614.250 24.240 2810.070 24.380 ;
        RECT 2614.250 24.180 2614.570 24.240 ;
        RECT 2809.750 24.180 2810.070 24.240 ;
      LAYER via ;
        RECT 2614.280 24.180 2614.540 24.440 ;
        RECT 2809.780 24.180 2810.040 24.440 ;
      LAYER met2 ;
        RECT 2614.340 24.470 2614.480 54.000 ;
        RECT 2614.280 24.150 2614.540 24.470 ;
        RECT 2809.780 24.150 2810.040 24.470 ;
        RECT 2809.840 2.400 2809.980 24.150 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2659.790 27.100 2660.110 27.160 ;
        RECT 2827.690 27.100 2828.010 27.160 ;
        RECT 2659.790 26.960 2828.010 27.100 ;
        RECT 2659.790 26.900 2660.110 26.960 ;
        RECT 2827.690 26.900 2828.010 26.960 ;
      LAYER via ;
        RECT 2659.820 26.900 2660.080 27.160 ;
        RECT 2827.720 26.900 2827.980 27.160 ;
      LAYER met2 ;
        RECT 2659.880 27.190 2660.020 54.000 ;
        RECT 2659.820 26.870 2660.080 27.190 ;
        RECT 2827.720 26.870 2827.980 27.190 ;
        RECT 2827.780 2.400 2827.920 26.870 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2642.310 30.840 2642.630 30.900 ;
        RECT 2845.170 30.840 2845.490 30.900 ;
        RECT 2642.310 30.700 2845.490 30.840 ;
        RECT 2642.310 30.640 2642.630 30.700 ;
        RECT 2845.170 30.640 2845.490 30.700 ;
      LAYER via ;
        RECT 2642.340 30.640 2642.600 30.900 ;
        RECT 2845.200 30.640 2845.460 30.900 ;
      LAYER met2 ;
        RECT 2642.400 30.930 2642.540 54.000 ;
        RECT 2642.340 30.610 2642.600 30.930 ;
        RECT 2845.200 30.610 2845.460 30.930 ;
        RECT 2845.260 2.400 2845.400 30.610 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2666.690 24.720 2667.010 24.780 ;
        RECT 2863.110 24.720 2863.430 24.780 ;
        RECT 2666.690 24.580 2863.430 24.720 ;
        RECT 2666.690 24.520 2667.010 24.580 ;
        RECT 2863.110 24.520 2863.430 24.580 ;
      LAYER via ;
        RECT 2666.720 24.520 2666.980 24.780 ;
        RECT 2863.140 24.520 2863.400 24.780 ;
      LAYER met2 ;
        RECT 2666.780 24.810 2666.920 54.000 ;
        RECT 2666.720 24.490 2666.980 24.810 ;
        RECT 2863.140 24.490 2863.400 24.810 ;
        RECT 2863.200 2.400 2863.340 24.490 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2680.490 24.040 2680.810 24.100 ;
        RECT 2881.050 24.040 2881.370 24.100 ;
        RECT 2680.490 23.900 2881.370 24.040 ;
        RECT 2680.490 23.840 2680.810 23.900 ;
        RECT 2881.050 23.840 2881.370 23.900 ;
      LAYER via ;
        RECT 2680.520 23.840 2680.780 24.100 ;
        RECT 2881.080 23.840 2881.340 24.100 ;
      LAYER met2 ;
        RECT 2680.580 24.130 2680.720 54.000 ;
        RECT 2680.520 23.810 2680.780 24.130 ;
        RECT 2881.080 23.810 2881.340 24.130 ;
        RECT 2881.140 2.400 2881.280 23.810 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2839.190 18.260 2839.510 18.320 ;
        RECT 2898.990 18.260 2899.310 18.320 ;
        RECT 2839.190 18.120 2899.310 18.260 ;
        RECT 2839.190 18.060 2839.510 18.120 ;
        RECT 2898.990 18.060 2899.310 18.120 ;
      LAYER via ;
        RECT 2839.220 18.060 2839.480 18.320 ;
        RECT 2899.020 18.060 2899.280 18.320 ;
      LAYER met2 ;
        RECT 2839.280 18.350 2839.420 54.000 ;
        RECT 2839.220 18.030 2839.480 18.350 ;
        RECT 2899.020 18.030 2899.280 18.350 ;
        RECT 2899.080 2.400 2899.220 18.030 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 848.400 17.410 848.540 54.000 ;
        RECT 847.020 17.270 848.540 17.410 ;
        RECT 847.020 2.400 847.160 17.270 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 864.870 17.580 865.190 17.640 ;
        RECT 869.010 17.580 869.330 17.640 ;
        RECT 864.870 17.440 869.330 17.580 ;
        RECT 864.870 17.380 865.190 17.440 ;
        RECT 869.010 17.380 869.330 17.440 ;
      LAYER via ;
        RECT 864.900 17.380 865.160 17.640 ;
        RECT 869.040 17.380 869.300 17.640 ;
      LAYER met2 ;
        RECT 869.100 17.670 869.240 54.000 ;
        RECT 864.900 17.350 865.160 17.670 ;
        RECT 869.040 17.350 869.300 17.670 ;
        RECT 864.960 2.400 865.100 17.350 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.900 2.400 883.040 54.000 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 900.750 17.580 901.070 17.640 ;
        RECT 903.510 17.580 903.830 17.640 ;
        RECT 900.750 17.440 903.830 17.580 ;
        RECT 900.750 17.380 901.070 17.440 ;
        RECT 903.510 17.380 903.830 17.440 ;
      LAYER via ;
        RECT 900.780 17.380 901.040 17.640 ;
        RECT 903.540 17.380 903.800 17.640 ;
      LAYER met2 ;
        RECT 903.600 17.670 903.740 54.000 ;
        RECT 900.780 17.350 901.040 17.670 ;
        RECT 903.540 17.350 903.800 17.670 ;
        RECT 900.840 2.400 900.980 17.350 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 918.690 17.580 919.010 17.640 ;
        RECT 923.750 17.580 924.070 17.640 ;
        RECT 918.690 17.440 924.070 17.580 ;
        RECT 918.690 17.380 919.010 17.440 ;
        RECT 923.750 17.380 924.070 17.440 ;
      LAYER via ;
        RECT 918.720 17.380 918.980 17.640 ;
        RECT 923.780 17.380 924.040 17.640 ;
      LAYER met2 ;
        RECT 923.840 17.670 923.980 54.000 ;
        RECT 918.720 17.350 918.980 17.670 ;
        RECT 923.780 17.350 924.040 17.670 ;
        RECT 918.780 2.400 918.920 17.350 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 938.100 17.410 938.240 54.000 ;
        RECT 936.260 17.270 938.240 17.410 ;
        RECT 936.260 2.400 936.400 17.270 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 954.110 15.200 954.430 15.260 ;
        RECT 958.710 15.200 959.030 15.260 ;
        RECT 954.110 15.060 959.030 15.200 ;
        RECT 954.110 15.000 954.430 15.060 ;
        RECT 958.710 15.000 959.030 15.060 ;
      LAYER via ;
        RECT 954.140 15.000 954.400 15.260 ;
        RECT 958.740 15.000 959.000 15.260 ;
      LAYER met2 ;
        RECT 958.800 15.290 958.940 54.000 ;
        RECT 954.140 14.970 954.400 15.290 ;
        RECT 958.740 14.970 959.000 15.290 ;
        RECT 954.200 2.400 954.340 14.970 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 972.140 2.400 972.280 54.000 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 650.970 17.580 651.290 17.640 ;
        RECT 650.970 17.440 728.020 17.580 ;
        RECT 650.970 17.380 651.290 17.440 ;
        RECT 727.880 16.900 728.020 17.440 ;
        RECT 753.090 16.900 753.410 16.960 ;
        RECT 727.880 16.760 753.410 16.900 ;
        RECT 753.090 16.700 753.410 16.760 ;
      LAYER via ;
        RECT 651.000 17.380 651.260 17.640 ;
        RECT 753.120 16.700 753.380 16.960 ;
      LAYER met2 ;
        RECT 651.000 17.350 651.260 17.670 ;
        RECT 651.060 2.400 651.200 17.350 ;
        RECT 753.180 16.990 753.320 54.000 ;
        RECT 753.120 16.670 753.380 16.990 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 989.990 17.580 990.310 17.640 ;
        RECT 993.210 17.580 993.530 17.640 ;
        RECT 989.990 17.440 993.530 17.580 ;
        RECT 989.990 17.380 990.310 17.440 ;
        RECT 993.210 17.380 993.530 17.440 ;
      LAYER via ;
        RECT 990.020 17.380 990.280 17.640 ;
        RECT 993.240 17.380 993.500 17.640 ;
      LAYER met2 ;
        RECT 993.300 17.670 993.440 54.000 ;
        RECT 990.020 17.350 990.280 17.670 ;
        RECT 993.240 17.350 993.500 17.670 ;
        RECT 990.080 2.400 990.220 17.350 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.470 17.920 1007.790 17.980 ;
        RECT 1013.450 17.920 1013.770 17.980 ;
        RECT 1007.470 17.780 1013.770 17.920 ;
        RECT 1007.470 17.720 1007.790 17.780 ;
        RECT 1013.450 17.720 1013.770 17.780 ;
      LAYER via ;
        RECT 1007.500 17.720 1007.760 17.980 ;
        RECT 1013.480 17.720 1013.740 17.980 ;
      LAYER met2 ;
        RECT 1013.540 18.010 1013.680 54.000 ;
        RECT 1007.500 17.690 1007.760 18.010 ;
        RECT 1013.480 17.690 1013.740 18.010 ;
        RECT 1007.560 2.400 1007.700 17.690 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1025.410 17.580 1025.730 17.640 ;
        RECT 1027.710 17.580 1028.030 17.640 ;
        RECT 1025.410 17.440 1028.030 17.580 ;
        RECT 1025.410 17.380 1025.730 17.440 ;
        RECT 1027.710 17.380 1028.030 17.440 ;
      LAYER via ;
        RECT 1025.440 17.380 1025.700 17.640 ;
        RECT 1027.740 17.380 1028.000 17.640 ;
      LAYER met2 ;
        RECT 1027.800 17.670 1027.940 54.000 ;
        RECT 1025.440 17.350 1025.700 17.670 ;
        RECT 1027.740 17.350 1028.000 17.670 ;
        RECT 1025.500 2.400 1025.640 17.350 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1043.350 17.580 1043.670 17.640 ;
        RECT 1048.410 17.580 1048.730 17.640 ;
        RECT 1043.350 17.440 1048.730 17.580 ;
        RECT 1043.350 17.380 1043.670 17.440 ;
        RECT 1048.410 17.380 1048.730 17.440 ;
      LAYER via ;
        RECT 1043.380 17.380 1043.640 17.640 ;
        RECT 1048.440 17.380 1048.700 17.640 ;
      LAYER met2 ;
        RECT 1048.500 17.670 1048.640 54.000 ;
        RECT 1043.380 17.350 1043.640 17.670 ;
        RECT 1048.440 17.350 1048.700 17.670 ;
        RECT 1043.440 2.400 1043.580 17.350 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1062.300 17.410 1062.440 54.000 ;
        RECT 1061.380 17.270 1062.440 17.410 ;
        RECT 1061.380 2.400 1061.520 17.270 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1079.230 17.580 1079.550 17.640 ;
        RECT 1082.910 17.580 1083.230 17.640 ;
        RECT 1079.230 17.440 1083.230 17.580 ;
        RECT 1079.230 17.380 1079.550 17.440 ;
        RECT 1082.910 17.380 1083.230 17.440 ;
      LAYER via ;
        RECT 1079.260 17.380 1079.520 17.640 ;
        RECT 1082.940 17.380 1083.200 17.640 ;
      LAYER met2 ;
        RECT 1083.000 17.670 1083.140 54.000 ;
        RECT 1079.260 17.350 1079.520 17.670 ;
        RECT 1082.940 17.350 1083.200 17.670 ;
        RECT 1079.320 2.400 1079.460 17.350 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.800 2.400 1096.940 54.000 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1114.650 17.580 1114.970 17.640 ;
        RECT 1117.410 17.580 1117.730 17.640 ;
        RECT 1114.650 17.440 1117.730 17.580 ;
        RECT 1114.650 17.380 1114.970 17.440 ;
        RECT 1117.410 17.380 1117.730 17.440 ;
      LAYER via ;
        RECT 1114.680 17.380 1114.940 17.640 ;
        RECT 1117.440 17.380 1117.700 17.640 ;
      LAYER met2 ;
        RECT 1117.500 17.670 1117.640 54.000 ;
        RECT 1114.680 17.350 1114.940 17.670 ;
        RECT 1117.440 17.350 1117.700 17.670 ;
        RECT 1114.740 2.400 1114.880 17.350 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1132.590 17.580 1132.910 17.640 ;
        RECT 1138.110 17.580 1138.430 17.640 ;
        RECT 1132.590 17.440 1138.430 17.580 ;
        RECT 1132.590 17.380 1132.910 17.440 ;
        RECT 1138.110 17.380 1138.430 17.440 ;
      LAYER via ;
        RECT 1132.620 17.380 1132.880 17.640 ;
        RECT 1138.140 17.380 1138.400 17.640 ;
      LAYER met2 ;
        RECT 1138.200 17.670 1138.340 54.000 ;
        RECT 1132.620 17.350 1132.880 17.670 ;
        RECT 1138.140 17.350 1138.400 17.670 ;
        RECT 1132.680 2.400 1132.820 17.350 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1152.000 17.410 1152.140 54.000 ;
        RECT 1150.620 17.270 1152.140 17.410 ;
        RECT 1150.620 2.400 1150.760 17.270 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 669.000 2.400 669.140 54.000 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1168.470 17.580 1168.790 17.640 ;
        RECT 1172.610 17.580 1172.930 17.640 ;
        RECT 1168.470 17.440 1172.930 17.580 ;
        RECT 1168.470 17.380 1168.790 17.440 ;
        RECT 1172.610 17.380 1172.930 17.440 ;
      LAYER via ;
        RECT 1168.500 17.380 1168.760 17.640 ;
        RECT 1172.640 17.380 1172.900 17.640 ;
      LAYER met2 ;
        RECT 1172.700 17.670 1172.840 54.000 ;
        RECT 1168.500 17.350 1168.760 17.670 ;
        RECT 1172.640 17.350 1172.900 17.670 ;
        RECT 1168.560 2.400 1168.700 17.350 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1186.040 2.400 1186.180 54.000 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1203.890 17.580 1204.210 17.640 ;
        RECT 1207.110 17.580 1207.430 17.640 ;
        RECT 1203.890 17.440 1207.430 17.580 ;
        RECT 1203.890 17.380 1204.210 17.440 ;
        RECT 1207.110 17.380 1207.430 17.440 ;
      LAYER via ;
        RECT 1203.920 17.380 1204.180 17.640 ;
        RECT 1207.140 17.380 1207.400 17.640 ;
      LAYER met2 ;
        RECT 1207.200 17.670 1207.340 54.000 ;
        RECT 1203.920 17.350 1204.180 17.670 ;
        RECT 1207.140 17.350 1207.400 17.670 ;
        RECT 1203.980 2.400 1204.120 17.350 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1221.830 17.920 1222.150 17.980 ;
        RECT 1227.810 17.920 1228.130 17.980 ;
        RECT 1221.830 17.780 1228.130 17.920 ;
        RECT 1221.830 17.720 1222.150 17.780 ;
        RECT 1227.810 17.720 1228.130 17.780 ;
      LAYER via ;
        RECT 1221.860 17.720 1222.120 17.980 ;
        RECT 1227.840 17.720 1228.100 17.980 ;
      LAYER met2 ;
        RECT 1227.900 18.010 1228.040 54.000 ;
        RECT 1221.860 17.690 1222.120 18.010 ;
        RECT 1227.840 17.690 1228.100 18.010 ;
        RECT 1221.920 2.400 1222.060 17.690 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1239.770 16.900 1240.090 16.960 ;
        RECT 1245.290 16.900 1245.610 16.960 ;
        RECT 1239.770 16.760 1245.610 16.900 ;
        RECT 1239.770 16.700 1240.090 16.760 ;
        RECT 1245.290 16.700 1245.610 16.760 ;
      LAYER via ;
        RECT 1239.800 16.700 1240.060 16.960 ;
        RECT 1245.320 16.700 1245.580 16.960 ;
      LAYER met2 ;
        RECT 1245.380 16.990 1245.520 54.000 ;
        RECT 1239.800 16.670 1240.060 16.990 ;
        RECT 1245.320 16.670 1245.580 16.990 ;
        RECT 1239.860 2.400 1240.000 16.670 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1257.250 17.580 1257.570 17.640 ;
        RECT 1262.310 17.580 1262.630 17.640 ;
        RECT 1257.250 17.440 1262.630 17.580 ;
        RECT 1257.250 17.380 1257.570 17.440 ;
        RECT 1262.310 17.380 1262.630 17.440 ;
      LAYER via ;
        RECT 1257.280 17.380 1257.540 17.640 ;
        RECT 1262.340 17.380 1262.600 17.640 ;
      LAYER met2 ;
        RECT 1262.400 17.670 1262.540 54.000 ;
        RECT 1257.280 17.350 1257.540 17.670 ;
        RECT 1262.340 17.350 1262.600 17.670 ;
        RECT 1257.340 2.400 1257.480 17.350 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1276.200 17.410 1276.340 54.000 ;
        RECT 1275.280 17.270 1276.340 17.410 ;
        RECT 1275.280 2.400 1275.420 17.270 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1293.130 17.580 1293.450 17.640 ;
        RECT 1296.810 17.580 1297.130 17.640 ;
        RECT 1293.130 17.440 1297.130 17.580 ;
        RECT 1293.130 17.380 1293.450 17.440 ;
        RECT 1296.810 17.380 1297.130 17.440 ;
      LAYER via ;
        RECT 1293.160 17.380 1293.420 17.640 ;
        RECT 1296.840 17.380 1297.100 17.640 ;
      LAYER met2 ;
        RECT 1296.900 17.670 1297.040 54.000 ;
        RECT 1293.160 17.350 1293.420 17.670 ;
        RECT 1296.840 17.350 1297.100 17.670 ;
        RECT 1293.220 2.400 1293.360 17.350 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.070 17.580 1311.390 17.640 ;
        RECT 1318.430 17.580 1318.750 17.640 ;
        RECT 1311.070 17.440 1318.750 17.580 ;
        RECT 1311.070 17.380 1311.390 17.440 ;
        RECT 1318.430 17.380 1318.750 17.440 ;
      LAYER via ;
        RECT 1311.100 17.380 1311.360 17.640 ;
        RECT 1318.460 17.380 1318.720 17.640 ;
      LAYER met2 ;
        RECT 1318.520 17.670 1318.660 54.000 ;
        RECT 1311.100 17.350 1311.360 17.670 ;
        RECT 1318.460 17.350 1318.720 17.670 ;
        RECT 1311.160 2.400 1311.300 17.350 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1329.010 17.580 1329.330 17.640 ;
        RECT 1331.310 17.580 1331.630 17.640 ;
        RECT 1329.010 17.440 1331.630 17.580 ;
        RECT 1329.010 17.380 1329.330 17.440 ;
        RECT 1331.310 17.380 1331.630 17.440 ;
      LAYER via ;
        RECT 1329.040 17.380 1329.300 17.640 ;
        RECT 1331.340 17.380 1331.600 17.640 ;
      LAYER met2 ;
        RECT 1331.400 17.670 1331.540 54.000 ;
        RECT 1329.040 17.350 1329.300 17.670 ;
        RECT 1331.340 17.350 1331.600 17.670 ;
        RECT 1329.100 2.400 1329.240 17.350 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 686.390 17.240 686.710 17.300 ;
        RECT 689.610 17.240 689.930 17.300 ;
        RECT 686.390 17.100 689.930 17.240 ;
        RECT 686.390 17.040 686.710 17.100 ;
        RECT 689.610 17.040 689.930 17.100 ;
      LAYER via ;
        RECT 686.420 17.040 686.680 17.300 ;
        RECT 689.640 17.040 689.900 17.300 ;
      LAYER met2 ;
        RECT 689.700 17.330 689.840 54.000 ;
        RECT 686.420 17.010 686.680 17.330 ;
        RECT 689.640 17.010 689.900 17.330 ;
        RECT 686.480 2.400 686.620 17.010 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.490 17.580 1346.810 17.640 ;
        RECT 1352.010 17.580 1352.330 17.640 ;
        RECT 1346.490 17.440 1352.330 17.580 ;
        RECT 1346.490 17.380 1346.810 17.440 ;
        RECT 1352.010 17.380 1352.330 17.440 ;
      LAYER via ;
        RECT 1346.520 17.380 1346.780 17.640 ;
        RECT 1352.040 17.380 1352.300 17.640 ;
      LAYER met2 ;
        RECT 1352.100 17.670 1352.240 54.000 ;
        RECT 1346.520 17.350 1346.780 17.670 ;
        RECT 1352.040 17.350 1352.300 17.670 ;
        RECT 1346.580 2.400 1346.720 17.350 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1364.430 17.580 1364.750 17.640 ;
        RECT 1366.730 17.580 1367.050 17.640 ;
        RECT 1364.430 17.440 1367.050 17.580 ;
        RECT 1364.430 17.380 1364.750 17.440 ;
        RECT 1366.730 17.380 1367.050 17.440 ;
      LAYER via ;
        RECT 1364.460 17.380 1364.720 17.640 ;
        RECT 1366.760 17.380 1367.020 17.640 ;
      LAYER met2 ;
        RECT 1366.820 17.670 1366.960 54.000 ;
        RECT 1364.460 17.350 1364.720 17.670 ;
        RECT 1366.760 17.350 1367.020 17.670 ;
        RECT 1364.520 2.400 1364.660 17.350 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1380.070 17.580 1380.390 17.640 ;
        RECT 1382.370 17.580 1382.690 17.640 ;
        RECT 1380.070 17.440 1382.690 17.580 ;
        RECT 1380.070 17.380 1380.390 17.440 ;
        RECT 1382.370 17.380 1382.690 17.440 ;
      LAYER via ;
        RECT 1380.100 17.380 1380.360 17.640 ;
        RECT 1382.400 17.380 1382.660 17.640 ;
      LAYER met2 ;
        RECT 1380.160 17.670 1380.300 54.000 ;
        RECT 1380.100 17.350 1380.360 17.670 ;
        RECT 1382.400 17.350 1382.660 17.670 ;
        RECT 1382.460 2.400 1382.600 17.350 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1394.330 17.920 1394.650 17.980 ;
        RECT 1400.310 17.920 1400.630 17.980 ;
        RECT 1394.330 17.780 1400.630 17.920 ;
        RECT 1394.330 17.720 1394.650 17.780 ;
        RECT 1400.310 17.720 1400.630 17.780 ;
      LAYER via ;
        RECT 1394.360 17.720 1394.620 17.980 ;
        RECT 1400.340 17.720 1400.600 17.980 ;
      LAYER met2 ;
        RECT 1394.420 18.010 1394.560 54.000 ;
        RECT 1394.360 17.690 1394.620 18.010 ;
        RECT 1400.340 17.690 1400.600 18.010 ;
        RECT 1400.400 2.400 1400.540 17.690 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1414.660 17.410 1414.800 54.000 ;
        RECT 1414.660 17.270 1418.480 17.410 ;
        RECT 1418.340 2.400 1418.480 17.270 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1434.900 20.640 1435.040 54.000 ;
        RECT 1434.900 20.500 1435.960 20.640 ;
        RECT 1435.820 2.400 1435.960 20.500 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1450.080 17.410 1450.220 54.000 ;
        RECT 1450.080 17.270 1453.900 17.410 ;
        RECT 1453.760 2.400 1453.900 17.270 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1462.410 17.580 1462.730 17.640 ;
        RECT 1471.610 17.580 1471.930 17.640 ;
        RECT 1462.410 17.440 1471.930 17.580 ;
        RECT 1462.410 17.380 1462.730 17.440 ;
        RECT 1471.610 17.380 1471.930 17.440 ;
      LAYER via ;
        RECT 1462.440 17.380 1462.700 17.640 ;
        RECT 1471.640 17.380 1471.900 17.640 ;
      LAYER met2 ;
        RECT 1462.500 17.670 1462.640 54.000 ;
        RECT 1462.440 17.350 1462.700 17.670 ;
        RECT 1471.640 17.350 1471.900 17.670 ;
        RECT 1471.700 2.400 1471.840 17.350 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1476.210 17.240 1476.530 17.300 ;
        RECT 1489.550 17.240 1489.870 17.300 ;
        RECT 1476.210 17.100 1489.870 17.240 ;
        RECT 1476.210 17.040 1476.530 17.100 ;
        RECT 1489.550 17.040 1489.870 17.100 ;
      LAYER via ;
        RECT 1476.240 17.040 1476.500 17.300 ;
        RECT 1489.580 17.040 1489.840 17.300 ;
      LAYER met2 ;
        RECT 1476.300 17.330 1476.440 54.000 ;
        RECT 1476.240 17.010 1476.500 17.330 ;
        RECT 1489.580 17.010 1489.840 17.330 ;
        RECT 1489.640 2.400 1489.780 17.010 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1496.910 15.200 1497.230 15.260 ;
        RECT 1507.030 15.200 1507.350 15.260 ;
        RECT 1496.910 15.060 1507.350 15.200 ;
        RECT 1496.910 15.000 1497.230 15.060 ;
        RECT 1507.030 15.000 1507.350 15.060 ;
      LAYER via ;
        RECT 1496.940 15.000 1497.200 15.260 ;
        RECT 1507.060 15.000 1507.320 15.260 ;
      LAYER met2 ;
        RECT 1497.000 15.290 1497.140 54.000 ;
        RECT 1496.940 14.970 1497.200 15.290 ;
        RECT 1507.060 14.970 1507.320 15.290 ;
        RECT 1507.120 2.400 1507.260 14.970 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 704.330 15.200 704.650 15.260 ;
        RECT 710.310 15.200 710.630 15.260 ;
        RECT 704.330 15.060 710.630 15.200 ;
        RECT 704.330 15.000 704.650 15.060 ;
        RECT 710.310 15.000 710.630 15.060 ;
      LAYER via ;
        RECT 704.360 15.000 704.620 15.260 ;
        RECT 710.340 15.000 710.600 15.260 ;
      LAYER met2 ;
        RECT 710.400 15.290 710.540 54.000 ;
        RECT 704.360 14.970 704.620 15.290 ;
        RECT 710.340 14.970 710.600 15.290 ;
        RECT 704.420 2.400 704.560 14.970 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1510.710 17.580 1511.030 17.640 ;
        RECT 1524.970 17.580 1525.290 17.640 ;
        RECT 1510.710 17.440 1525.290 17.580 ;
        RECT 1510.710 17.380 1511.030 17.440 ;
        RECT 1524.970 17.380 1525.290 17.440 ;
      LAYER via ;
        RECT 1510.740 17.380 1511.000 17.640 ;
        RECT 1525.000 17.380 1525.260 17.640 ;
      LAYER met2 ;
        RECT 1510.800 17.670 1510.940 54.000 ;
        RECT 1510.740 17.350 1511.000 17.670 ;
        RECT 1525.000 17.350 1525.260 17.670 ;
        RECT 1525.060 2.400 1525.200 17.350 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.510 20.640 1524.830 20.700 ;
        RECT 1542.910 20.640 1543.230 20.700 ;
        RECT 1524.510 20.500 1543.230 20.640 ;
        RECT 1524.510 20.440 1524.830 20.500 ;
        RECT 1542.910 20.440 1543.230 20.500 ;
      LAYER via ;
        RECT 1524.540 20.440 1524.800 20.700 ;
        RECT 1542.940 20.440 1543.200 20.700 ;
      LAYER met2 ;
        RECT 1524.600 20.730 1524.740 54.000 ;
        RECT 1524.540 20.410 1524.800 20.730 ;
        RECT 1542.940 20.410 1543.200 20.730 ;
        RECT 1543.000 2.400 1543.140 20.410 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1538.310 16.220 1538.630 16.280 ;
        RECT 1560.850 16.220 1561.170 16.280 ;
        RECT 1538.310 16.080 1561.170 16.220 ;
        RECT 1538.310 16.020 1538.630 16.080 ;
        RECT 1560.850 16.020 1561.170 16.080 ;
      LAYER via ;
        RECT 1538.340 16.020 1538.600 16.280 ;
        RECT 1560.880 16.020 1561.140 16.280 ;
      LAYER met2 ;
        RECT 1538.400 16.310 1538.540 54.000 ;
        RECT 1538.340 15.990 1538.600 16.310 ;
        RECT 1560.880 15.990 1561.140 16.310 ;
        RECT 1560.940 2.400 1561.080 15.990 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1551.650 16.900 1551.970 16.960 ;
        RECT 1578.790 16.900 1579.110 16.960 ;
        RECT 1551.650 16.760 1579.110 16.900 ;
        RECT 1551.650 16.700 1551.970 16.760 ;
        RECT 1578.790 16.700 1579.110 16.760 ;
      LAYER via ;
        RECT 1551.680 16.700 1551.940 16.960 ;
        RECT 1578.820 16.700 1579.080 16.960 ;
      LAYER met2 ;
        RECT 1551.740 16.990 1551.880 54.000 ;
        RECT 1551.680 16.670 1551.940 16.990 ;
        RECT 1578.820 16.670 1579.080 16.990 ;
        RECT 1578.880 2.400 1579.020 16.670 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1572.350 18.260 1572.670 18.320 ;
        RECT 1596.270 18.260 1596.590 18.320 ;
        RECT 1572.350 18.120 1596.590 18.260 ;
        RECT 1572.350 18.060 1572.670 18.120 ;
        RECT 1596.270 18.060 1596.590 18.120 ;
      LAYER via ;
        RECT 1572.380 18.060 1572.640 18.320 ;
        RECT 1596.300 18.060 1596.560 18.320 ;
      LAYER met2 ;
        RECT 1572.440 18.350 1572.580 54.000 ;
        RECT 1572.380 18.030 1572.640 18.350 ;
        RECT 1596.300 18.030 1596.560 18.350 ;
        RECT 1596.360 2.400 1596.500 18.030 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1586.610 17.580 1586.930 17.640 ;
        RECT 1614.210 17.580 1614.530 17.640 ;
        RECT 1586.610 17.440 1614.530 17.580 ;
        RECT 1586.610 17.380 1586.930 17.440 ;
        RECT 1614.210 17.380 1614.530 17.440 ;
      LAYER via ;
        RECT 1586.640 17.380 1586.900 17.640 ;
        RECT 1614.240 17.380 1614.500 17.640 ;
      LAYER met2 ;
        RECT 1586.700 17.670 1586.840 54.000 ;
        RECT 1586.640 17.350 1586.900 17.670 ;
        RECT 1614.240 17.350 1614.500 17.670 ;
        RECT 1614.300 2.400 1614.440 17.350 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1600.410 20.640 1600.730 20.700 ;
        RECT 1632.150 20.640 1632.470 20.700 ;
        RECT 1600.410 20.500 1632.470 20.640 ;
        RECT 1600.410 20.440 1600.730 20.500 ;
        RECT 1632.150 20.440 1632.470 20.500 ;
      LAYER via ;
        RECT 1600.440 20.440 1600.700 20.700 ;
        RECT 1632.180 20.440 1632.440 20.700 ;
      LAYER met2 ;
        RECT 1600.500 20.730 1600.640 54.000 ;
        RECT 1600.440 20.410 1600.700 20.730 ;
        RECT 1632.180 20.410 1632.440 20.730 ;
        RECT 1632.240 2.400 1632.380 20.410 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1613.750 17.240 1614.070 17.300 ;
        RECT 1650.090 17.240 1650.410 17.300 ;
        RECT 1613.750 17.100 1650.410 17.240 ;
        RECT 1613.750 17.040 1614.070 17.100 ;
        RECT 1650.090 17.040 1650.410 17.100 ;
      LAYER via ;
        RECT 1613.780 17.040 1614.040 17.300 ;
        RECT 1650.120 17.040 1650.380 17.300 ;
      LAYER met2 ;
        RECT 1613.840 17.330 1613.980 54.000 ;
        RECT 1613.780 17.010 1614.040 17.330 ;
        RECT 1650.120 17.010 1650.380 17.330 ;
        RECT 1650.180 2.400 1650.320 17.010 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1634.450 16.900 1634.770 16.960 ;
        RECT 1668.030 16.900 1668.350 16.960 ;
        RECT 1634.450 16.760 1668.350 16.900 ;
        RECT 1634.450 16.700 1634.770 16.760 ;
        RECT 1668.030 16.700 1668.350 16.760 ;
      LAYER via ;
        RECT 1634.480 16.700 1634.740 16.960 ;
        RECT 1668.060 16.700 1668.320 16.960 ;
      LAYER met2 ;
        RECT 1634.540 16.990 1634.680 54.000 ;
        RECT 1634.480 16.670 1634.740 16.990 ;
        RECT 1668.060 16.670 1668.320 16.990 ;
        RECT 1668.120 2.400 1668.260 16.670 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1648.710 14.860 1649.030 14.920 ;
        RECT 1685.510 14.860 1685.830 14.920 ;
        RECT 1648.710 14.720 1685.830 14.860 ;
        RECT 1648.710 14.660 1649.030 14.720 ;
        RECT 1685.510 14.660 1685.830 14.720 ;
      LAYER via ;
        RECT 1648.740 14.660 1649.000 14.920 ;
        RECT 1685.540 14.660 1685.800 14.920 ;
      LAYER met2 ;
        RECT 1648.800 14.950 1648.940 54.000 ;
        RECT 1648.740 14.630 1649.000 14.950 ;
        RECT 1685.540 14.630 1685.800 14.950 ;
        RECT 1685.600 2.400 1685.740 14.630 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 724.200 16.730 724.340 54.000 ;
        RECT 722.360 16.590 724.340 16.730 ;
        RECT 722.360 2.400 722.500 16.590 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1662.510 19.960 1662.830 20.020 ;
        RECT 1703.450 19.960 1703.770 20.020 ;
        RECT 1662.510 19.820 1703.770 19.960 ;
        RECT 1662.510 19.760 1662.830 19.820 ;
        RECT 1703.450 19.760 1703.770 19.820 ;
      LAYER via ;
        RECT 1662.540 19.760 1662.800 20.020 ;
        RECT 1703.480 19.760 1703.740 20.020 ;
      LAYER met2 ;
        RECT 1662.600 20.050 1662.740 54.000 ;
        RECT 1662.540 19.730 1662.800 20.050 ;
        RECT 1703.480 19.730 1703.740 20.050 ;
        RECT 1703.540 2.400 1703.680 19.730 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1676.310 19.620 1676.630 19.680 ;
        RECT 1721.390 19.620 1721.710 19.680 ;
        RECT 1676.310 19.480 1721.710 19.620 ;
        RECT 1676.310 19.420 1676.630 19.480 ;
        RECT 1721.390 19.420 1721.710 19.480 ;
      LAYER via ;
        RECT 1676.340 19.420 1676.600 19.680 ;
        RECT 1721.420 19.420 1721.680 19.680 ;
      LAYER met2 ;
        RECT 1676.400 19.710 1676.540 54.000 ;
        RECT 1676.340 19.390 1676.600 19.710 ;
        RECT 1721.420 19.390 1721.680 19.710 ;
        RECT 1721.480 2.400 1721.620 19.390 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1690.110 17.240 1690.430 17.300 ;
        RECT 1739.330 17.240 1739.650 17.300 ;
        RECT 1690.110 17.100 1739.650 17.240 ;
        RECT 1690.110 17.040 1690.430 17.100 ;
        RECT 1739.330 17.040 1739.650 17.100 ;
      LAYER via ;
        RECT 1690.140 17.040 1690.400 17.300 ;
        RECT 1739.360 17.040 1739.620 17.300 ;
      LAYER met2 ;
        RECT 1690.200 17.330 1690.340 54.000 ;
        RECT 1690.140 17.010 1690.400 17.330 ;
        RECT 1739.360 17.010 1739.620 17.330 ;
        RECT 1739.420 2.400 1739.560 17.010 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1710.350 19.960 1710.670 20.020 ;
        RECT 1756.810 19.960 1757.130 20.020 ;
        RECT 1710.350 19.820 1757.130 19.960 ;
        RECT 1710.350 19.760 1710.670 19.820 ;
        RECT 1756.810 19.760 1757.130 19.820 ;
      LAYER via ;
        RECT 1710.380 19.760 1710.640 20.020 ;
        RECT 1756.840 19.760 1757.100 20.020 ;
      LAYER met2 ;
        RECT 1710.440 20.050 1710.580 54.000 ;
        RECT 1710.380 19.730 1710.640 20.050 ;
        RECT 1756.840 19.730 1757.100 20.050 ;
        RECT 1756.900 2.400 1757.040 19.730 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1724.610 17.920 1724.930 17.980 ;
        RECT 1774.750 17.920 1775.070 17.980 ;
        RECT 1724.610 17.780 1775.070 17.920 ;
        RECT 1724.610 17.720 1724.930 17.780 ;
        RECT 1774.750 17.720 1775.070 17.780 ;
      LAYER via ;
        RECT 1724.640 17.720 1724.900 17.980 ;
        RECT 1774.780 17.720 1775.040 17.980 ;
      LAYER met2 ;
        RECT 1724.700 18.010 1724.840 54.000 ;
        RECT 1724.640 17.690 1724.900 18.010 ;
        RECT 1774.780 17.690 1775.040 18.010 ;
        RECT 1774.840 2.400 1774.980 17.690 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1738.410 19.620 1738.730 19.680 ;
        RECT 1792.690 19.620 1793.010 19.680 ;
        RECT 1738.410 19.480 1793.010 19.620 ;
        RECT 1738.410 19.420 1738.730 19.480 ;
        RECT 1792.690 19.420 1793.010 19.480 ;
      LAYER via ;
        RECT 1738.440 19.420 1738.700 19.680 ;
        RECT 1792.720 19.420 1792.980 19.680 ;
      LAYER met2 ;
        RECT 1738.500 19.710 1738.640 54.000 ;
        RECT 1738.440 19.390 1738.700 19.710 ;
        RECT 1792.720 19.390 1792.980 19.710 ;
        RECT 1792.780 2.400 1792.920 19.390 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1752.210 17.240 1752.530 17.300 ;
        RECT 1810.630 17.240 1810.950 17.300 ;
        RECT 1752.210 17.100 1810.950 17.240 ;
        RECT 1752.210 17.040 1752.530 17.100 ;
        RECT 1810.630 17.040 1810.950 17.100 ;
      LAYER via ;
        RECT 1752.240 17.040 1752.500 17.300 ;
        RECT 1810.660 17.040 1810.920 17.300 ;
      LAYER met2 ;
        RECT 1752.300 17.330 1752.440 54.000 ;
        RECT 1752.240 17.010 1752.500 17.330 ;
        RECT 1810.660 17.010 1810.920 17.330 ;
        RECT 1810.720 2.400 1810.860 17.010 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 19.960 1773.230 20.020 ;
        RECT 1828.570 19.960 1828.890 20.020 ;
        RECT 1772.910 19.820 1828.890 19.960 ;
        RECT 1772.910 19.760 1773.230 19.820 ;
        RECT 1828.570 19.760 1828.890 19.820 ;
      LAYER via ;
        RECT 1772.940 19.760 1773.200 20.020 ;
        RECT 1828.600 19.760 1828.860 20.020 ;
      LAYER met2 ;
        RECT 1773.000 20.050 1773.140 54.000 ;
        RECT 1772.940 19.730 1773.200 20.050 ;
        RECT 1828.600 19.730 1828.860 20.050 ;
        RECT 1828.660 2.400 1828.800 19.730 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1786.250 18.940 1786.570 19.000 ;
        RECT 1846.050 18.940 1846.370 19.000 ;
        RECT 1786.250 18.800 1846.370 18.940 ;
        RECT 1786.250 18.740 1786.570 18.800 ;
        RECT 1846.050 18.740 1846.370 18.800 ;
      LAYER via ;
        RECT 1786.280 18.740 1786.540 19.000 ;
        RECT 1846.080 18.740 1846.340 19.000 ;
      LAYER met2 ;
        RECT 1786.340 19.030 1786.480 54.000 ;
        RECT 1786.280 18.710 1786.540 19.030 ;
        RECT 1846.080 18.710 1846.340 19.030 ;
        RECT 1846.140 2.400 1846.280 18.710 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1800.510 19.620 1800.830 19.680 ;
        RECT 1863.990 19.620 1864.310 19.680 ;
        RECT 1800.510 19.480 1864.310 19.620 ;
        RECT 1800.510 19.420 1800.830 19.480 ;
        RECT 1863.990 19.420 1864.310 19.480 ;
      LAYER via ;
        RECT 1800.540 19.420 1800.800 19.680 ;
        RECT 1864.020 19.420 1864.280 19.680 ;
      LAYER met2 ;
        RECT 1800.600 19.710 1800.740 54.000 ;
        RECT 1800.540 19.390 1800.800 19.710 ;
        RECT 1864.020 19.390 1864.280 19.710 ;
        RECT 1864.080 2.400 1864.220 19.390 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 740.210 17.580 740.530 17.640 ;
        RECT 744.810 17.580 745.130 17.640 ;
        RECT 740.210 17.440 745.130 17.580 ;
        RECT 740.210 17.380 740.530 17.440 ;
        RECT 744.810 17.380 745.130 17.440 ;
      LAYER via ;
        RECT 740.240 17.380 740.500 17.640 ;
        RECT 744.840 17.380 745.100 17.640 ;
      LAYER met2 ;
        RECT 744.900 17.670 745.040 54.000 ;
        RECT 740.240 17.350 740.500 17.670 ;
        RECT 744.840 17.350 745.100 17.670 ;
        RECT 740.300 2.400 740.440 17.350 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1814.310 20.640 1814.630 20.700 ;
        RECT 1881.930 20.640 1882.250 20.700 ;
        RECT 1814.310 20.500 1882.250 20.640 ;
        RECT 1814.310 20.440 1814.630 20.500 ;
        RECT 1881.930 20.440 1882.250 20.500 ;
      LAYER via ;
        RECT 1814.340 20.440 1814.600 20.700 ;
        RECT 1881.960 20.440 1882.220 20.700 ;
      LAYER met2 ;
        RECT 1814.400 20.730 1814.540 54.000 ;
        RECT 1814.340 20.410 1814.600 20.730 ;
        RECT 1881.960 20.410 1882.220 20.730 ;
        RECT 1882.020 2.400 1882.160 20.410 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1828.110 17.240 1828.430 17.300 ;
        RECT 1899.870 17.240 1900.190 17.300 ;
        RECT 1828.110 17.100 1900.190 17.240 ;
        RECT 1828.110 17.040 1828.430 17.100 ;
        RECT 1899.870 17.040 1900.190 17.100 ;
      LAYER via ;
        RECT 1828.140 17.040 1828.400 17.300 ;
        RECT 1899.900 17.040 1900.160 17.300 ;
      LAYER met2 ;
        RECT 1828.200 17.330 1828.340 54.000 ;
        RECT 1828.140 17.010 1828.400 17.330 ;
        RECT 1899.900 17.010 1900.160 17.330 ;
        RECT 1899.960 2.400 1900.100 17.010 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1848.350 16.560 1848.670 16.620 ;
        RECT 1917.810 16.560 1918.130 16.620 ;
        RECT 1848.350 16.420 1918.130 16.560 ;
        RECT 1848.350 16.360 1848.670 16.420 ;
        RECT 1917.810 16.360 1918.130 16.420 ;
      LAYER via ;
        RECT 1848.380 16.360 1848.640 16.620 ;
        RECT 1917.840 16.360 1918.100 16.620 ;
      LAYER met2 ;
        RECT 1848.440 16.650 1848.580 54.000 ;
        RECT 1848.380 16.330 1848.640 16.650 ;
        RECT 1917.840 16.330 1918.100 16.650 ;
        RECT 1917.900 2.400 1918.040 16.330 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1862.610 17.920 1862.930 17.980 ;
        RECT 1935.290 17.920 1935.610 17.980 ;
        RECT 1862.610 17.780 1935.610 17.920 ;
        RECT 1862.610 17.720 1862.930 17.780 ;
        RECT 1935.290 17.720 1935.610 17.780 ;
      LAYER via ;
        RECT 1862.640 17.720 1862.900 17.980 ;
        RECT 1935.320 17.720 1935.580 17.980 ;
      LAYER met2 ;
        RECT 1862.700 18.010 1862.840 54.000 ;
        RECT 1862.640 17.690 1862.900 18.010 ;
        RECT 1935.320 17.690 1935.580 18.010 ;
        RECT 1935.380 2.400 1935.520 17.690 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1876.410 18.600 1876.730 18.660 ;
        RECT 1953.230 18.600 1953.550 18.660 ;
        RECT 1876.410 18.460 1953.550 18.600 ;
        RECT 1876.410 18.400 1876.730 18.460 ;
        RECT 1953.230 18.400 1953.550 18.460 ;
      LAYER via ;
        RECT 1876.440 18.400 1876.700 18.660 ;
        RECT 1953.260 18.400 1953.520 18.660 ;
      LAYER met2 ;
        RECT 1876.500 18.690 1876.640 54.000 ;
        RECT 1876.440 18.370 1876.700 18.690 ;
        RECT 1953.260 18.370 1953.520 18.690 ;
        RECT 1953.320 2.400 1953.460 18.370 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1890.210 19.620 1890.530 19.680 ;
        RECT 1971.170 19.620 1971.490 19.680 ;
        RECT 1890.210 19.480 1971.490 19.620 ;
        RECT 1890.210 19.420 1890.530 19.480 ;
        RECT 1971.170 19.420 1971.490 19.480 ;
      LAYER via ;
        RECT 1890.240 19.420 1890.500 19.680 ;
        RECT 1971.200 19.420 1971.460 19.680 ;
      LAYER met2 ;
        RECT 1890.300 19.710 1890.440 54.000 ;
        RECT 1890.240 19.390 1890.500 19.710 ;
        RECT 1971.200 19.390 1971.460 19.710 ;
        RECT 1971.260 2.400 1971.400 19.390 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1903.550 17.240 1903.870 17.300 ;
        RECT 1989.110 17.240 1989.430 17.300 ;
        RECT 1903.550 17.100 1989.430 17.240 ;
        RECT 1903.550 17.040 1903.870 17.100 ;
        RECT 1989.110 17.040 1989.430 17.100 ;
      LAYER via ;
        RECT 1903.580 17.040 1903.840 17.300 ;
        RECT 1989.140 17.040 1989.400 17.300 ;
      LAYER met2 ;
        RECT 1903.640 17.330 1903.780 54.000 ;
        RECT 1903.580 17.010 1903.840 17.330 ;
        RECT 1989.140 17.010 1989.400 17.330 ;
        RECT 1989.200 2.400 1989.340 17.010 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1924.250 14.860 1924.570 14.920 ;
        RECT 2006.590 14.860 2006.910 14.920 ;
        RECT 1924.250 14.720 2006.910 14.860 ;
        RECT 1924.250 14.660 1924.570 14.720 ;
        RECT 2006.590 14.660 2006.910 14.720 ;
      LAYER via ;
        RECT 1924.280 14.660 1924.540 14.920 ;
        RECT 2006.620 14.660 2006.880 14.920 ;
      LAYER met2 ;
        RECT 1924.340 14.950 1924.480 54.000 ;
        RECT 1924.280 14.630 1924.540 14.950 ;
        RECT 2006.620 14.630 2006.880 14.950 ;
        RECT 2006.680 2.400 2006.820 14.630 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1938.510 18.940 1938.830 19.000 ;
        RECT 2024.530 18.940 2024.850 19.000 ;
        RECT 1938.510 18.800 2024.850 18.940 ;
        RECT 1938.510 18.740 1938.830 18.800 ;
        RECT 2024.530 18.740 2024.850 18.800 ;
      LAYER via ;
        RECT 1938.540 18.740 1938.800 19.000 ;
        RECT 2024.560 18.740 2024.820 19.000 ;
      LAYER met2 ;
        RECT 1938.600 19.030 1938.740 54.000 ;
        RECT 1938.540 18.710 1938.800 19.030 ;
        RECT 2024.560 18.710 2024.820 19.030 ;
        RECT 2024.620 2.400 2024.760 18.710 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1952.310 19.960 1952.630 20.020 ;
        RECT 2042.470 19.960 2042.790 20.020 ;
        RECT 1952.310 19.820 2042.790 19.960 ;
        RECT 1952.310 19.760 1952.630 19.820 ;
        RECT 2042.470 19.760 2042.790 19.820 ;
      LAYER via ;
        RECT 1952.340 19.760 1952.600 20.020 ;
        RECT 2042.500 19.760 2042.760 20.020 ;
      LAYER met2 ;
        RECT 1952.400 20.050 1952.540 54.000 ;
        RECT 1952.340 19.730 1952.600 20.050 ;
        RECT 2042.500 19.730 2042.760 20.050 ;
        RECT 2042.560 2.400 2042.700 19.730 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 758.240 17.410 758.380 54.000 ;
        RECT 757.780 17.270 758.380 17.410 ;
        RECT 757.780 2.400 757.920 17.270 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1965.650 17.580 1965.970 17.640 ;
        RECT 2060.410 17.580 2060.730 17.640 ;
        RECT 1965.650 17.440 2060.730 17.580 ;
        RECT 1965.650 17.380 1965.970 17.440 ;
        RECT 2060.410 17.380 2060.730 17.440 ;
      LAYER via ;
        RECT 1965.680 17.380 1965.940 17.640 ;
        RECT 2060.440 17.380 2060.700 17.640 ;
      LAYER met2 ;
        RECT 1965.740 17.670 1965.880 54.000 ;
        RECT 1965.680 17.350 1965.940 17.670 ;
        RECT 2060.440 17.350 2060.700 17.670 ;
        RECT 2060.500 2.400 2060.640 17.350 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1986.350 19.620 1986.670 19.680 ;
        RECT 2078.350 19.620 2078.670 19.680 ;
        RECT 1986.350 19.480 2078.670 19.620 ;
        RECT 1986.350 19.420 1986.670 19.480 ;
        RECT 2078.350 19.420 2078.670 19.480 ;
      LAYER via ;
        RECT 1986.380 19.420 1986.640 19.680 ;
        RECT 2078.380 19.420 2078.640 19.680 ;
      LAYER met2 ;
        RECT 1986.440 19.710 1986.580 54.000 ;
        RECT 1986.380 19.390 1986.640 19.710 ;
        RECT 2078.380 19.390 2078.640 19.710 ;
        RECT 2078.440 2.400 2078.580 19.390 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2091.230 2.960 2091.550 3.020 ;
        RECT 2095.830 2.960 2096.150 3.020 ;
        RECT 2091.230 2.820 2096.150 2.960 ;
        RECT 2091.230 2.760 2091.550 2.820 ;
        RECT 2095.830 2.760 2096.150 2.820 ;
      LAYER via ;
        RECT 2091.260 2.760 2091.520 3.020 ;
        RECT 2095.860 2.760 2096.120 3.020 ;
      LAYER met2 ;
        RECT 2091.320 3.050 2091.460 54.000 ;
        RECT 2091.260 2.730 2091.520 3.050 ;
        RECT 2095.860 2.730 2096.120 3.050 ;
        RECT 2095.920 2.400 2096.060 2.730 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2112.020 3.130 2112.160 54.000 ;
        RECT 2112.020 2.990 2114.000 3.130 ;
        RECT 2113.860 2.400 2114.000 2.990 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2125.730 17.240 2126.050 17.300 ;
        RECT 2131.710 17.240 2132.030 17.300 ;
        RECT 2125.730 17.100 2132.030 17.240 ;
        RECT 2125.730 17.040 2126.050 17.100 ;
        RECT 2131.710 17.040 2132.030 17.100 ;
      LAYER via ;
        RECT 2125.760 17.040 2126.020 17.300 ;
        RECT 2131.740 17.040 2132.000 17.300 ;
      LAYER met2 ;
        RECT 2125.820 17.330 2125.960 54.000 ;
        RECT 2125.760 17.010 2126.020 17.330 ;
        RECT 2131.740 17.010 2132.000 17.330 ;
        RECT 2131.800 2.400 2131.940 17.010 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2145.970 2.960 2146.290 3.020 ;
        RECT 2149.650 2.960 2149.970 3.020 ;
        RECT 2145.970 2.820 2149.970 2.960 ;
        RECT 2145.970 2.760 2146.290 2.820 ;
        RECT 2149.650 2.760 2149.970 2.820 ;
      LAYER via ;
        RECT 2146.000 2.760 2146.260 3.020 ;
        RECT 2149.680 2.760 2149.940 3.020 ;
      LAYER met2 ;
        RECT 2146.060 3.050 2146.200 54.000 ;
        RECT 2146.000 2.730 2146.260 3.050 ;
        RECT 2149.680 2.730 2149.940 3.050 ;
        RECT 2149.740 2.400 2149.880 2.730 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.220 17.410 2167.360 54.000 ;
        RECT 2167.220 17.270 2167.820 17.410 ;
        RECT 2167.680 2.400 2167.820 17.270 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.930 2.960 2181.250 3.020 ;
        RECT 2185.070 2.960 2185.390 3.020 ;
        RECT 2180.930 2.820 2185.390 2.960 ;
        RECT 2180.930 2.760 2181.250 2.820 ;
        RECT 2185.070 2.760 2185.390 2.820 ;
      LAYER via ;
        RECT 2180.960 2.760 2181.220 3.020 ;
        RECT 2185.100 2.760 2185.360 3.020 ;
      LAYER met2 ;
        RECT 2181.020 3.050 2181.160 54.000 ;
        RECT 2180.960 2.730 2181.220 3.050 ;
        RECT 2185.100 2.730 2185.360 3.050 ;
        RECT 2185.160 2.400 2185.300 2.730 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2201.720 3.130 2201.860 54.000 ;
        RECT 2201.720 2.990 2203.240 3.130 ;
        RECT 2203.100 2.400 2203.240 2.990 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2215.980 16.050 2216.120 54.000 ;
        RECT 2215.980 15.910 2221.180 16.050 ;
        RECT 2221.040 2.400 2221.180 15.910 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 775.630 17.580 775.950 17.640 ;
        RECT 779.310 17.580 779.630 17.640 ;
        RECT 775.630 17.440 779.630 17.580 ;
        RECT 775.630 17.380 775.950 17.440 ;
        RECT 779.310 17.380 779.630 17.440 ;
      LAYER via ;
        RECT 775.660 17.380 775.920 17.640 ;
        RECT 779.340 17.380 779.600 17.640 ;
      LAYER met2 ;
        RECT 779.400 17.670 779.540 54.000 ;
        RECT 775.660 17.350 775.920 17.670 ;
        RECT 779.340 17.350 779.600 17.670 ;
        RECT 775.720 2.400 775.860 17.350 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2235.670 2.960 2235.990 3.020 ;
        RECT 2238.890 2.960 2239.210 3.020 ;
        RECT 2235.670 2.820 2239.210 2.960 ;
        RECT 2235.670 2.760 2235.990 2.820 ;
        RECT 2238.890 2.760 2239.210 2.820 ;
      LAYER via ;
        RECT 2235.700 2.760 2235.960 3.020 ;
        RECT 2238.920 2.760 2239.180 3.020 ;
      LAYER met2 ;
        RECT 2235.760 3.050 2235.900 54.000 ;
        RECT 2235.700 2.730 2235.960 3.050 ;
        RECT 2238.920 2.730 2239.180 3.050 ;
        RECT 2238.980 2.400 2239.120 2.730 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2257.380 3.130 2257.520 54.000 ;
        RECT 2256.920 2.990 2257.520 3.130 ;
        RECT 2256.920 2.960 2257.060 2.990 ;
        RECT 2256.460 2.820 2257.060 2.960 ;
        RECT 2256.460 2.400 2256.600 2.820 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2271.090 2.960 2271.410 3.020 ;
        RECT 2274.310 2.960 2274.630 3.020 ;
        RECT 2271.090 2.820 2274.630 2.960 ;
        RECT 2271.090 2.760 2271.410 2.820 ;
        RECT 2274.310 2.760 2274.630 2.820 ;
      LAYER via ;
        RECT 2271.120 2.760 2271.380 3.020 ;
        RECT 2274.340 2.760 2274.600 3.020 ;
      LAYER met2 ;
        RECT 2271.180 3.050 2271.320 54.000 ;
        RECT 2271.120 2.730 2271.380 3.050 ;
        RECT 2274.340 2.730 2274.600 3.050 ;
        RECT 2274.400 2.400 2274.540 2.730 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2291.880 2.960 2292.020 54.000 ;
        RECT 2291.880 2.820 2292.480 2.960 ;
        RECT 2292.340 2.400 2292.480 2.820 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2305.130 2.960 2305.450 3.020 ;
        RECT 2310.190 2.960 2310.510 3.020 ;
        RECT 2305.130 2.820 2310.510 2.960 ;
        RECT 2305.130 2.760 2305.450 2.820 ;
        RECT 2310.190 2.760 2310.510 2.820 ;
      LAYER via ;
        RECT 2305.160 2.760 2305.420 3.020 ;
        RECT 2310.220 2.760 2310.480 3.020 ;
      LAYER met2 ;
        RECT 2305.220 3.050 2305.360 54.000 ;
        RECT 2305.160 2.730 2305.420 3.050 ;
        RECT 2310.220 2.730 2310.480 3.050 ;
        RECT 2310.280 2.400 2310.420 2.730 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2325.920 3.130 2326.060 54.000 ;
        RECT 2325.920 2.990 2328.360 3.130 ;
        RECT 2328.220 2.400 2328.360 2.990 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2339.630 17.580 2339.950 17.640 ;
        RECT 2345.610 17.580 2345.930 17.640 ;
        RECT 2339.630 17.440 2345.930 17.580 ;
        RECT 2339.630 17.380 2339.950 17.440 ;
        RECT 2345.610 17.380 2345.930 17.440 ;
      LAYER via ;
        RECT 2339.660 17.380 2339.920 17.640 ;
        RECT 2345.640 17.380 2345.900 17.640 ;
      LAYER met2 ;
        RECT 2339.720 17.670 2339.860 54.000 ;
        RECT 2339.660 17.350 2339.920 17.670 ;
        RECT 2345.640 17.350 2345.900 17.670 ;
        RECT 2345.700 2.400 2345.840 17.350 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2360.330 2.960 2360.650 3.020 ;
        RECT 2363.550 2.960 2363.870 3.020 ;
        RECT 2360.330 2.820 2363.870 2.960 ;
        RECT 2360.330 2.760 2360.650 2.820 ;
        RECT 2363.550 2.760 2363.870 2.820 ;
      LAYER via ;
        RECT 2360.360 2.760 2360.620 3.020 ;
        RECT 2363.580 2.760 2363.840 3.020 ;
      LAYER met2 ;
        RECT 2360.420 3.050 2360.560 54.000 ;
        RECT 2360.360 2.730 2360.620 3.050 ;
        RECT 2363.580 2.730 2363.840 3.050 ;
        RECT 2363.640 2.400 2363.780 2.730 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2241.650 24.040 2241.970 24.100 ;
        RECT 2381.490 24.040 2381.810 24.100 ;
        RECT 2241.650 23.900 2381.810 24.040 ;
        RECT 2241.650 23.840 2241.970 23.900 ;
        RECT 2381.490 23.840 2381.810 23.900 ;
      LAYER via ;
        RECT 2241.680 23.840 2241.940 24.100 ;
        RECT 2381.520 23.840 2381.780 24.100 ;
      LAYER met2 ;
        RECT 2241.740 24.130 2241.880 54.000 ;
        RECT 2241.680 23.810 2241.940 24.130 ;
        RECT 2381.520 23.810 2381.780 24.130 ;
        RECT 2381.580 2.400 2381.720 23.810 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2261.430 15.200 2261.750 15.260 ;
        RECT 2399.430 15.200 2399.750 15.260 ;
        RECT 2261.430 15.060 2399.750 15.200 ;
        RECT 2261.430 15.000 2261.750 15.060 ;
        RECT 2399.430 15.000 2399.750 15.060 ;
      LAYER via ;
        RECT 2261.460 15.000 2261.720 15.260 ;
        RECT 2399.460 15.000 2399.720 15.260 ;
      LAYER met2 ;
        RECT 2262.440 34.410 2262.580 54.000 ;
        RECT 2261.520 34.270 2262.580 34.410 ;
        RECT 2261.520 15.290 2261.660 34.270 ;
        RECT 2261.460 14.970 2261.720 15.290 ;
        RECT 2399.460 14.970 2399.720 15.290 ;
        RECT 2399.520 2.400 2399.660 14.970 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.570 17.920 793.890 17.980 ;
        RECT 799.550 17.920 799.870 17.980 ;
        RECT 793.570 17.780 799.870 17.920 ;
        RECT 793.570 17.720 793.890 17.780 ;
        RECT 799.550 17.720 799.870 17.780 ;
      LAYER via ;
        RECT 793.600 17.720 793.860 17.980 ;
        RECT 799.580 17.720 799.840 17.980 ;
      LAYER met2 ;
        RECT 799.640 18.010 799.780 54.000 ;
        RECT 793.600 17.690 793.860 18.010 ;
        RECT 799.580 17.690 799.840 18.010 ;
        RECT 793.660 2.400 793.800 17.690 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 639.010 17.920 639.330 17.980 ;
        RECT 745.270 17.920 745.590 17.980 ;
        RECT 639.010 17.780 745.590 17.920 ;
        RECT 639.010 17.720 639.330 17.780 ;
        RECT 745.270 17.720 745.590 17.780 ;
      LAYER via ;
        RECT 639.040 17.720 639.300 17.980 ;
        RECT 745.300 17.720 745.560 17.980 ;
      LAYER met2 ;
        RECT 745.360 18.010 745.500 54.000 ;
        RECT 639.040 17.690 639.300 18.010 ;
        RECT 745.300 17.690 745.560 18.010 ;
        RECT 639.100 2.400 639.240 17.690 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2276.610 17.240 2276.930 17.300 ;
        RECT 2422.890 17.240 2423.210 17.300 ;
        RECT 2276.610 17.100 2423.210 17.240 ;
        RECT 2276.610 17.040 2276.930 17.100 ;
        RECT 2422.890 17.040 2423.210 17.100 ;
      LAYER via ;
        RECT 2276.640 17.040 2276.900 17.300 ;
        RECT 2422.920 17.040 2423.180 17.300 ;
      LAYER met2 ;
        RECT 2276.700 17.330 2276.840 54.000 ;
        RECT 2276.640 17.010 2276.900 17.330 ;
        RECT 2422.920 17.010 2423.180 17.330 ;
        RECT 2422.980 2.400 2423.120 17.010 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2296.850 15.540 2297.170 15.600 ;
        RECT 2440.830 15.540 2441.150 15.600 ;
        RECT 2296.850 15.400 2441.150 15.540 ;
        RECT 2296.850 15.340 2297.170 15.400 ;
        RECT 2440.830 15.340 2441.150 15.400 ;
      LAYER via ;
        RECT 2296.880 15.340 2297.140 15.600 ;
        RECT 2440.860 15.340 2441.120 15.600 ;
      LAYER met2 ;
        RECT 2296.940 15.630 2297.080 54.000 ;
        RECT 2296.880 15.310 2297.140 15.630 ;
        RECT 2440.860 15.310 2441.120 15.630 ;
        RECT 2440.920 2.400 2441.060 15.310 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2346.990 16.900 2347.310 16.960 ;
        RECT 2458.770 16.900 2459.090 16.960 ;
        RECT 2346.990 16.760 2459.090 16.900 ;
        RECT 2346.990 16.700 2347.310 16.760 ;
        RECT 2458.770 16.700 2459.090 16.760 ;
        RECT 2311.110 15.880 2311.430 15.940 ;
        RECT 2346.990 15.880 2347.310 15.940 ;
        RECT 2311.110 15.740 2347.310 15.880 ;
        RECT 2311.110 15.680 2311.430 15.740 ;
        RECT 2346.990 15.680 2347.310 15.740 ;
      LAYER via ;
        RECT 2347.020 16.700 2347.280 16.960 ;
        RECT 2458.800 16.700 2459.060 16.960 ;
        RECT 2311.140 15.680 2311.400 15.940 ;
        RECT 2347.020 15.680 2347.280 15.940 ;
      LAYER met2 ;
        RECT 2311.200 15.970 2311.340 54.000 ;
        RECT 2347.020 16.670 2347.280 16.990 ;
        RECT 2458.800 16.670 2459.060 16.990 ;
        RECT 2347.080 15.970 2347.220 16.670 ;
        RECT 2311.140 15.650 2311.400 15.970 ;
        RECT 2347.020 15.650 2347.280 15.970 ;
        RECT 2458.860 2.400 2459.000 16.670 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2324.910 19.960 2325.230 20.020 ;
        RECT 2347.450 19.960 2347.770 20.020 ;
        RECT 2324.910 19.820 2347.770 19.960 ;
        RECT 2324.910 19.760 2325.230 19.820 ;
        RECT 2347.450 19.760 2347.770 19.820 ;
        RECT 2347.450 15.880 2347.770 15.940 ;
        RECT 2476.710 15.880 2477.030 15.940 ;
        RECT 2347.450 15.740 2477.030 15.880 ;
        RECT 2347.450 15.680 2347.770 15.740 ;
        RECT 2476.710 15.680 2477.030 15.740 ;
      LAYER via ;
        RECT 2324.940 19.760 2325.200 20.020 ;
        RECT 2347.480 19.760 2347.740 20.020 ;
        RECT 2347.480 15.680 2347.740 15.940 ;
        RECT 2476.740 15.680 2477.000 15.940 ;
      LAYER met2 ;
        RECT 2325.000 20.050 2325.140 54.000 ;
        RECT 2324.940 19.730 2325.200 20.050 ;
        RECT 2347.480 19.730 2347.740 20.050 ;
        RECT 2347.540 15.970 2347.680 19.730 ;
        RECT 2347.480 15.650 2347.740 15.970 ;
        RECT 2476.740 15.650 2477.000 15.970 ;
        RECT 2476.800 2.400 2476.940 15.650 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2338.710 17.920 2339.030 17.980 ;
        RECT 2338.710 17.780 2346.300 17.920 ;
        RECT 2338.710 17.720 2339.030 17.780 ;
        RECT 2346.160 17.580 2346.300 17.780 ;
        RECT 2494.650 17.580 2494.970 17.640 ;
        RECT 2346.160 17.440 2494.970 17.580 ;
        RECT 2494.650 17.380 2494.970 17.440 ;
      LAYER via ;
        RECT 2338.740 17.720 2339.000 17.980 ;
        RECT 2494.680 17.380 2494.940 17.640 ;
      LAYER met2 ;
        RECT 2338.800 18.010 2338.940 54.000 ;
        RECT 2338.740 17.690 2339.000 18.010 ;
        RECT 2494.680 17.350 2494.940 17.670 ;
        RECT 2494.740 2.400 2494.880 17.350 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2359.410 19.960 2359.730 20.020 ;
        RECT 2512.130 19.960 2512.450 20.020 ;
        RECT 2359.410 19.820 2512.450 19.960 ;
        RECT 2359.410 19.760 2359.730 19.820 ;
        RECT 2512.130 19.760 2512.450 19.820 ;
      LAYER via ;
        RECT 2359.440 19.760 2359.700 20.020 ;
        RECT 2512.160 19.760 2512.420 20.020 ;
      LAYER met2 ;
        RECT 2359.500 20.050 2359.640 54.000 ;
        RECT 2359.440 19.730 2359.700 20.050 ;
        RECT 2512.160 19.730 2512.420 20.050 ;
        RECT 2512.220 2.400 2512.360 19.730 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2373.210 20.300 2373.530 20.360 ;
        RECT 2530.070 20.300 2530.390 20.360 ;
        RECT 2373.210 20.160 2530.390 20.300 ;
        RECT 2373.210 20.100 2373.530 20.160 ;
        RECT 2530.070 20.100 2530.390 20.160 ;
      LAYER via ;
        RECT 2373.240 20.100 2373.500 20.360 ;
        RECT 2530.100 20.100 2530.360 20.360 ;
      LAYER met2 ;
        RECT 2373.300 20.390 2373.440 54.000 ;
        RECT 2373.240 20.070 2373.500 20.390 ;
        RECT 2530.100 20.070 2530.360 20.390 ;
        RECT 2530.160 2.400 2530.300 20.070 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2536.510 19.960 2536.830 20.020 ;
        RECT 2521.880 19.820 2536.830 19.960 ;
        RECT 2387.010 19.620 2387.330 19.680 ;
        RECT 2521.880 19.620 2522.020 19.820 ;
        RECT 2536.510 19.760 2536.830 19.820 ;
        RECT 2387.010 19.480 2522.020 19.620 ;
        RECT 2387.010 19.420 2387.330 19.480 ;
        RECT 2536.510 16.900 2536.830 16.960 ;
        RECT 2548.010 16.900 2548.330 16.960 ;
        RECT 2536.510 16.760 2548.330 16.900 ;
        RECT 2536.510 16.700 2536.830 16.760 ;
        RECT 2548.010 16.700 2548.330 16.760 ;
      LAYER via ;
        RECT 2387.040 19.420 2387.300 19.680 ;
        RECT 2536.540 19.760 2536.800 20.020 ;
        RECT 2536.540 16.700 2536.800 16.960 ;
        RECT 2548.040 16.700 2548.300 16.960 ;
      LAYER met2 ;
        RECT 2387.100 19.710 2387.240 54.000 ;
        RECT 2536.540 19.730 2536.800 20.050 ;
        RECT 2387.040 19.390 2387.300 19.710 ;
        RECT 2536.600 16.990 2536.740 19.730 ;
        RECT 2536.540 16.670 2536.800 16.990 ;
        RECT 2548.040 16.670 2548.300 16.990 ;
        RECT 2548.100 2.400 2548.240 16.670 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2400.810 20.640 2401.130 20.700 ;
        RECT 2400.810 20.500 2537.660 20.640 ;
        RECT 2400.810 20.440 2401.130 20.500 ;
        RECT 2537.520 19.620 2537.660 20.500 ;
        RECT 2565.950 19.620 2566.270 19.680 ;
        RECT 2537.520 19.480 2566.270 19.620 ;
        RECT 2565.950 19.420 2566.270 19.480 ;
      LAYER via ;
        RECT 2400.840 20.440 2401.100 20.700 ;
        RECT 2565.980 19.420 2566.240 19.680 ;
      LAYER met2 ;
        RECT 2400.900 20.730 2401.040 54.000 ;
        RECT 2400.840 20.410 2401.100 20.730 ;
        RECT 2565.980 19.390 2566.240 19.710 ;
        RECT 2566.040 2.400 2566.180 19.390 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2414.610 18.260 2414.930 18.320 ;
        RECT 2583.890 18.260 2584.210 18.320 ;
        RECT 2414.610 18.120 2584.210 18.260 ;
        RECT 2414.610 18.060 2414.930 18.120 ;
        RECT 2583.890 18.060 2584.210 18.120 ;
      LAYER via ;
        RECT 2414.640 18.060 2414.900 18.320 ;
        RECT 2583.920 18.060 2584.180 18.320 ;
      LAYER met2 ;
        RECT 2414.700 18.350 2414.840 54.000 ;
        RECT 2414.640 18.030 2414.900 18.350 ;
        RECT 2583.920 18.030 2584.180 18.350 ;
        RECT 2583.980 2.400 2584.120 18.030 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 817.490 17.580 817.810 17.640 ;
        RECT 820.710 17.580 821.030 17.640 ;
        RECT 817.490 17.440 821.030 17.580 ;
        RECT 817.490 17.380 817.810 17.440 ;
        RECT 820.710 17.380 821.030 17.440 ;
      LAYER via ;
        RECT 817.520 17.380 817.780 17.640 ;
        RECT 820.740 17.380 821.000 17.640 ;
      LAYER met2 ;
        RECT 820.800 17.670 820.940 54.000 ;
        RECT 817.520 17.350 817.780 17.670 ;
        RECT 820.740 17.350 821.000 17.670 ;
        RECT 817.580 2.400 817.720 17.350 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2435.310 18.940 2435.630 19.000 ;
        RECT 2572.390 18.940 2572.710 19.000 ;
        RECT 2435.310 18.800 2572.710 18.940 ;
        RECT 2435.310 18.740 2435.630 18.800 ;
        RECT 2572.390 18.740 2572.710 18.800 ;
        RECT 2572.390 16.220 2572.710 16.280 ;
        RECT 2601.370 16.220 2601.690 16.280 ;
        RECT 2572.390 16.080 2601.690 16.220 ;
        RECT 2572.390 16.020 2572.710 16.080 ;
        RECT 2601.370 16.020 2601.690 16.080 ;
      LAYER via ;
        RECT 2435.340 18.740 2435.600 19.000 ;
        RECT 2572.420 18.740 2572.680 19.000 ;
        RECT 2572.420 16.020 2572.680 16.280 ;
        RECT 2601.400 16.020 2601.660 16.280 ;
      LAYER met2 ;
        RECT 2435.400 19.030 2435.540 54.000 ;
        RECT 2435.340 18.710 2435.600 19.030 ;
        RECT 2572.420 18.710 2572.680 19.030 ;
        RECT 2572.480 16.310 2572.620 18.710 ;
        RECT 2572.420 15.990 2572.680 16.310 ;
        RECT 2601.400 15.990 2601.660 16.310 ;
        RECT 2601.460 2.400 2601.600 15.990 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2449.110 19.280 2449.430 19.340 ;
        RECT 2619.310 19.280 2619.630 19.340 ;
        RECT 2449.110 19.140 2619.630 19.280 ;
        RECT 2449.110 19.080 2449.430 19.140 ;
        RECT 2619.310 19.080 2619.630 19.140 ;
      LAYER via ;
        RECT 2449.140 19.080 2449.400 19.340 ;
        RECT 2619.340 19.080 2619.600 19.340 ;
      LAYER met2 ;
        RECT 2449.200 19.370 2449.340 54.000 ;
        RECT 2449.140 19.050 2449.400 19.370 ;
        RECT 2619.340 19.050 2619.600 19.370 ;
        RECT 2619.400 2.400 2619.540 19.050 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2462.910 17.240 2463.230 17.300 ;
        RECT 2637.250 17.240 2637.570 17.300 ;
        RECT 2462.910 17.100 2637.570 17.240 ;
        RECT 2462.910 17.040 2463.230 17.100 ;
        RECT 2637.250 17.040 2637.570 17.100 ;
      LAYER via ;
        RECT 2462.940 17.040 2463.200 17.300 ;
        RECT 2637.280 17.040 2637.540 17.300 ;
      LAYER met2 ;
        RECT 2463.000 17.330 2463.140 54.000 ;
        RECT 2462.940 17.010 2463.200 17.330 ;
        RECT 2637.280 17.010 2637.540 17.330 ;
        RECT 2637.340 2.400 2637.480 17.010 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2476.710 17.920 2477.030 17.980 ;
        RECT 2655.190 17.920 2655.510 17.980 ;
        RECT 2476.710 17.780 2655.510 17.920 ;
        RECT 2476.710 17.720 2477.030 17.780 ;
        RECT 2655.190 17.720 2655.510 17.780 ;
      LAYER via ;
        RECT 2476.740 17.720 2477.000 17.980 ;
        RECT 2655.220 17.720 2655.480 17.980 ;
      LAYER met2 ;
        RECT 2476.800 18.010 2476.940 54.000 ;
        RECT 2476.740 17.690 2477.000 18.010 ;
        RECT 2655.220 17.690 2655.480 18.010 ;
        RECT 2655.280 2.400 2655.420 17.690 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2497.410 15.880 2497.730 15.940 ;
        RECT 2672.670 15.880 2672.990 15.940 ;
        RECT 2497.410 15.740 2672.990 15.880 ;
        RECT 2497.410 15.680 2497.730 15.740 ;
        RECT 2672.670 15.680 2672.990 15.740 ;
      LAYER via ;
        RECT 2497.440 15.680 2497.700 15.940 ;
        RECT 2672.700 15.680 2672.960 15.940 ;
      LAYER met2 ;
        RECT 2497.500 15.970 2497.640 54.000 ;
        RECT 2497.440 15.650 2497.700 15.970 ;
        RECT 2672.700 15.650 2672.960 15.970 ;
        RECT 2672.760 2.400 2672.900 15.650 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2511.210 16.560 2511.530 16.620 ;
        RECT 2690.610 16.560 2690.930 16.620 ;
        RECT 2511.210 16.420 2690.930 16.560 ;
        RECT 2511.210 16.360 2511.530 16.420 ;
        RECT 2690.610 16.360 2690.930 16.420 ;
      LAYER via ;
        RECT 2511.240 16.360 2511.500 16.620 ;
        RECT 2690.640 16.360 2690.900 16.620 ;
      LAYER met2 ;
        RECT 2511.300 16.650 2511.440 54.000 ;
        RECT 2511.240 16.330 2511.500 16.650 ;
        RECT 2690.640 16.330 2690.900 16.650 ;
        RECT 2690.700 2.400 2690.840 16.330 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2525.010 18.600 2525.330 18.660 ;
        RECT 2708.550 18.600 2708.870 18.660 ;
        RECT 2525.010 18.460 2708.870 18.600 ;
        RECT 2525.010 18.400 2525.330 18.460 ;
        RECT 2708.550 18.400 2708.870 18.460 ;
      LAYER via ;
        RECT 2525.040 18.400 2525.300 18.660 ;
        RECT 2708.580 18.400 2708.840 18.660 ;
      LAYER met2 ;
        RECT 2525.100 18.690 2525.240 54.000 ;
        RECT 2525.040 18.370 2525.300 18.690 ;
        RECT 2708.580 18.370 2708.840 18.690 ;
        RECT 2708.640 2.400 2708.780 18.370 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2538.810 20.300 2539.130 20.360 ;
        RECT 2584.350 20.300 2584.670 20.360 ;
        RECT 2538.810 20.160 2584.670 20.300 ;
        RECT 2538.810 20.100 2539.130 20.160 ;
        RECT 2584.350 20.100 2584.670 20.160 ;
        RECT 2642.310 20.300 2642.630 20.360 ;
        RECT 2726.490 20.300 2726.810 20.360 ;
        RECT 2642.310 20.160 2726.810 20.300 ;
        RECT 2642.310 20.100 2642.630 20.160 ;
        RECT 2726.490 20.100 2726.810 20.160 ;
        RECT 2584.350 14.860 2584.670 14.920 ;
        RECT 2642.310 14.860 2642.630 14.920 ;
        RECT 2584.350 14.720 2642.630 14.860 ;
        RECT 2584.350 14.660 2584.670 14.720 ;
        RECT 2642.310 14.660 2642.630 14.720 ;
      LAYER via ;
        RECT 2538.840 20.100 2539.100 20.360 ;
        RECT 2584.380 20.100 2584.640 20.360 ;
        RECT 2642.340 20.100 2642.600 20.360 ;
        RECT 2726.520 20.100 2726.780 20.360 ;
        RECT 2584.380 14.660 2584.640 14.920 ;
        RECT 2642.340 14.660 2642.600 14.920 ;
      LAYER met2 ;
        RECT 2538.900 20.390 2539.040 54.000 ;
        RECT 2538.840 20.070 2539.100 20.390 ;
        RECT 2584.380 20.070 2584.640 20.390 ;
        RECT 2642.340 20.070 2642.600 20.390 ;
        RECT 2726.520 20.070 2726.780 20.390 ;
        RECT 2584.440 14.950 2584.580 20.070 ;
        RECT 2642.400 14.950 2642.540 20.070 ;
        RECT 2584.380 14.630 2584.640 14.950 ;
        RECT 2642.340 14.630 2642.600 14.950 ;
        RECT 2726.580 2.400 2726.720 20.070 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2552.610 19.960 2552.930 20.020 ;
        RECT 2574.230 19.960 2574.550 20.020 ;
        RECT 2552.610 19.820 2574.550 19.960 ;
        RECT 2552.610 19.760 2552.930 19.820 ;
        RECT 2574.230 19.760 2574.550 19.820 ;
        RECT 2641.850 19.960 2642.170 20.020 ;
        RECT 2714.990 19.960 2715.310 20.020 ;
        RECT 2641.850 19.820 2715.310 19.960 ;
        RECT 2641.850 19.760 2642.170 19.820 ;
        RECT 2714.990 19.760 2715.310 19.820 ;
        RECT 2714.990 18.600 2715.310 18.660 ;
        RECT 2744.430 18.600 2744.750 18.660 ;
        RECT 2714.990 18.460 2744.750 18.600 ;
        RECT 2714.990 18.400 2715.310 18.460 ;
        RECT 2744.430 18.400 2744.750 18.460 ;
        RECT 2574.230 14.520 2574.550 14.580 ;
        RECT 2641.850 14.520 2642.170 14.580 ;
        RECT 2574.230 14.380 2642.170 14.520 ;
        RECT 2574.230 14.320 2574.550 14.380 ;
        RECT 2641.850 14.320 2642.170 14.380 ;
      LAYER via ;
        RECT 2552.640 19.760 2552.900 20.020 ;
        RECT 2574.260 19.760 2574.520 20.020 ;
        RECT 2641.880 19.760 2642.140 20.020 ;
        RECT 2715.020 19.760 2715.280 20.020 ;
        RECT 2715.020 18.400 2715.280 18.660 ;
        RECT 2744.460 18.400 2744.720 18.660 ;
        RECT 2574.260 14.320 2574.520 14.580 ;
        RECT 2641.880 14.320 2642.140 14.580 ;
      LAYER met2 ;
        RECT 2552.700 20.050 2552.840 54.000 ;
        RECT 2552.640 19.730 2552.900 20.050 ;
        RECT 2574.260 19.730 2574.520 20.050 ;
        RECT 2641.880 19.730 2642.140 20.050 ;
        RECT 2715.020 19.730 2715.280 20.050 ;
        RECT 2574.320 14.610 2574.460 19.730 ;
        RECT 2641.940 14.610 2642.080 19.730 ;
        RECT 2715.080 18.690 2715.220 19.730 ;
        RECT 2715.020 18.370 2715.280 18.690 ;
        RECT 2744.460 18.370 2744.720 18.690 ;
        RECT 2574.260 14.290 2574.520 14.610 ;
        RECT 2641.880 14.290 2642.140 14.610 ;
        RECT 2744.520 2.400 2744.660 18.370 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2573.310 20.640 2573.630 20.700 ;
        RECT 2761.910 20.640 2762.230 20.700 ;
        RECT 2573.310 20.500 2762.230 20.640 ;
        RECT 2573.310 20.440 2573.630 20.500 ;
        RECT 2761.910 20.440 2762.230 20.500 ;
      LAYER via ;
        RECT 2573.340 20.440 2573.600 20.700 ;
        RECT 2761.940 20.440 2762.200 20.700 ;
      LAYER met2 ;
        RECT 2573.400 20.730 2573.540 54.000 ;
        RECT 2573.340 20.410 2573.600 20.730 ;
        RECT 2761.940 20.410 2762.200 20.730 ;
        RECT 2762.000 2.400 2762.140 20.410 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 835.430 17.920 835.750 17.980 ;
        RECT 840.950 17.920 841.270 17.980 ;
        RECT 835.430 17.780 841.270 17.920 ;
        RECT 835.430 17.720 835.750 17.780 ;
        RECT 840.950 17.720 841.270 17.780 ;
      LAYER via ;
        RECT 835.460 17.720 835.720 17.980 ;
        RECT 840.980 17.720 841.240 17.980 ;
      LAYER met2 ;
        RECT 841.040 18.010 841.180 54.000 ;
        RECT 835.460 17.690 835.720 18.010 ;
        RECT 840.980 17.690 841.240 18.010 ;
        RECT 835.520 2.400 835.660 17.690 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2597.230 18.260 2597.550 18.320 ;
        RECT 2601.830 18.260 2602.150 18.320 ;
        RECT 2597.230 18.120 2602.150 18.260 ;
        RECT 2597.230 18.060 2597.550 18.120 ;
        RECT 2601.830 18.060 2602.150 18.120 ;
        RECT 2601.830 16.220 2602.150 16.280 ;
        RECT 2779.850 16.220 2780.170 16.280 ;
        RECT 2601.830 16.080 2780.170 16.220 ;
        RECT 2601.830 16.020 2602.150 16.080 ;
        RECT 2779.850 16.020 2780.170 16.080 ;
      LAYER via ;
        RECT 2597.260 18.060 2597.520 18.320 ;
        RECT 2601.860 18.060 2602.120 18.320 ;
        RECT 2601.860 16.020 2602.120 16.280 ;
        RECT 2779.880 16.020 2780.140 16.280 ;
      LAYER met2 ;
        RECT 2597.780 52.770 2597.920 54.000 ;
        RECT 2597.320 52.630 2597.920 52.770 ;
        RECT 2597.320 18.350 2597.460 52.630 ;
        RECT 2597.260 18.030 2597.520 18.350 ;
        RECT 2601.860 18.030 2602.120 18.350 ;
        RECT 2601.920 16.310 2602.060 18.030 ;
        RECT 2601.860 15.990 2602.120 16.310 ;
        RECT 2779.880 15.990 2780.140 16.310 ;
        RECT 2779.940 2.400 2780.080 15.990 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2632.190 15.200 2632.510 15.260 ;
        RECT 2797.790 15.200 2798.110 15.260 ;
        RECT 2632.190 15.060 2798.110 15.200 ;
        RECT 2632.190 15.000 2632.510 15.060 ;
        RECT 2797.790 15.000 2798.110 15.060 ;
      LAYER via ;
        RECT 2632.220 15.000 2632.480 15.260 ;
        RECT 2797.820 15.000 2798.080 15.260 ;
      LAYER met2 ;
        RECT 2632.280 15.290 2632.420 54.000 ;
        RECT 2632.220 14.970 2632.480 15.290 ;
        RECT 2797.820 14.970 2798.080 15.290 ;
        RECT 2797.880 2.400 2798.020 14.970 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2614.710 18.260 2615.030 18.320 ;
        RECT 2815.730 18.260 2816.050 18.320 ;
        RECT 2614.710 18.120 2816.050 18.260 ;
        RECT 2614.710 18.060 2615.030 18.120 ;
        RECT 2815.730 18.060 2816.050 18.120 ;
      LAYER via ;
        RECT 2614.740 18.060 2615.000 18.320 ;
        RECT 2815.760 18.060 2816.020 18.320 ;
      LAYER met2 ;
        RECT 2614.800 18.350 2614.940 54.000 ;
        RECT 2614.740 18.030 2615.000 18.350 ;
        RECT 2815.760 18.030 2816.020 18.350 ;
        RECT 2815.820 2.400 2815.960 18.030 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2673.590 15.540 2673.910 15.600 ;
        RECT 2833.670 15.540 2833.990 15.600 ;
        RECT 2673.590 15.400 2833.990 15.540 ;
        RECT 2673.590 15.340 2673.910 15.400 ;
        RECT 2833.670 15.340 2833.990 15.400 ;
      LAYER via ;
        RECT 2673.620 15.340 2673.880 15.600 ;
        RECT 2833.700 15.340 2833.960 15.600 ;
      LAYER met2 ;
        RECT 2673.680 15.630 2673.820 54.000 ;
        RECT 2673.620 15.310 2673.880 15.630 ;
        RECT 2833.700 15.310 2833.960 15.630 ;
        RECT 2833.760 2.400 2833.900 15.310 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2687.390 15.880 2687.710 15.940 ;
        RECT 2851.150 15.880 2851.470 15.940 ;
        RECT 2687.390 15.740 2851.470 15.880 ;
        RECT 2687.390 15.680 2687.710 15.740 ;
        RECT 2851.150 15.680 2851.470 15.740 ;
      LAYER via ;
        RECT 2687.420 15.680 2687.680 15.940 ;
        RECT 2851.180 15.680 2851.440 15.940 ;
      LAYER met2 ;
        RECT 2687.480 15.970 2687.620 54.000 ;
        RECT 2687.420 15.650 2687.680 15.970 ;
        RECT 2851.180 15.650 2851.440 15.970 ;
        RECT 2851.240 2.400 2851.380 15.650 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2663.010 17.920 2663.330 17.980 ;
        RECT 2869.090 17.920 2869.410 17.980 ;
        RECT 2663.010 17.780 2869.410 17.920 ;
        RECT 2663.010 17.720 2663.330 17.780 ;
        RECT 2869.090 17.720 2869.410 17.780 ;
      LAYER via ;
        RECT 2663.040 17.720 2663.300 17.980 ;
        RECT 2869.120 17.720 2869.380 17.980 ;
      LAYER met2 ;
        RECT 2663.100 18.010 2663.240 54.000 ;
        RECT 2663.040 17.690 2663.300 18.010 ;
        RECT 2869.120 17.690 2869.380 18.010 ;
        RECT 2869.180 2.400 2869.320 17.690 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2732.930 16.560 2733.250 16.620 ;
        RECT 2887.030 16.560 2887.350 16.620 ;
        RECT 2732.930 16.420 2887.350 16.560 ;
        RECT 2732.930 16.360 2733.250 16.420 ;
        RECT 2887.030 16.360 2887.350 16.420 ;
        RECT 2701.190 14.860 2701.510 14.920 ;
        RECT 2732.930 14.860 2733.250 14.920 ;
        RECT 2701.190 14.720 2733.250 14.860 ;
        RECT 2701.190 14.660 2701.510 14.720 ;
        RECT 2732.930 14.660 2733.250 14.720 ;
      LAYER via ;
        RECT 2732.960 16.360 2733.220 16.620 ;
        RECT 2887.060 16.360 2887.320 16.620 ;
        RECT 2701.220 14.660 2701.480 14.920 ;
        RECT 2732.960 14.660 2733.220 14.920 ;
      LAYER met2 ;
        RECT 2701.280 14.950 2701.420 54.000 ;
        RECT 2732.960 16.330 2733.220 16.650 ;
        RECT 2887.060 16.330 2887.320 16.650 ;
        RECT 2733.020 14.950 2733.160 16.330 ;
        RECT 2701.220 14.630 2701.480 14.950 ;
        RECT 2732.960 14.630 2733.220 14.950 ;
        RECT 2887.120 2.400 2887.260 16.330 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2763.290 18.600 2763.610 18.660 ;
        RECT 2904.970 18.600 2905.290 18.660 ;
        RECT 2763.290 18.460 2905.290 18.600 ;
        RECT 2763.290 18.400 2763.610 18.460 ;
        RECT 2904.970 18.400 2905.290 18.460 ;
        RECT 2763.290 14.860 2763.610 14.920 ;
        RECT 2733.480 14.720 2763.610 14.860 ;
        RECT 2708.090 14.520 2708.410 14.580 ;
        RECT 2733.480 14.520 2733.620 14.720 ;
        RECT 2763.290 14.660 2763.610 14.720 ;
        RECT 2708.090 14.380 2733.620 14.520 ;
        RECT 2708.090 14.320 2708.410 14.380 ;
      LAYER via ;
        RECT 2763.320 18.400 2763.580 18.660 ;
        RECT 2905.000 18.400 2905.260 18.660 ;
        RECT 2708.120 14.320 2708.380 14.580 ;
        RECT 2763.320 14.660 2763.580 14.920 ;
      LAYER met2 ;
        RECT 2708.180 14.610 2708.320 54.000 ;
        RECT 2763.320 18.370 2763.580 18.690 ;
        RECT 2905.000 18.370 2905.260 18.690 ;
        RECT 2763.380 14.950 2763.520 18.370 ;
        RECT 2763.320 14.630 2763.580 14.950 ;
        RECT 2708.120 14.290 2708.380 14.610 ;
        RECT 2905.060 2.400 2905.200 18.370 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 852.910 16.900 853.230 16.960 ;
        RECT 855.210 16.900 855.530 16.960 ;
        RECT 852.910 16.760 855.530 16.900 ;
        RECT 852.910 16.700 853.230 16.760 ;
        RECT 855.210 16.700 855.530 16.760 ;
      LAYER via ;
        RECT 852.940 16.700 853.200 16.960 ;
        RECT 855.240 16.700 855.500 16.960 ;
      LAYER met2 ;
        RECT 855.300 16.990 855.440 54.000 ;
        RECT 852.940 16.670 853.200 16.990 ;
        RECT 855.240 16.670 855.500 16.990 ;
        RECT 853.000 2.400 853.140 16.670 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 870.850 16.560 871.170 16.620 ;
        RECT 875.910 16.560 876.230 16.620 ;
        RECT 870.850 16.420 876.230 16.560 ;
        RECT 870.850 16.360 871.170 16.420 ;
        RECT 875.910 16.360 876.230 16.420 ;
      LAYER via ;
        RECT 870.880 16.360 871.140 16.620 ;
        RECT 875.940 16.360 876.200 16.620 ;
      LAYER met2 ;
        RECT 876.000 16.650 876.140 54.000 ;
        RECT 870.880 16.330 871.140 16.650 ;
        RECT 875.940 16.330 876.200 16.650 ;
        RECT 870.940 2.400 871.080 16.330 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 889.800 17.410 889.940 54.000 ;
        RECT 888.880 17.270 889.940 17.410 ;
        RECT 888.880 2.400 889.020 17.270 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 906.730 15.540 907.050 15.600 ;
        RECT 910.410 15.540 910.730 15.600 ;
        RECT 906.730 15.400 910.730 15.540 ;
        RECT 906.730 15.340 907.050 15.400 ;
        RECT 910.410 15.340 910.730 15.400 ;
      LAYER via ;
        RECT 906.760 15.340 907.020 15.600 ;
        RECT 910.440 15.340 910.700 15.600 ;
      LAYER met2 ;
        RECT 910.500 15.630 910.640 54.000 ;
        RECT 906.760 15.310 907.020 15.630 ;
        RECT 910.440 15.310 910.700 15.630 ;
        RECT 906.820 2.400 906.960 15.310 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.300 2.400 924.440 54.000 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 942.150 17.580 942.470 17.640 ;
        RECT 944.910 17.580 945.230 17.640 ;
        RECT 942.150 17.440 945.230 17.580 ;
        RECT 942.150 17.380 942.470 17.440 ;
        RECT 944.910 17.380 945.230 17.440 ;
      LAYER via ;
        RECT 942.180 17.380 942.440 17.640 ;
        RECT 944.940 17.380 945.200 17.640 ;
      LAYER met2 ;
        RECT 945.000 17.670 945.140 54.000 ;
        RECT 942.180 17.350 942.440 17.670 ;
        RECT 944.940 17.350 945.200 17.670 ;
        RECT 942.240 2.400 942.380 17.350 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 960.090 17.580 960.410 17.640 ;
        RECT 965.610 17.580 965.930 17.640 ;
        RECT 960.090 17.440 965.930 17.580 ;
        RECT 960.090 17.380 960.410 17.440 ;
        RECT 965.610 17.380 965.930 17.440 ;
      LAYER via ;
        RECT 960.120 17.380 960.380 17.640 ;
        RECT 965.640 17.380 965.900 17.640 ;
      LAYER met2 ;
        RECT 965.700 17.670 965.840 54.000 ;
        RECT 960.120 17.350 960.380 17.670 ;
        RECT 965.640 17.350 965.900 17.670 ;
        RECT 960.180 2.400 960.320 17.350 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 979.500 17.410 979.640 54.000 ;
        RECT 978.120 17.270 979.640 17.410 ;
        RECT 978.120 2.400 978.260 17.270 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 16.900 657.270 16.960 ;
        RECT 662.010 16.900 662.330 16.960 ;
        RECT 656.950 16.760 662.330 16.900 ;
        RECT 656.950 16.700 657.270 16.760 ;
        RECT 662.010 16.700 662.330 16.760 ;
      LAYER via ;
        RECT 656.980 16.700 657.240 16.960 ;
        RECT 662.040 16.700 662.300 16.960 ;
      LAYER met2 ;
        RECT 662.100 16.990 662.240 54.000 ;
        RECT 656.980 16.670 657.240 16.990 ;
        RECT 662.040 16.670 662.300 16.990 ;
        RECT 657.040 2.400 657.180 16.670 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 995.970 17.580 996.290 17.640 ;
        RECT 1000.110 17.580 1000.430 17.640 ;
        RECT 995.970 17.440 1000.430 17.580 ;
        RECT 995.970 17.380 996.290 17.440 ;
        RECT 1000.110 17.380 1000.430 17.440 ;
      LAYER via ;
        RECT 996.000 17.380 996.260 17.640 ;
        RECT 1000.140 17.380 1000.400 17.640 ;
      LAYER met2 ;
        RECT 1000.200 17.670 1000.340 54.000 ;
        RECT 996.000 17.350 996.260 17.670 ;
        RECT 1000.140 17.350 1000.400 17.670 ;
        RECT 996.060 2.400 996.200 17.350 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1014.000 17.410 1014.140 54.000 ;
        RECT 1013.540 17.270 1014.140 17.410 ;
        RECT 1013.540 2.400 1013.680 17.270 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1031.390 15.200 1031.710 15.260 ;
        RECT 1034.610 15.200 1034.930 15.260 ;
        RECT 1031.390 15.060 1034.930 15.200 ;
        RECT 1031.390 15.000 1031.710 15.060 ;
        RECT 1034.610 15.000 1034.930 15.060 ;
      LAYER via ;
        RECT 1031.420 15.000 1031.680 15.260 ;
        RECT 1034.640 15.000 1034.900 15.260 ;
      LAYER met2 ;
        RECT 1034.700 15.290 1034.840 54.000 ;
        RECT 1031.420 14.970 1031.680 15.290 ;
        RECT 1034.640 14.970 1034.900 15.290 ;
        RECT 1031.480 2.400 1031.620 14.970 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1049.330 17.580 1049.650 17.640 ;
        RECT 1055.310 17.580 1055.630 17.640 ;
        RECT 1049.330 17.440 1055.630 17.580 ;
        RECT 1049.330 17.380 1049.650 17.440 ;
        RECT 1055.310 17.380 1055.630 17.440 ;
      LAYER via ;
        RECT 1049.360 17.380 1049.620 17.640 ;
        RECT 1055.340 17.380 1055.600 17.640 ;
      LAYER met2 ;
        RECT 1055.400 17.670 1055.540 54.000 ;
        RECT 1049.360 17.350 1049.620 17.670 ;
        RECT 1055.340 17.350 1055.600 17.670 ;
        RECT 1049.420 2.400 1049.560 17.350 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1069.200 17.410 1069.340 54.000 ;
        RECT 1067.360 17.270 1069.340 17.410 ;
        RECT 1067.360 2.400 1067.500 17.270 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1085.210 17.580 1085.530 17.640 ;
        RECT 1089.810 17.580 1090.130 17.640 ;
        RECT 1085.210 17.440 1090.130 17.580 ;
        RECT 1085.210 17.380 1085.530 17.440 ;
        RECT 1089.810 17.380 1090.130 17.440 ;
      LAYER via ;
        RECT 1085.240 17.380 1085.500 17.640 ;
        RECT 1089.840 17.380 1090.100 17.640 ;
      LAYER met2 ;
        RECT 1089.900 17.670 1090.040 54.000 ;
        RECT 1085.240 17.350 1085.500 17.670 ;
        RECT 1089.840 17.350 1090.100 17.670 ;
        RECT 1085.300 2.400 1085.440 17.350 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1103.700 17.410 1103.840 54.000 ;
        RECT 1102.780 17.270 1103.840 17.410 ;
        RECT 1102.780 2.400 1102.920 17.270 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1120.630 17.580 1120.950 17.640 ;
        RECT 1124.310 17.580 1124.630 17.640 ;
        RECT 1120.630 17.440 1124.630 17.580 ;
        RECT 1120.630 17.380 1120.950 17.440 ;
        RECT 1124.310 17.380 1124.630 17.440 ;
      LAYER via ;
        RECT 1120.660 17.380 1120.920 17.640 ;
        RECT 1124.340 17.380 1124.600 17.640 ;
      LAYER met2 ;
        RECT 1124.400 17.670 1124.540 54.000 ;
        RECT 1120.660 17.350 1120.920 17.670 ;
        RECT 1124.340 17.350 1124.600 17.670 ;
        RECT 1120.720 2.400 1120.860 17.350 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1138.570 17.920 1138.890 17.980 ;
        RECT 1144.550 17.920 1144.870 17.980 ;
        RECT 1138.570 17.780 1144.870 17.920 ;
        RECT 1138.570 17.720 1138.890 17.780 ;
        RECT 1144.550 17.720 1144.870 17.780 ;
      LAYER via ;
        RECT 1138.600 17.720 1138.860 17.980 ;
        RECT 1144.580 17.720 1144.840 17.980 ;
      LAYER met2 ;
        RECT 1144.640 18.010 1144.780 54.000 ;
        RECT 1138.600 17.690 1138.860 18.010 ;
        RECT 1144.580 17.690 1144.840 18.010 ;
        RECT 1138.660 2.400 1138.800 17.690 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1156.510 17.580 1156.830 17.640 ;
        RECT 1158.810 17.580 1159.130 17.640 ;
        RECT 1156.510 17.440 1159.130 17.580 ;
        RECT 1156.510 17.380 1156.830 17.440 ;
        RECT 1158.810 17.380 1159.130 17.440 ;
      LAYER via ;
        RECT 1156.540 17.380 1156.800 17.640 ;
        RECT 1158.840 17.380 1159.100 17.640 ;
      LAYER met2 ;
        RECT 1158.900 17.670 1159.040 54.000 ;
        RECT 1156.540 17.350 1156.800 17.670 ;
        RECT 1158.840 17.350 1159.100 17.670 ;
        RECT 1156.600 2.400 1156.740 17.350 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 675.900 17.410 676.040 54.000 ;
        RECT 674.520 17.270 676.040 17.410 ;
        RECT 674.520 2.400 674.660 17.270 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1173.990 16.560 1174.310 16.620 ;
        RECT 1179.510 16.560 1179.830 16.620 ;
        RECT 1173.990 16.420 1179.830 16.560 ;
        RECT 1173.990 16.360 1174.310 16.420 ;
        RECT 1179.510 16.360 1179.830 16.420 ;
      LAYER via ;
        RECT 1174.020 16.360 1174.280 16.620 ;
        RECT 1179.540 16.360 1179.800 16.620 ;
      LAYER met2 ;
        RECT 1179.600 16.650 1179.740 54.000 ;
        RECT 1174.020 16.330 1174.280 16.650 ;
        RECT 1179.540 16.330 1179.800 16.650 ;
        RECT 1174.080 2.400 1174.220 16.330 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1193.400 17.410 1193.540 54.000 ;
        RECT 1192.020 17.270 1193.540 17.410 ;
        RECT 1192.020 2.400 1192.160 17.270 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1209.870 17.240 1210.190 17.300 ;
        RECT 1214.010 17.240 1214.330 17.300 ;
        RECT 1209.870 17.100 1214.330 17.240 ;
        RECT 1209.870 17.040 1210.190 17.100 ;
        RECT 1214.010 17.040 1214.330 17.100 ;
      LAYER via ;
        RECT 1209.900 17.040 1210.160 17.300 ;
        RECT 1214.040 17.040 1214.300 17.300 ;
      LAYER met2 ;
        RECT 1214.100 17.330 1214.240 54.000 ;
        RECT 1209.900 17.010 1210.160 17.330 ;
        RECT 1214.040 17.010 1214.300 17.330 ;
        RECT 1209.960 2.400 1210.100 17.010 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.440 17.410 1227.580 54.000 ;
        RECT 1227.440 17.270 1228.040 17.410 ;
        RECT 1227.900 2.400 1228.040 17.270 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1245.750 17.580 1246.070 17.640 ;
        RECT 1248.510 17.580 1248.830 17.640 ;
        RECT 1245.750 17.440 1248.830 17.580 ;
        RECT 1245.750 17.380 1246.070 17.440 ;
        RECT 1248.510 17.380 1248.830 17.440 ;
      LAYER via ;
        RECT 1245.780 17.380 1246.040 17.640 ;
        RECT 1248.540 17.380 1248.800 17.640 ;
      LAYER met2 ;
        RECT 1248.600 17.670 1248.740 54.000 ;
        RECT 1245.780 17.350 1246.040 17.670 ;
        RECT 1248.540 17.350 1248.800 17.670 ;
        RECT 1245.840 2.400 1245.980 17.350 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1263.230 17.920 1263.550 17.980 ;
        RECT 1269.210 17.920 1269.530 17.980 ;
        RECT 1263.230 17.780 1269.530 17.920 ;
        RECT 1263.230 17.720 1263.550 17.780 ;
        RECT 1269.210 17.720 1269.530 17.780 ;
      LAYER via ;
        RECT 1263.260 17.720 1263.520 17.980 ;
        RECT 1269.240 17.720 1269.500 17.980 ;
      LAYER met2 ;
        RECT 1269.300 18.010 1269.440 54.000 ;
        RECT 1263.260 17.690 1263.520 18.010 ;
        RECT 1269.240 17.690 1269.500 18.010 ;
        RECT 1263.320 2.400 1263.460 17.690 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1283.100 17.410 1283.240 54.000 ;
        RECT 1281.260 17.270 1283.240 17.410 ;
        RECT 1281.260 2.400 1281.400 17.270 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1299.110 15.200 1299.430 15.260 ;
        RECT 1303.710 15.200 1304.030 15.260 ;
        RECT 1299.110 15.060 1304.030 15.200 ;
        RECT 1299.110 15.000 1299.430 15.060 ;
        RECT 1303.710 15.000 1304.030 15.060 ;
      LAYER via ;
        RECT 1299.140 15.000 1299.400 15.260 ;
        RECT 1303.740 15.000 1304.000 15.260 ;
      LAYER met2 ;
        RECT 1303.800 15.290 1303.940 54.000 ;
        RECT 1299.140 14.970 1299.400 15.290 ;
        RECT 1303.740 14.970 1304.000 15.290 ;
        RECT 1299.200 2.400 1299.340 14.970 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1317.600 17.410 1317.740 54.000 ;
        RECT 1317.140 17.270 1317.740 17.410 ;
        RECT 1317.140 2.400 1317.280 17.270 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1334.990 16.220 1335.310 16.280 ;
        RECT 1339.130 16.220 1339.450 16.280 ;
        RECT 1334.990 16.080 1339.450 16.220 ;
        RECT 1334.990 16.020 1335.310 16.080 ;
        RECT 1339.130 16.020 1339.450 16.080 ;
      LAYER via ;
        RECT 1335.020 16.020 1335.280 16.280 ;
        RECT 1339.160 16.020 1339.420 16.280 ;
      LAYER met2 ;
        RECT 1339.220 16.310 1339.360 54.000 ;
        RECT 1335.020 15.990 1335.280 16.310 ;
        RECT 1339.160 15.990 1339.420 16.310 ;
        RECT 1335.080 2.400 1335.220 15.990 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 692.370 17.240 692.690 17.300 ;
        RECT 696.510 17.240 696.830 17.300 ;
        RECT 692.370 17.100 696.830 17.240 ;
        RECT 692.370 17.040 692.690 17.100 ;
        RECT 696.510 17.040 696.830 17.100 ;
      LAYER via ;
        RECT 692.400 17.040 692.660 17.300 ;
        RECT 696.540 17.040 696.800 17.300 ;
      LAYER met2 ;
        RECT 696.600 17.330 696.740 54.000 ;
        RECT 692.400 17.010 692.660 17.330 ;
        RECT 696.540 17.010 696.800 17.330 ;
        RECT 692.460 2.400 692.600 17.010 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1353.480 17.410 1353.620 54.000 ;
        RECT 1352.560 17.270 1353.620 17.410 ;
        RECT 1352.560 2.400 1352.700 17.270 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1370.410 14.520 1370.730 14.580 ;
        RECT 1372.710 14.520 1373.030 14.580 ;
        RECT 1370.410 14.380 1373.030 14.520 ;
        RECT 1370.410 14.320 1370.730 14.380 ;
        RECT 1372.710 14.320 1373.030 14.380 ;
      LAYER via ;
        RECT 1370.440 14.320 1370.700 14.580 ;
        RECT 1372.740 14.320 1373.000 14.580 ;
      LAYER met2 ;
        RECT 1372.800 14.610 1372.940 54.000 ;
        RECT 1370.440 14.290 1370.700 14.610 ;
        RECT 1372.740 14.290 1373.000 14.610 ;
        RECT 1370.500 2.400 1370.640 14.290 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1387.060 17.410 1387.200 54.000 ;
        RECT 1387.060 17.270 1388.580 17.410 ;
        RECT 1388.440 2.400 1388.580 17.270 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1400.770 16.560 1401.090 16.620 ;
        RECT 1406.290 16.560 1406.610 16.620 ;
        RECT 1400.770 16.420 1406.610 16.560 ;
        RECT 1400.770 16.360 1401.090 16.420 ;
        RECT 1406.290 16.360 1406.610 16.420 ;
      LAYER via ;
        RECT 1400.800 16.360 1401.060 16.620 ;
        RECT 1406.320 16.360 1406.580 16.620 ;
      LAYER met2 ;
        RECT 1400.860 16.650 1401.000 54.000 ;
        RECT 1400.800 16.330 1401.060 16.650 ;
        RECT 1406.320 16.330 1406.580 16.650 ;
        RECT 1406.380 2.400 1406.520 16.330 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1422.020 17.410 1422.160 54.000 ;
        RECT 1422.020 17.270 1424.000 17.410 ;
        RECT 1423.860 2.400 1424.000 17.270 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1436.280 17.410 1436.420 54.000 ;
        RECT 1436.280 17.270 1441.940 17.410 ;
        RECT 1441.800 2.400 1441.940 17.270 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1455.510 17.580 1455.830 17.640 ;
        RECT 1459.650 17.580 1459.970 17.640 ;
        RECT 1455.510 17.440 1459.970 17.580 ;
        RECT 1455.510 17.380 1455.830 17.440 ;
        RECT 1459.650 17.380 1459.970 17.440 ;
      LAYER via ;
        RECT 1455.540 17.380 1455.800 17.640 ;
        RECT 1459.680 17.380 1459.940 17.640 ;
      LAYER met2 ;
        RECT 1455.600 17.670 1455.740 54.000 ;
        RECT 1455.540 17.350 1455.800 17.670 ;
        RECT 1459.680 17.350 1459.940 17.670 ;
        RECT 1459.740 2.400 1459.880 17.350 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1469.310 17.920 1469.630 17.980 ;
        RECT 1477.590 17.920 1477.910 17.980 ;
        RECT 1469.310 17.780 1477.910 17.920 ;
        RECT 1469.310 17.720 1469.630 17.780 ;
        RECT 1477.590 17.720 1477.910 17.780 ;
      LAYER via ;
        RECT 1469.340 17.720 1469.600 17.980 ;
        RECT 1477.620 17.720 1477.880 17.980 ;
      LAYER met2 ;
        RECT 1469.400 18.010 1469.540 54.000 ;
        RECT 1469.340 17.690 1469.600 18.010 ;
        RECT 1477.620 17.690 1477.880 18.010 ;
        RECT 1477.680 2.400 1477.820 17.690 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1483.110 20.640 1483.430 20.700 ;
        RECT 1495.530 20.640 1495.850 20.700 ;
        RECT 1483.110 20.500 1495.850 20.640 ;
        RECT 1483.110 20.440 1483.430 20.500 ;
        RECT 1495.530 20.440 1495.850 20.500 ;
      LAYER via ;
        RECT 1483.140 20.440 1483.400 20.700 ;
        RECT 1495.560 20.440 1495.820 20.700 ;
      LAYER met2 ;
        RECT 1483.200 20.730 1483.340 54.000 ;
        RECT 1483.140 20.410 1483.400 20.730 ;
        RECT 1495.560 20.410 1495.820 20.730 ;
        RECT 1495.620 2.400 1495.760 20.410 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1496.450 14.860 1496.770 14.920 ;
        RECT 1513.010 14.860 1513.330 14.920 ;
        RECT 1496.450 14.720 1513.330 14.860 ;
        RECT 1496.450 14.660 1496.770 14.720 ;
        RECT 1513.010 14.660 1513.330 14.720 ;
      LAYER via ;
        RECT 1496.480 14.660 1496.740 14.920 ;
        RECT 1513.040 14.660 1513.300 14.920 ;
      LAYER met2 ;
        RECT 1496.540 14.950 1496.680 54.000 ;
        RECT 1496.480 14.630 1496.740 14.950 ;
        RECT 1513.040 14.630 1513.300 14.950 ;
        RECT 1513.100 2.400 1513.240 14.630 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 709.940 7.890 710.080 54.000 ;
        RECT 709.940 7.750 710.540 7.890 ;
        RECT 710.400 2.400 710.540 7.750 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1517.610 15.880 1517.930 15.940 ;
        RECT 1530.950 15.880 1531.270 15.940 ;
        RECT 1517.610 15.740 1531.270 15.880 ;
        RECT 1517.610 15.680 1517.930 15.740 ;
        RECT 1530.950 15.680 1531.270 15.740 ;
      LAYER via ;
        RECT 1517.640 15.680 1517.900 15.940 ;
        RECT 1530.980 15.680 1531.240 15.940 ;
      LAYER met2 ;
        RECT 1517.700 15.970 1517.840 54.000 ;
        RECT 1517.640 15.650 1517.900 15.970 ;
        RECT 1530.980 15.650 1531.240 15.970 ;
        RECT 1531.040 2.400 1531.180 15.650 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1531.410 18.600 1531.730 18.660 ;
        RECT 1548.890 18.600 1549.210 18.660 ;
        RECT 1531.410 18.460 1549.210 18.600 ;
        RECT 1531.410 18.400 1531.730 18.460 ;
        RECT 1548.890 18.400 1549.210 18.460 ;
      LAYER via ;
        RECT 1531.440 18.400 1531.700 18.660 ;
        RECT 1548.920 18.400 1549.180 18.660 ;
      LAYER met2 ;
        RECT 1531.500 18.690 1531.640 54.000 ;
        RECT 1531.440 18.370 1531.700 18.690 ;
        RECT 1548.920 18.370 1549.180 18.690 ;
        RECT 1548.980 2.400 1549.120 18.370 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1545.210 17.580 1545.530 17.640 ;
        RECT 1566.830 17.580 1567.150 17.640 ;
        RECT 1545.210 17.440 1567.150 17.580 ;
        RECT 1545.210 17.380 1545.530 17.440 ;
        RECT 1566.830 17.380 1567.150 17.440 ;
      LAYER via ;
        RECT 1545.240 17.380 1545.500 17.640 ;
        RECT 1566.860 17.380 1567.120 17.640 ;
      LAYER met2 ;
        RECT 1545.300 17.670 1545.440 54.000 ;
        RECT 1545.240 17.350 1545.500 17.670 ;
        RECT 1566.860 17.350 1567.120 17.670 ;
        RECT 1566.920 2.400 1567.060 17.350 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1559.010 15.200 1559.330 15.260 ;
        RECT 1584.770 15.200 1585.090 15.260 ;
        RECT 1559.010 15.060 1585.090 15.200 ;
        RECT 1559.010 15.000 1559.330 15.060 ;
        RECT 1584.770 15.000 1585.090 15.060 ;
      LAYER via ;
        RECT 1559.040 15.000 1559.300 15.260 ;
        RECT 1584.800 15.000 1585.060 15.260 ;
      LAYER met2 ;
        RECT 1559.100 15.290 1559.240 54.000 ;
        RECT 1559.040 14.970 1559.300 15.290 ;
        RECT 1584.800 14.970 1585.060 15.290 ;
        RECT 1584.860 2.400 1585.000 14.970 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1572.810 17.920 1573.130 17.980 ;
        RECT 1602.250 17.920 1602.570 17.980 ;
        RECT 1572.810 17.780 1602.570 17.920 ;
        RECT 1572.810 17.720 1573.130 17.780 ;
        RECT 1602.250 17.720 1602.570 17.780 ;
      LAYER via ;
        RECT 1572.840 17.720 1573.100 17.980 ;
        RECT 1602.280 17.720 1602.540 17.980 ;
      LAYER met2 ;
        RECT 1572.900 18.010 1573.040 54.000 ;
        RECT 1572.840 17.690 1573.100 18.010 ;
        RECT 1602.280 17.690 1602.540 18.010 ;
        RECT 1602.340 2.400 1602.480 17.690 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1593.510 14.520 1593.830 14.580 ;
        RECT 1620.190 14.520 1620.510 14.580 ;
        RECT 1593.510 14.380 1620.510 14.520 ;
        RECT 1593.510 14.320 1593.830 14.380 ;
        RECT 1620.190 14.320 1620.510 14.380 ;
      LAYER via ;
        RECT 1593.540 14.320 1593.800 14.580 ;
        RECT 1620.220 14.320 1620.480 14.580 ;
      LAYER met2 ;
        RECT 1593.600 14.610 1593.740 54.000 ;
        RECT 1593.540 14.290 1593.800 14.610 ;
        RECT 1620.220 14.290 1620.480 14.610 ;
        RECT 1620.280 2.400 1620.420 14.290 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1607.310 15.200 1607.630 15.260 ;
        RECT 1638.130 15.200 1638.450 15.260 ;
        RECT 1607.310 15.060 1638.450 15.200 ;
        RECT 1607.310 15.000 1607.630 15.060 ;
        RECT 1638.130 15.000 1638.450 15.060 ;
      LAYER via ;
        RECT 1607.340 15.000 1607.600 15.260 ;
        RECT 1638.160 15.000 1638.420 15.260 ;
      LAYER met2 ;
        RECT 1607.400 15.290 1607.540 54.000 ;
        RECT 1607.340 14.970 1607.600 15.290 ;
        RECT 1638.160 14.970 1638.420 15.290 ;
        RECT 1638.220 2.400 1638.360 14.970 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1621.110 17.920 1621.430 17.980 ;
        RECT 1656.070 17.920 1656.390 17.980 ;
        RECT 1621.110 17.780 1656.390 17.920 ;
        RECT 1621.110 17.720 1621.430 17.780 ;
        RECT 1656.070 17.720 1656.390 17.780 ;
      LAYER via ;
        RECT 1621.140 17.720 1621.400 17.980 ;
        RECT 1656.100 17.720 1656.360 17.980 ;
      LAYER met2 ;
        RECT 1621.200 18.010 1621.340 54.000 ;
        RECT 1621.140 17.690 1621.400 18.010 ;
        RECT 1656.100 17.690 1656.360 18.010 ;
        RECT 1656.160 2.400 1656.300 17.690 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1634.910 14.520 1635.230 14.580 ;
        RECT 1673.550 14.520 1673.870 14.580 ;
        RECT 1634.910 14.380 1673.870 14.520 ;
        RECT 1634.910 14.320 1635.230 14.380 ;
        RECT 1673.550 14.320 1673.870 14.380 ;
      LAYER via ;
        RECT 1634.940 14.320 1635.200 14.580 ;
        RECT 1673.580 14.320 1673.840 14.580 ;
      LAYER met2 ;
        RECT 1635.000 14.610 1635.140 54.000 ;
        RECT 1634.940 14.290 1635.200 14.610 ;
        RECT 1673.580 14.290 1673.840 14.610 ;
        RECT 1673.640 2.400 1673.780 14.290 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1655.610 18.260 1655.930 18.320 ;
        RECT 1691.490 18.260 1691.810 18.320 ;
        RECT 1655.610 18.120 1691.810 18.260 ;
        RECT 1655.610 18.060 1655.930 18.120 ;
        RECT 1691.490 18.060 1691.810 18.120 ;
      LAYER via ;
        RECT 1655.640 18.060 1655.900 18.320 ;
        RECT 1691.520 18.060 1691.780 18.320 ;
      LAYER met2 ;
        RECT 1655.700 18.350 1655.840 54.000 ;
        RECT 1655.640 18.030 1655.900 18.350 ;
        RECT 1691.520 18.030 1691.780 18.350 ;
        RECT 1691.580 2.400 1691.720 18.030 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 728.250 17.580 728.570 17.640 ;
        RECT 731.010 17.580 731.330 17.640 ;
        RECT 728.250 17.440 731.330 17.580 ;
        RECT 728.250 17.380 728.570 17.440 ;
        RECT 731.010 17.380 731.330 17.440 ;
      LAYER via ;
        RECT 728.280 17.380 728.540 17.640 ;
        RECT 731.040 17.380 731.300 17.640 ;
      LAYER met2 ;
        RECT 731.100 17.670 731.240 54.000 ;
        RECT 728.280 17.350 728.540 17.670 ;
        RECT 731.040 17.350 731.300 17.670 ;
        RECT 728.340 2.400 728.480 17.350 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1669.410 19.280 1669.730 19.340 ;
        RECT 1709.430 19.280 1709.750 19.340 ;
        RECT 1669.410 19.140 1709.750 19.280 ;
        RECT 1669.410 19.080 1669.730 19.140 ;
        RECT 1709.430 19.080 1709.750 19.140 ;
      LAYER via ;
        RECT 1669.440 19.080 1669.700 19.340 ;
        RECT 1709.460 19.080 1709.720 19.340 ;
      LAYER met2 ;
        RECT 1669.500 19.370 1669.640 54.000 ;
        RECT 1669.440 19.050 1669.700 19.370 ;
        RECT 1709.460 19.050 1709.720 19.370 ;
        RECT 1709.520 2.400 1709.660 19.050 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1683.210 18.940 1683.530 19.000 ;
        RECT 1727.370 18.940 1727.690 19.000 ;
        RECT 1683.210 18.800 1727.690 18.940 ;
        RECT 1683.210 18.740 1683.530 18.800 ;
        RECT 1727.370 18.740 1727.690 18.800 ;
      LAYER via ;
        RECT 1683.240 18.740 1683.500 19.000 ;
        RECT 1727.400 18.740 1727.660 19.000 ;
      LAYER met2 ;
        RECT 1683.300 19.030 1683.440 54.000 ;
        RECT 1683.240 18.710 1683.500 19.030 ;
        RECT 1727.400 18.710 1727.660 19.030 ;
        RECT 1727.460 2.400 1727.600 18.710 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1697.010 20.640 1697.330 20.700 ;
        RECT 1744.850 20.640 1745.170 20.700 ;
        RECT 1697.010 20.500 1745.170 20.640 ;
        RECT 1697.010 20.440 1697.330 20.500 ;
        RECT 1744.850 20.440 1745.170 20.500 ;
      LAYER via ;
        RECT 1697.040 20.440 1697.300 20.700 ;
        RECT 1744.880 20.440 1745.140 20.700 ;
      LAYER met2 ;
        RECT 1697.100 20.730 1697.240 54.000 ;
        RECT 1697.040 20.410 1697.300 20.730 ;
        RECT 1744.880 20.410 1745.140 20.730 ;
        RECT 1744.940 20.130 1745.080 20.410 ;
        RECT 1744.940 19.990 1745.540 20.130 ;
        RECT 1745.400 2.400 1745.540 19.990 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1710.810 19.280 1711.130 19.340 ;
        RECT 1762.790 19.280 1763.110 19.340 ;
        RECT 1710.810 19.140 1763.110 19.280 ;
        RECT 1710.810 19.080 1711.130 19.140 ;
        RECT 1762.790 19.080 1763.110 19.140 ;
      LAYER via ;
        RECT 1710.840 19.080 1711.100 19.340 ;
        RECT 1762.820 19.080 1763.080 19.340 ;
      LAYER met2 ;
        RECT 1710.900 19.370 1711.040 54.000 ;
        RECT 1710.840 19.050 1711.100 19.370 ;
        RECT 1762.820 19.050 1763.080 19.370 ;
        RECT 1762.880 2.400 1763.020 19.050 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1731.510 18.940 1731.830 19.000 ;
        RECT 1780.730 18.940 1781.050 19.000 ;
        RECT 1731.510 18.800 1781.050 18.940 ;
        RECT 1731.510 18.740 1731.830 18.800 ;
        RECT 1780.730 18.740 1781.050 18.800 ;
      LAYER via ;
        RECT 1731.540 18.740 1731.800 19.000 ;
        RECT 1780.760 18.740 1781.020 19.000 ;
      LAYER met2 ;
        RECT 1731.600 19.030 1731.740 54.000 ;
        RECT 1731.540 18.710 1731.800 19.030 ;
        RECT 1780.760 18.710 1781.020 19.030 ;
        RECT 1780.820 2.400 1780.960 18.710 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1745.310 20.640 1745.630 20.700 ;
        RECT 1798.670 20.640 1798.990 20.700 ;
        RECT 1745.310 20.500 1798.990 20.640 ;
        RECT 1745.310 20.440 1745.630 20.500 ;
        RECT 1798.670 20.440 1798.990 20.500 ;
      LAYER via ;
        RECT 1745.340 20.440 1745.600 20.700 ;
        RECT 1798.700 20.440 1798.960 20.700 ;
      LAYER met2 ;
        RECT 1745.400 20.730 1745.540 54.000 ;
        RECT 1745.340 20.410 1745.600 20.730 ;
        RECT 1798.700 20.410 1798.960 20.730 ;
        RECT 1798.760 2.400 1798.900 20.410 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1759.110 20.300 1759.430 20.360 ;
        RECT 1816.610 20.300 1816.930 20.360 ;
        RECT 1759.110 20.160 1816.930 20.300 ;
        RECT 1759.110 20.100 1759.430 20.160 ;
        RECT 1816.610 20.100 1816.930 20.160 ;
      LAYER via ;
        RECT 1759.140 20.100 1759.400 20.360 ;
        RECT 1816.640 20.100 1816.900 20.360 ;
      LAYER met2 ;
        RECT 1759.200 20.390 1759.340 54.000 ;
        RECT 1759.140 20.070 1759.400 20.390 ;
        RECT 1816.640 20.070 1816.900 20.390 ;
        RECT 1816.700 2.400 1816.840 20.070 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.450 18.260 1772.770 18.320 ;
        RECT 1834.550 18.260 1834.870 18.320 ;
        RECT 1772.450 18.120 1834.870 18.260 ;
        RECT 1772.450 18.060 1772.770 18.120 ;
        RECT 1834.550 18.060 1834.870 18.120 ;
      LAYER via ;
        RECT 1772.480 18.060 1772.740 18.320 ;
        RECT 1834.580 18.060 1834.840 18.320 ;
      LAYER met2 ;
        RECT 1772.540 18.350 1772.680 54.000 ;
        RECT 1772.480 18.030 1772.740 18.350 ;
        RECT 1834.580 18.030 1834.840 18.350 ;
        RECT 1834.640 2.400 1834.780 18.030 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1786.250 17.920 1786.570 17.980 ;
        RECT 1852.030 17.920 1852.350 17.980 ;
        RECT 1786.250 17.780 1852.350 17.920 ;
        RECT 1786.250 17.720 1786.570 17.780 ;
        RECT 1852.030 17.720 1852.350 17.780 ;
      LAYER via ;
        RECT 1786.280 17.720 1786.540 17.980 ;
        RECT 1852.060 17.720 1852.320 17.980 ;
      LAYER met2 ;
        RECT 1786.800 18.090 1786.940 54.000 ;
        RECT 1786.340 18.010 1786.940 18.090 ;
        RECT 1786.280 17.950 1786.940 18.010 ;
        RECT 1786.280 17.690 1786.540 17.950 ;
        RECT 1852.060 17.690 1852.320 18.010 ;
        RECT 1852.120 2.400 1852.260 17.690 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1807.410 15.880 1807.730 15.940 ;
        RECT 1869.970 15.880 1870.290 15.940 ;
        RECT 1807.410 15.740 1870.290 15.880 ;
        RECT 1807.410 15.680 1807.730 15.740 ;
        RECT 1869.970 15.680 1870.290 15.740 ;
      LAYER via ;
        RECT 1807.440 15.680 1807.700 15.940 ;
        RECT 1870.000 15.680 1870.260 15.940 ;
      LAYER met2 ;
        RECT 1807.500 15.970 1807.640 54.000 ;
        RECT 1807.440 15.650 1807.700 15.970 ;
        RECT 1870.000 15.650 1870.260 15.970 ;
        RECT 1870.060 2.400 1870.200 15.650 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 746.190 16.560 746.510 16.620 ;
        RECT 751.710 16.560 752.030 16.620 ;
        RECT 746.190 16.420 752.030 16.560 ;
        RECT 746.190 16.360 746.510 16.420 ;
        RECT 751.710 16.360 752.030 16.420 ;
      LAYER via ;
        RECT 746.220 16.360 746.480 16.620 ;
        RECT 751.740 16.360 752.000 16.620 ;
      LAYER met2 ;
        RECT 751.800 16.650 751.940 54.000 ;
        RECT 746.220 16.330 746.480 16.650 ;
        RECT 751.740 16.330 752.000 16.650 ;
        RECT 746.280 2.400 746.420 16.330 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1821.210 16.220 1821.530 16.280 ;
        RECT 1887.910 16.220 1888.230 16.280 ;
        RECT 1821.210 16.080 1888.230 16.220 ;
        RECT 1821.210 16.020 1821.530 16.080 ;
        RECT 1887.910 16.020 1888.230 16.080 ;
      LAYER via ;
        RECT 1821.240 16.020 1821.500 16.280 ;
        RECT 1887.940 16.020 1888.200 16.280 ;
      LAYER met2 ;
        RECT 1821.300 16.310 1821.440 54.000 ;
        RECT 1821.240 15.990 1821.500 16.310 ;
        RECT 1887.940 15.990 1888.200 16.310 ;
        RECT 1888.000 2.400 1888.140 15.990 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1835.010 20.300 1835.330 20.360 ;
        RECT 1905.850 20.300 1906.170 20.360 ;
        RECT 1835.010 20.160 1906.170 20.300 ;
        RECT 1835.010 20.100 1835.330 20.160 ;
        RECT 1905.850 20.100 1906.170 20.160 ;
      LAYER via ;
        RECT 1835.040 20.100 1835.300 20.360 ;
        RECT 1905.880 20.100 1906.140 20.360 ;
      LAYER met2 ;
        RECT 1835.100 20.390 1835.240 54.000 ;
        RECT 1835.040 20.070 1835.300 20.390 ;
        RECT 1905.880 20.070 1906.140 20.390 ;
        RECT 1905.940 2.400 1906.080 20.070 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1848.810 16.900 1849.130 16.960 ;
        RECT 1923.330 16.900 1923.650 16.960 ;
        RECT 1848.810 16.760 1923.650 16.900 ;
        RECT 1848.810 16.700 1849.130 16.760 ;
        RECT 1923.330 16.700 1923.650 16.760 ;
      LAYER via ;
        RECT 1848.840 16.700 1849.100 16.960 ;
        RECT 1923.360 16.700 1923.620 16.960 ;
      LAYER met2 ;
        RECT 1848.900 16.990 1849.040 54.000 ;
        RECT 1848.840 16.670 1849.100 16.990 ;
        RECT 1923.360 16.670 1923.620 16.990 ;
        RECT 1923.420 2.400 1923.560 16.670 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1869.510 19.960 1869.830 20.020 ;
        RECT 1941.270 19.960 1941.590 20.020 ;
        RECT 1869.510 19.820 1941.590 19.960 ;
        RECT 1869.510 19.760 1869.830 19.820 ;
        RECT 1941.270 19.760 1941.590 19.820 ;
      LAYER via ;
        RECT 1869.540 19.760 1869.800 20.020 ;
        RECT 1941.300 19.760 1941.560 20.020 ;
      LAYER met2 ;
        RECT 1869.600 20.050 1869.740 54.000 ;
        RECT 1869.540 19.730 1869.800 20.050 ;
        RECT 1941.300 19.730 1941.560 20.050 ;
        RECT 1941.360 2.400 1941.500 19.730 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1883.310 15.540 1883.630 15.600 ;
        RECT 1959.210 15.540 1959.530 15.600 ;
        RECT 1883.310 15.400 1959.530 15.540 ;
        RECT 1883.310 15.340 1883.630 15.400 ;
        RECT 1959.210 15.340 1959.530 15.400 ;
      LAYER via ;
        RECT 1883.340 15.340 1883.600 15.600 ;
        RECT 1959.240 15.340 1959.500 15.600 ;
      LAYER met2 ;
        RECT 1883.400 15.630 1883.540 54.000 ;
        RECT 1883.340 15.310 1883.600 15.630 ;
        RECT 1959.240 15.310 1959.500 15.630 ;
        RECT 1959.300 2.400 1959.440 15.310 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1897.110 19.280 1897.430 19.340 ;
        RECT 1977.150 19.280 1977.470 19.340 ;
        RECT 1897.110 19.140 1977.470 19.280 ;
        RECT 1897.110 19.080 1897.430 19.140 ;
        RECT 1977.150 19.080 1977.470 19.140 ;
      LAYER via ;
        RECT 1897.140 19.080 1897.400 19.340 ;
        RECT 1977.180 19.080 1977.440 19.340 ;
      LAYER met2 ;
        RECT 1897.200 19.370 1897.340 54.000 ;
        RECT 1897.140 19.050 1897.400 19.370 ;
        RECT 1977.180 19.050 1977.440 19.370 ;
        RECT 1977.240 2.400 1977.380 19.050 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1910.910 20.300 1911.230 20.360 ;
        RECT 1995.090 20.300 1995.410 20.360 ;
        RECT 1910.910 20.160 1995.410 20.300 ;
        RECT 1910.910 20.100 1911.230 20.160 ;
        RECT 1995.090 20.100 1995.410 20.160 ;
      LAYER via ;
        RECT 1910.940 20.100 1911.200 20.360 ;
        RECT 1995.120 20.100 1995.380 20.360 ;
      LAYER met2 ;
        RECT 1911.000 20.390 1911.140 54.000 ;
        RECT 1910.940 20.070 1911.200 20.390 ;
        RECT 1995.120 20.070 1995.380 20.390 ;
        RECT 1995.180 2.400 1995.320 20.070 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1924.710 15.200 1925.030 15.260 ;
        RECT 2012.570 15.200 2012.890 15.260 ;
        RECT 1924.710 15.060 2012.890 15.200 ;
        RECT 1924.710 15.000 1925.030 15.060 ;
        RECT 2012.570 15.000 2012.890 15.060 ;
      LAYER via ;
        RECT 1924.740 15.000 1925.000 15.260 ;
        RECT 2012.600 15.000 2012.860 15.260 ;
      LAYER met2 ;
        RECT 1924.800 15.290 1924.940 54.000 ;
        RECT 1924.740 14.970 1925.000 15.290 ;
        RECT 2012.600 14.970 2012.860 15.290 ;
        RECT 2012.660 2.400 2012.800 14.970 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1945.410 16.560 1945.730 16.620 ;
        RECT 2030.510 16.560 2030.830 16.620 ;
        RECT 1945.410 16.420 2030.830 16.560 ;
        RECT 1945.410 16.360 1945.730 16.420 ;
        RECT 2030.510 16.360 2030.830 16.420 ;
      LAYER via ;
        RECT 1945.440 16.360 1945.700 16.620 ;
        RECT 2030.540 16.360 2030.800 16.620 ;
      LAYER met2 ;
        RECT 1945.500 16.650 1945.640 54.000 ;
        RECT 1945.440 16.330 1945.700 16.650 ;
        RECT 2030.540 16.330 2030.800 16.650 ;
        RECT 2030.600 2.400 2030.740 16.330 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1959.210 16.900 1959.530 16.960 ;
        RECT 2048.450 16.900 2048.770 16.960 ;
        RECT 1959.210 16.760 2048.770 16.900 ;
        RECT 1959.210 16.700 1959.530 16.760 ;
        RECT 2048.450 16.700 2048.770 16.760 ;
      LAYER via ;
        RECT 1959.240 16.700 1959.500 16.960 ;
        RECT 2048.480 16.700 2048.740 16.960 ;
      LAYER met2 ;
        RECT 1959.300 16.990 1959.440 54.000 ;
        RECT 1959.240 16.670 1959.500 16.990 ;
        RECT 2048.480 16.670 2048.740 16.990 ;
        RECT 2048.540 2.400 2048.680 16.670 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 765.600 17.410 765.740 54.000 ;
        RECT 763.760 17.270 765.740 17.410 ;
        RECT 763.760 2.400 763.900 17.270 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1973.010 18.600 1973.330 18.660 ;
        RECT 2066.390 18.600 2066.710 18.660 ;
        RECT 1973.010 18.460 2066.710 18.600 ;
        RECT 1973.010 18.400 1973.330 18.460 ;
        RECT 2066.390 18.400 2066.710 18.460 ;
      LAYER via ;
        RECT 1973.040 18.400 1973.300 18.660 ;
        RECT 2066.420 18.400 2066.680 18.660 ;
      LAYER met2 ;
        RECT 1973.100 18.690 1973.240 54.000 ;
        RECT 1973.040 18.370 1973.300 18.690 ;
        RECT 2066.420 18.370 2066.680 18.690 ;
        RECT 2066.480 2.400 2066.620 18.370 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1986.810 19.280 1987.130 19.340 ;
        RECT 2084.330 19.280 2084.650 19.340 ;
        RECT 1986.810 19.140 2084.650 19.280 ;
        RECT 1986.810 19.080 1987.130 19.140 ;
        RECT 2084.330 19.080 2084.650 19.140 ;
      LAYER via ;
        RECT 1986.840 19.080 1987.100 19.340 ;
        RECT 2084.360 19.080 2084.620 19.340 ;
      LAYER met2 ;
        RECT 1986.900 19.370 1987.040 54.000 ;
        RECT 1986.840 19.050 1987.100 19.370 ;
        RECT 2084.360 19.050 2084.620 19.370 ;
        RECT 2084.420 2.400 2084.560 19.050 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2007.050 20.300 2007.370 20.360 ;
        RECT 2101.810 20.300 2102.130 20.360 ;
        RECT 2007.050 20.160 2102.130 20.300 ;
        RECT 2007.050 20.100 2007.370 20.160 ;
        RECT 2101.810 20.100 2102.130 20.160 ;
      LAYER via ;
        RECT 2007.080 20.100 2007.340 20.360 ;
        RECT 2101.840 20.100 2102.100 20.360 ;
      LAYER met2 ;
        RECT 2007.140 20.390 2007.280 54.000 ;
        RECT 2007.080 20.070 2007.340 20.390 ;
        RECT 2101.840 20.070 2102.100 20.390 ;
        RECT 2101.900 2.400 2102.040 20.070 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2021.310 16.220 2021.630 16.280 ;
        RECT 2119.750 16.220 2120.070 16.280 ;
        RECT 2021.310 16.080 2120.070 16.220 ;
        RECT 2021.310 16.020 2021.630 16.080 ;
        RECT 2119.750 16.020 2120.070 16.080 ;
      LAYER via ;
        RECT 2021.340 16.020 2021.600 16.280 ;
        RECT 2119.780 16.020 2120.040 16.280 ;
      LAYER met2 ;
        RECT 2021.400 16.310 2021.540 54.000 ;
        RECT 2021.340 15.990 2021.600 16.310 ;
        RECT 2119.780 15.990 2120.040 16.310 ;
        RECT 2119.840 2.400 2119.980 15.990 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2035.110 16.560 2035.430 16.620 ;
        RECT 2137.690 16.560 2138.010 16.620 ;
        RECT 2035.110 16.420 2138.010 16.560 ;
        RECT 2035.110 16.360 2035.430 16.420 ;
        RECT 2137.690 16.360 2138.010 16.420 ;
      LAYER via ;
        RECT 2035.140 16.360 2035.400 16.620 ;
        RECT 2137.720 16.360 2137.980 16.620 ;
      LAYER met2 ;
        RECT 2035.200 16.650 2035.340 54.000 ;
        RECT 2035.140 16.330 2035.400 16.650 ;
        RECT 2137.720 16.330 2137.980 16.650 ;
        RECT 2137.780 2.400 2137.920 16.330 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2048.910 17.920 2049.230 17.980 ;
        RECT 2155.630 17.920 2155.950 17.980 ;
        RECT 2048.910 17.780 2155.950 17.920 ;
        RECT 2048.910 17.720 2049.230 17.780 ;
        RECT 2155.630 17.720 2155.950 17.780 ;
      LAYER via ;
        RECT 2048.940 17.720 2049.200 17.980 ;
        RECT 2155.660 17.720 2155.920 17.980 ;
      LAYER met2 ;
        RECT 2049.000 18.010 2049.140 54.000 ;
        RECT 2048.940 17.690 2049.200 18.010 ;
        RECT 2155.660 17.690 2155.920 18.010 ;
        RECT 2155.720 2.400 2155.860 17.690 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2062.710 16.900 2063.030 16.960 ;
        RECT 2111.470 16.900 2111.790 16.960 ;
        RECT 2062.710 16.760 2111.790 16.900 ;
        RECT 2062.710 16.700 2063.030 16.760 ;
        RECT 2111.470 16.700 2111.790 16.760 ;
        RECT 2173.110 16.560 2173.430 16.620 ;
        RECT 2138.240 16.420 2173.430 16.560 ;
        RECT 2111.470 15.880 2111.790 15.940 ;
        RECT 2138.240 15.880 2138.380 16.420 ;
        RECT 2173.110 16.360 2173.430 16.420 ;
        RECT 2111.470 15.740 2138.380 15.880 ;
        RECT 2111.470 15.680 2111.790 15.740 ;
      LAYER via ;
        RECT 2062.740 16.700 2063.000 16.960 ;
        RECT 2111.500 16.700 2111.760 16.960 ;
        RECT 2111.500 15.680 2111.760 15.940 ;
        RECT 2173.140 16.360 2173.400 16.620 ;
      LAYER met2 ;
        RECT 2062.800 16.990 2062.940 54.000 ;
        RECT 2062.740 16.670 2063.000 16.990 ;
        RECT 2111.500 16.670 2111.760 16.990 ;
        RECT 2111.560 15.970 2111.700 16.670 ;
        RECT 2173.140 16.330 2173.400 16.650 ;
        RECT 2111.500 15.650 2111.760 15.970 ;
        RECT 2173.200 2.400 2173.340 16.330 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2083.410 15.200 2083.730 15.260 ;
        RECT 2191.050 15.200 2191.370 15.260 ;
        RECT 2083.410 15.060 2191.370 15.200 ;
        RECT 2083.410 15.000 2083.730 15.060 ;
        RECT 2191.050 15.000 2191.370 15.060 ;
      LAYER via ;
        RECT 2083.440 15.000 2083.700 15.260 ;
        RECT 2191.080 15.000 2191.340 15.260 ;
      LAYER met2 ;
        RECT 2083.500 15.290 2083.640 54.000 ;
        RECT 2083.440 14.970 2083.700 15.290 ;
        RECT 2191.080 14.970 2191.340 15.290 ;
        RECT 2191.140 2.400 2191.280 14.970 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2097.210 19.620 2097.530 19.680 ;
        RECT 2208.990 19.620 2209.310 19.680 ;
        RECT 2097.210 19.480 2209.310 19.620 ;
        RECT 2097.210 19.420 2097.530 19.480 ;
        RECT 2208.990 19.420 2209.310 19.480 ;
      LAYER via ;
        RECT 2097.240 19.420 2097.500 19.680 ;
        RECT 2209.020 19.420 2209.280 19.680 ;
      LAYER met2 ;
        RECT 2097.300 19.710 2097.440 54.000 ;
        RECT 2097.240 19.390 2097.500 19.710 ;
        RECT 2209.020 19.390 2209.280 19.710 ;
        RECT 2209.080 2.400 2209.220 19.390 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2111.010 15.540 2111.330 15.600 ;
        RECT 2226.930 15.540 2227.250 15.600 ;
        RECT 2111.010 15.400 2227.250 15.540 ;
        RECT 2111.010 15.340 2111.330 15.400 ;
        RECT 2226.930 15.340 2227.250 15.400 ;
      LAYER via ;
        RECT 2111.040 15.340 2111.300 15.600 ;
        RECT 2226.960 15.340 2227.220 15.600 ;
      LAYER met2 ;
        RECT 2111.100 15.630 2111.240 54.000 ;
        RECT 2111.040 15.310 2111.300 15.630 ;
        RECT 2226.960 15.310 2227.220 15.630 ;
        RECT 2227.020 2.400 2227.160 15.310 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 781.610 17.580 781.930 17.640 ;
        RECT 786.210 17.580 786.530 17.640 ;
        RECT 781.610 17.440 786.530 17.580 ;
        RECT 781.610 17.380 781.930 17.440 ;
        RECT 786.210 17.380 786.530 17.440 ;
      LAYER via ;
        RECT 781.640 17.380 781.900 17.640 ;
        RECT 786.240 17.380 786.500 17.640 ;
      LAYER met2 ;
        RECT 786.300 17.670 786.440 54.000 ;
        RECT 781.640 17.350 781.900 17.670 ;
        RECT 786.240 17.350 786.500 17.670 ;
        RECT 781.700 2.400 781.840 17.350 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2124.810 19.280 2125.130 19.340 ;
        RECT 2244.870 19.280 2245.190 19.340 ;
        RECT 2124.810 19.140 2245.190 19.280 ;
        RECT 2124.810 19.080 2125.130 19.140 ;
        RECT 2244.870 19.080 2245.190 19.140 ;
      LAYER via ;
        RECT 2124.840 19.080 2125.100 19.340 ;
        RECT 2244.900 19.080 2245.160 19.340 ;
      LAYER met2 ;
        RECT 2124.900 19.370 2125.040 54.000 ;
        RECT 2124.840 19.050 2125.100 19.370 ;
        RECT 2244.900 19.050 2245.160 19.370 ;
        RECT 2244.960 2.400 2245.100 19.050 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2138.610 16.220 2138.930 16.280 ;
        RECT 2262.350 16.220 2262.670 16.280 ;
        RECT 2138.610 16.080 2262.670 16.220 ;
        RECT 2138.610 16.020 2138.930 16.080 ;
        RECT 2262.350 16.020 2262.670 16.080 ;
      LAYER via ;
        RECT 2138.640 16.020 2138.900 16.280 ;
        RECT 2262.380 16.020 2262.640 16.280 ;
      LAYER met2 ;
        RECT 2138.700 16.310 2138.840 54.000 ;
        RECT 2138.640 15.990 2138.900 16.310 ;
        RECT 2262.380 15.990 2262.640 16.310 ;
        RECT 2262.440 2.400 2262.580 15.990 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2159.310 18.940 2159.630 19.000 ;
        RECT 2280.290 18.940 2280.610 19.000 ;
        RECT 2159.310 18.800 2280.610 18.940 ;
        RECT 2159.310 18.740 2159.630 18.800 ;
        RECT 2280.290 18.740 2280.610 18.800 ;
      LAYER via ;
        RECT 2159.340 18.740 2159.600 19.000 ;
        RECT 2280.320 18.740 2280.580 19.000 ;
      LAYER met2 ;
        RECT 2159.400 19.030 2159.540 54.000 ;
        RECT 2159.340 18.710 2159.600 19.030 ;
        RECT 2280.320 18.710 2280.580 19.030 ;
        RECT 2280.380 2.400 2280.520 18.710 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2173.570 16.900 2173.890 16.960 ;
        RECT 2298.230 16.900 2298.550 16.960 ;
        RECT 2173.570 16.760 2298.550 16.900 ;
        RECT 2173.570 16.700 2173.890 16.760 ;
        RECT 2298.230 16.700 2298.550 16.760 ;
      LAYER via ;
        RECT 2173.600 16.700 2173.860 16.960 ;
        RECT 2298.260 16.700 2298.520 16.960 ;
      LAYER met2 ;
        RECT 2173.200 17.410 2173.340 54.000 ;
        RECT 2173.200 17.270 2173.800 17.410 ;
        RECT 2173.660 16.990 2173.800 17.270 ;
        RECT 2173.600 16.670 2173.860 16.990 ;
        RECT 2298.260 16.670 2298.520 16.990 ;
        RECT 2298.320 2.400 2298.460 16.670 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2186.910 16.560 2187.230 16.620 ;
        RECT 2316.170 16.560 2316.490 16.620 ;
        RECT 2186.910 16.420 2316.490 16.560 ;
        RECT 2186.910 16.360 2187.230 16.420 ;
        RECT 2316.170 16.360 2316.490 16.420 ;
      LAYER via ;
        RECT 2186.940 16.360 2187.200 16.620 ;
        RECT 2316.200 16.360 2316.460 16.620 ;
      LAYER met2 ;
        RECT 2187.000 16.650 2187.140 54.000 ;
        RECT 2186.940 16.330 2187.200 16.650 ;
        RECT 2316.200 16.330 2316.460 16.650 ;
        RECT 2316.260 2.400 2316.400 16.330 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2200.710 17.580 2201.030 17.640 ;
        RECT 2334.110 17.580 2334.430 17.640 ;
        RECT 2200.710 17.440 2334.430 17.580 ;
        RECT 2200.710 17.380 2201.030 17.440 ;
        RECT 2334.110 17.380 2334.430 17.440 ;
      LAYER via ;
        RECT 2200.740 17.380 2201.000 17.640 ;
        RECT 2334.140 17.380 2334.400 17.640 ;
      LAYER met2 ;
        RECT 2200.800 17.670 2200.940 54.000 ;
        RECT 2200.740 17.350 2201.000 17.670 ;
        RECT 2334.140 17.350 2334.400 17.670 ;
        RECT 2334.200 2.400 2334.340 17.350 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2221.410 14.180 2221.730 14.240 ;
        RECT 2351.590 14.180 2351.910 14.240 ;
        RECT 2221.410 14.040 2351.910 14.180 ;
        RECT 2221.410 13.980 2221.730 14.040 ;
        RECT 2351.590 13.980 2351.910 14.040 ;
      LAYER via ;
        RECT 2221.440 13.980 2221.700 14.240 ;
        RECT 2351.620 13.980 2351.880 14.240 ;
      LAYER met2 ;
        RECT 2221.500 14.270 2221.640 54.000 ;
        RECT 2221.440 13.950 2221.700 14.270 ;
        RECT 2351.620 13.950 2351.880 14.270 ;
        RECT 2351.680 2.400 2351.820 13.950 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2235.210 20.300 2235.530 20.360 ;
        RECT 2369.530 20.300 2369.850 20.360 ;
        RECT 2235.210 20.160 2369.850 20.300 ;
        RECT 2235.210 20.100 2235.530 20.160 ;
        RECT 2369.530 20.100 2369.850 20.160 ;
      LAYER via ;
        RECT 2235.240 20.100 2235.500 20.360 ;
        RECT 2369.560 20.100 2369.820 20.360 ;
      LAYER met2 ;
        RECT 2235.300 20.390 2235.440 54.000 ;
        RECT 2235.240 20.070 2235.500 20.390 ;
        RECT 2369.560 20.070 2369.820 20.390 ;
        RECT 2369.620 2.400 2369.760 20.070 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2249.010 20.640 2249.330 20.700 ;
        RECT 2387.470 20.640 2387.790 20.700 ;
        RECT 2249.010 20.500 2387.790 20.640 ;
        RECT 2249.010 20.440 2249.330 20.500 ;
        RECT 2387.470 20.440 2387.790 20.500 ;
      LAYER via ;
        RECT 2249.040 20.440 2249.300 20.700 ;
        RECT 2387.500 20.440 2387.760 20.700 ;
      LAYER met2 ;
        RECT 2249.100 20.730 2249.240 54.000 ;
        RECT 2249.040 20.410 2249.300 20.730 ;
        RECT 2387.500 20.410 2387.760 20.730 ;
        RECT 2387.560 2.400 2387.700 20.410 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2262.810 16.220 2263.130 16.280 ;
        RECT 2405.410 16.220 2405.730 16.280 ;
        RECT 2262.810 16.080 2405.730 16.220 ;
        RECT 2262.810 16.020 2263.130 16.080 ;
        RECT 2405.410 16.020 2405.730 16.080 ;
      LAYER via ;
        RECT 2262.840 16.020 2263.100 16.280 ;
        RECT 2405.440 16.020 2405.700 16.280 ;
      LAYER met2 ;
        RECT 2262.900 16.310 2263.040 54.000 ;
        RECT 2262.840 15.990 2263.100 16.310 ;
        RECT 2405.440 15.990 2405.700 16.310 ;
        RECT 2405.500 2.400 2405.640 15.990 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 800.100 17.410 800.240 54.000 ;
        RECT 799.640 17.270 800.240 17.410 ;
        RECT 799.640 2.400 799.780 17.270 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 644.990 17.580 645.310 17.640 ;
        RECT 648.210 17.580 648.530 17.640 ;
        RECT 644.990 17.440 648.530 17.580 ;
        RECT 644.990 17.380 645.310 17.440 ;
        RECT 648.210 17.380 648.530 17.440 ;
      LAYER via ;
        RECT 645.020 17.380 645.280 17.640 ;
        RECT 648.240 17.380 648.500 17.640 ;
      LAYER met2 ;
        RECT 648.300 17.670 648.440 54.000 ;
        RECT 645.020 17.350 645.280 17.670 ;
        RECT 648.240 17.350 648.500 17.670 ;
        RECT 645.080 2.400 645.220 17.350 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2283.510 18.940 2283.830 19.000 ;
        RECT 2428.870 18.940 2429.190 19.000 ;
        RECT 2283.510 18.800 2429.190 18.940 ;
        RECT 2283.510 18.740 2283.830 18.800 ;
        RECT 2428.870 18.740 2429.190 18.800 ;
      LAYER via ;
        RECT 2283.540 18.740 2283.800 19.000 ;
        RECT 2428.900 18.740 2429.160 19.000 ;
      LAYER met2 ;
        RECT 2283.600 19.030 2283.740 54.000 ;
        RECT 2283.540 18.710 2283.800 19.030 ;
        RECT 2428.900 18.710 2429.160 19.030 ;
        RECT 2428.960 2.400 2429.100 18.710 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2297.310 19.280 2297.630 19.340 ;
        RECT 2446.810 19.280 2447.130 19.340 ;
        RECT 2297.310 19.140 2447.130 19.280 ;
        RECT 2297.310 19.080 2297.630 19.140 ;
        RECT 2446.810 19.080 2447.130 19.140 ;
      LAYER via ;
        RECT 2297.340 19.080 2297.600 19.340 ;
        RECT 2446.840 19.080 2447.100 19.340 ;
      LAYER met2 ;
        RECT 2297.400 19.370 2297.540 54.000 ;
        RECT 2297.340 19.050 2297.600 19.370 ;
        RECT 2446.840 19.050 2447.100 19.370 ;
        RECT 2446.900 2.400 2447.040 19.050 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2346.530 17.920 2346.850 17.980 ;
        RECT 2464.750 17.920 2465.070 17.980 ;
        RECT 2346.530 17.780 2465.070 17.920 ;
        RECT 2346.530 17.720 2346.850 17.780 ;
        RECT 2464.750 17.720 2465.070 17.780 ;
        RECT 2318.010 16.900 2318.330 16.960 ;
        RECT 2346.530 16.900 2346.850 16.960 ;
        RECT 2318.010 16.760 2346.850 16.900 ;
        RECT 2318.010 16.700 2318.330 16.760 ;
        RECT 2346.530 16.700 2346.850 16.760 ;
      LAYER via ;
        RECT 2346.560 17.720 2346.820 17.980 ;
        RECT 2464.780 17.720 2465.040 17.980 ;
        RECT 2318.040 16.700 2318.300 16.960 ;
        RECT 2346.560 16.700 2346.820 16.960 ;
      LAYER met2 ;
        RECT 2318.100 16.990 2318.240 54.000 ;
        RECT 2346.560 17.690 2346.820 18.010 ;
        RECT 2464.780 17.690 2465.040 18.010 ;
        RECT 2346.620 16.990 2346.760 17.690 ;
        RECT 2318.040 16.670 2318.300 16.990 ;
        RECT 2346.560 16.670 2346.820 16.990 ;
        RECT 2464.840 2.400 2464.980 17.690 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2331.810 16.560 2332.130 16.620 ;
        RECT 2482.690 16.560 2483.010 16.620 ;
        RECT 2331.810 16.420 2483.010 16.560 ;
        RECT 2331.810 16.360 2332.130 16.420 ;
        RECT 2482.690 16.360 2483.010 16.420 ;
      LAYER via ;
        RECT 2331.840 16.360 2332.100 16.620 ;
        RECT 2482.720 16.360 2482.980 16.620 ;
      LAYER met2 ;
        RECT 2331.900 16.650 2332.040 54.000 ;
        RECT 2331.840 16.330 2332.100 16.650 ;
        RECT 2482.720 16.330 2482.980 16.650 ;
        RECT 2482.780 2.400 2482.920 16.330 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2345.610 18.600 2345.930 18.660 ;
        RECT 2500.630 18.600 2500.950 18.660 ;
        RECT 2345.610 18.460 2500.950 18.600 ;
        RECT 2345.610 18.400 2345.930 18.460 ;
        RECT 2500.630 18.400 2500.950 18.460 ;
      LAYER via ;
        RECT 2345.640 18.400 2345.900 18.660 ;
        RECT 2500.660 18.400 2500.920 18.660 ;
      LAYER met2 ;
        RECT 2345.700 18.690 2345.840 54.000 ;
        RECT 2345.640 18.370 2345.900 18.690 ;
        RECT 2500.660 18.370 2500.920 18.690 ;
        RECT 2500.720 2.400 2500.860 18.370 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2418.290 15.200 2418.610 15.260 ;
        RECT 2518.110 15.200 2518.430 15.260 ;
        RECT 2418.290 15.060 2518.430 15.200 ;
        RECT 2418.290 15.000 2418.610 15.060 ;
        RECT 2518.110 15.000 2518.430 15.060 ;
      LAYER via ;
        RECT 2418.320 15.000 2418.580 15.260 ;
        RECT 2518.140 15.000 2518.400 15.260 ;
      LAYER met2 ;
        RECT 2418.380 15.290 2418.520 54.000 ;
        RECT 2418.320 14.970 2418.580 15.290 ;
        RECT 2518.140 14.970 2518.400 15.290 ;
        RECT 2518.200 2.400 2518.340 14.970 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2480.390 16.900 2480.710 16.960 ;
        RECT 2536.050 16.900 2536.370 16.960 ;
        RECT 2480.390 16.760 2536.370 16.900 ;
        RECT 2480.390 16.700 2480.710 16.760 ;
        RECT 2536.050 16.700 2536.370 16.760 ;
      LAYER via ;
        RECT 2480.420 16.700 2480.680 16.960 ;
        RECT 2536.080 16.700 2536.340 16.960 ;
      LAYER met2 ;
        RECT 2480.480 16.990 2480.620 54.000 ;
        RECT 2480.420 16.670 2480.680 16.990 ;
        RECT 2536.080 16.670 2536.340 16.990 ;
        RECT 2536.140 2.400 2536.280 16.670 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2542.490 20.640 2542.810 20.700 ;
        RECT 2553.990 20.640 2554.310 20.700 ;
        RECT 2542.490 20.500 2554.310 20.640 ;
        RECT 2542.490 20.440 2542.810 20.500 ;
        RECT 2553.990 20.440 2554.310 20.500 ;
      LAYER via ;
        RECT 2542.520 20.440 2542.780 20.700 ;
        RECT 2554.020 20.440 2554.280 20.700 ;
      LAYER met2 ;
        RECT 2542.580 20.730 2542.720 54.000 ;
        RECT 2542.520 20.410 2542.780 20.730 ;
        RECT 2554.020 20.410 2554.280 20.730 ;
        RECT 2554.080 2.400 2554.220 20.410 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2407.710 16.220 2408.030 16.280 ;
        RECT 2571.930 16.220 2572.250 16.280 ;
        RECT 2407.710 16.080 2572.250 16.220 ;
        RECT 2407.710 16.020 2408.030 16.080 ;
        RECT 2571.930 16.020 2572.250 16.080 ;
      LAYER via ;
        RECT 2407.740 16.020 2408.000 16.280 ;
        RECT 2571.960 16.020 2572.220 16.280 ;
      LAYER met2 ;
        RECT 2407.800 16.310 2407.940 54.000 ;
        RECT 2407.740 15.990 2408.000 16.310 ;
        RECT 2571.960 15.990 2572.220 16.310 ;
        RECT 2572.020 2.400 2572.160 15.990 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2563.190 15.200 2563.510 15.260 ;
        RECT 2589.410 15.200 2589.730 15.260 ;
        RECT 2563.190 15.060 2589.730 15.200 ;
        RECT 2563.190 15.000 2563.510 15.060 ;
        RECT 2589.410 15.000 2589.730 15.060 ;
      LAYER via ;
        RECT 2563.220 15.000 2563.480 15.260 ;
        RECT 2589.440 15.000 2589.700 15.260 ;
      LAYER met2 ;
        RECT 2563.280 15.290 2563.420 54.000 ;
        RECT 2563.220 14.970 2563.480 15.290 ;
        RECT 2589.440 14.970 2589.700 15.290 ;
        RECT 2589.500 2.400 2589.640 14.970 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 823.470 17.240 823.790 17.300 ;
        RECT 827.610 17.240 827.930 17.300 ;
        RECT 823.470 17.100 827.930 17.240 ;
        RECT 823.470 17.040 823.790 17.100 ;
        RECT 827.610 17.040 827.930 17.100 ;
      LAYER via ;
        RECT 823.500 17.040 823.760 17.300 ;
        RECT 827.640 17.040 827.900 17.300 ;
      LAYER met2 ;
        RECT 827.700 17.330 827.840 54.000 ;
        RECT 823.500 17.010 823.760 17.330 ;
        RECT 827.640 17.010 827.900 17.330 ;
        RECT 823.560 2.400 823.700 17.010 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2584.810 20.300 2585.130 20.360 ;
        RECT 2607.350 20.300 2607.670 20.360 ;
        RECT 2584.810 20.160 2607.670 20.300 ;
        RECT 2584.810 20.100 2585.130 20.160 ;
        RECT 2607.350 20.100 2607.670 20.160 ;
      LAYER via ;
        RECT 2584.840 20.100 2585.100 20.360 ;
        RECT 2607.380 20.100 2607.640 20.360 ;
      LAYER met2 ;
        RECT 2584.900 20.390 2585.040 54.000 ;
        RECT 2584.840 20.070 2585.100 20.390 ;
        RECT 2607.380 20.070 2607.640 20.390 ;
        RECT 2607.440 2.400 2607.580 20.070 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2605.510 15.200 2605.830 15.260 ;
        RECT 2625.290 15.200 2625.610 15.260 ;
        RECT 2605.510 15.060 2625.610 15.200 ;
        RECT 2605.510 15.000 2605.830 15.060 ;
        RECT 2625.290 15.000 2625.610 15.060 ;
      LAYER via ;
        RECT 2605.540 15.000 2605.800 15.260 ;
        RECT 2625.320 15.000 2625.580 15.260 ;
      LAYER met2 ;
        RECT 2605.600 15.290 2605.740 54.000 ;
        RECT 2605.540 14.970 2605.800 15.290 ;
        RECT 2625.320 14.970 2625.580 15.290 ;
        RECT 2625.380 2.400 2625.520 14.970 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2469.810 15.540 2470.130 15.600 ;
        RECT 2643.230 15.540 2643.550 15.600 ;
        RECT 2469.810 15.400 2643.550 15.540 ;
        RECT 2469.810 15.340 2470.130 15.400 ;
        RECT 2643.230 15.340 2643.550 15.400 ;
      LAYER via ;
        RECT 2469.840 15.340 2470.100 15.600 ;
        RECT 2643.260 15.340 2643.520 15.600 ;
      LAYER met2 ;
        RECT 2469.900 15.630 2470.040 54.000 ;
        RECT 2469.840 15.310 2470.100 15.630 ;
        RECT 2643.260 15.310 2643.520 15.630 ;
        RECT 2643.320 2.400 2643.460 15.310 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2645.990 14.520 2646.310 14.580 ;
        RECT 2661.170 14.520 2661.490 14.580 ;
        RECT 2645.990 14.380 2661.490 14.520 ;
        RECT 2645.990 14.320 2646.310 14.380 ;
        RECT 2661.170 14.320 2661.490 14.380 ;
      LAYER via ;
        RECT 2646.020 14.320 2646.280 14.580 ;
        RECT 2661.200 14.320 2661.460 14.580 ;
      LAYER met2 ;
        RECT 2646.080 14.610 2646.220 54.000 ;
        RECT 2646.020 14.290 2646.280 14.610 ;
        RECT 2661.200 14.290 2661.460 14.610 ;
        RECT 2661.260 2.400 2661.400 14.290 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2496.950 17.580 2497.270 17.640 ;
        RECT 2678.650 17.580 2678.970 17.640 ;
        RECT 2496.950 17.440 2678.970 17.580 ;
        RECT 2496.950 17.380 2497.270 17.440 ;
        RECT 2678.650 17.380 2678.970 17.440 ;
      LAYER via ;
        RECT 2496.980 17.380 2497.240 17.640 ;
        RECT 2678.680 17.380 2678.940 17.640 ;
      LAYER met2 ;
        RECT 2497.040 17.670 2497.180 54.000 ;
        RECT 2496.980 17.350 2497.240 17.670 ;
        RECT 2678.680 17.350 2678.940 17.670 ;
        RECT 2678.740 2.400 2678.880 17.350 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2691.530 2.960 2691.850 3.020 ;
        RECT 2696.590 2.960 2696.910 3.020 ;
        RECT 2691.530 2.820 2696.910 2.960 ;
        RECT 2691.530 2.760 2691.850 2.820 ;
        RECT 2696.590 2.760 2696.910 2.820 ;
      LAYER via ;
        RECT 2691.560 2.760 2691.820 3.020 ;
        RECT 2696.620 2.760 2696.880 3.020 ;
      LAYER met2 ;
        RECT 2691.620 3.050 2691.760 54.000 ;
        RECT 2691.560 2.730 2691.820 3.050 ;
        RECT 2696.620 2.730 2696.880 3.050 ;
        RECT 2696.680 2.400 2696.820 2.730 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2711.770 2.960 2712.090 3.020 ;
        RECT 2714.530 2.960 2714.850 3.020 ;
        RECT 2711.770 2.820 2714.850 2.960 ;
        RECT 2711.770 2.760 2712.090 2.820 ;
        RECT 2714.530 2.760 2714.850 2.820 ;
      LAYER via ;
        RECT 2711.800 2.760 2712.060 3.020 ;
        RECT 2714.560 2.760 2714.820 3.020 ;
      LAYER met2 ;
        RECT 2711.860 3.050 2712.000 54.000 ;
        RECT 2711.800 2.730 2712.060 3.050 ;
        RECT 2714.560 2.730 2714.820 3.050 ;
        RECT 2714.620 2.400 2714.760 2.730 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2721.890 16.560 2722.210 16.620 ;
        RECT 2732.470 16.560 2732.790 16.620 ;
        RECT 2721.890 16.420 2732.790 16.560 ;
        RECT 2721.890 16.360 2722.210 16.420 ;
        RECT 2732.470 16.360 2732.790 16.420 ;
      LAYER via ;
        RECT 2721.920 16.360 2722.180 16.620 ;
        RECT 2732.500 16.360 2732.760 16.620 ;
      LAYER met2 ;
        RECT 2721.980 16.650 2722.120 54.000 ;
        RECT 2721.920 16.330 2722.180 16.650 ;
        RECT 2732.500 16.330 2732.760 16.650 ;
        RECT 2732.560 2.400 2732.700 16.330 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2559.510 16.900 2559.830 16.960 ;
        RECT 2750.410 16.900 2750.730 16.960 ;
        RECT 2559.510 16.760 2750.730 16.900 ;
        RECT 2559.510 16.700 2559.830 16.760 ;
        RECT 2750.410 16.700 2750.730 16.760 ;
      LAYER via ;
        RECT 2559.540 16.700 2559.800 16.960 ;
        RECT 2750.440 16.700 2750.700 16.960 ;
      LAYER met2 ;
        RECT 2559.600 16.990 2559.740 54.000 ;
        RECT 2559.540 16.670 2559.800 16.990 ;
        RECT 2750.440 16.670 2750.700 16.990 ;
        RECT 2750.500 2.400 2750.640 16.670 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2728.790 14.180 2729.110 14.240 ;
        RECT 2767.890 14.180 2768.210 14.240 ;
        RECT 2728.790 14.040 2768.210 14.180 ;
        RECT 2728.790 13.980 2729.110 14.040 ;
        RECT 2767.890 13.980 2768.210 14.040 ;
      LAYER via ;
        RECT 2728.820 13.980 2729.080 14.240 ;
        RECT 2767.920 13.980 2768.180 14.240 ;
      LAYER met2 ;
        RECT 2728.880 14.270 2729.020 54.000 ;
        RECT 2728.820 13.950 2729.080 14.270 ;
        RECT 2767.920 13.950 2768.180 14.270 ;
        RECT 2767.980 2.400 2768.120 13.950 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 841.500 17.410 841.640 54.000 ;
        RECT 841.040 17.270 841.640 17.410 ;
        RECT 841.040 2.400 841.180 17.270 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2594.010 19.620 2594.330 19.680 ;
        RECT 2785.830 19.620 2786.150 19.680 ;
        RECT 2594.010 19.480 2786.150 19.620 ;
        RECT 2594.010 19.420 2594.330 19.480 ;
        RECT 2785.830 19.420 2786.150 19.480 ;
      LAYER via ;
        RECT 2594.040 19.420 2594.300 19.680 ;
        RECT 2785.860 19.420 2786.120 19.680 ;
      LAYER met2 ;
        RECT 2594.100 19.710 2594.240 54.000 ;
        RECT 2594.040 19.390 2594.300 19.710 ;
        RECT 2785.860 19.390 2786.120 19.710 ;
        RECT 2785.920 2.400 2786.060 19.390 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2607.810 18.940 2608.130 19.000 ;
        RECT 2803.770 18.940 2804.090 19.000 ;
        RECT 2607.810 18.800 2804.090 18.940 ;
        RECT 2607.810 18.740 2608.130 18.800 ;
        RECT 2803.770 18.740 2804.090 18.800 ;
      LAYER via ;
        RECT 2607.840 18.740 2608.100 19.000 ;
        RECT 2803.800 18.740 2804.060 19.000 ;
      LAYER met2 ;
        RECT 2607.900 19.030 2608.040 54.000 ;
        RECT 2607.840 18.710 2608.100 19.030 ;
        RECT 2803.800 18.710 2804.060 19.030 ;
        RECT 2803.860 2.400 2804.000 18.710 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2621.610 19.280 2621.930 19.340 ;
        RECT 2821.710 19.280 2822.030 19.340 ;
        RECT 2621.610 19.140 2822.030 19.280 ;
        RECT 2621.610 19.080 2621.930 19.140 ;
        RECT 2821.710 19.080 2822.030 19.140 ;
      LAYER via ;
        RECT 2621.640 19.080 2621.900 19.340 ;
        RECT 2821.740 19.080 2822.000 19.340 ;
      LAYER met2 ;
        RECT 2621.700 19.370 2621.840 54.000 ;
        RECT 2621.640 19.050 2621.900 19.370 ;
        RECT 2821.740 19.050 2822.000 19.370 ;
        RECT 2821.800 2.400 2821.940 19.050 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2839.190 14.860 2839.510 14.920 ;
        RECT 2763.840 14.720 2839.510 14.860 ;
        RECT 2736.150 14.520 2736.470 14.580 ;
        RECT 2763.840 14.520 2763.980 14.720 ;
        RECT 2839.190 14.660 2839.510 14.720 ;
        RECT 2736.150 14.380 2763.980 14.520 ;
        RECT 2736.150 14.320 2736.470 14.380 ;
      LAYER via ;
        RECT 2736.180 14.320 2736.440 14.580 ;
        RECT 2839.220 14.660 2839.480 14.920 ;
      LAYER met2 ;
        RECT 2736.240 14.610 2736.380 54.000 ;
        RECT 2839.220 14.630 2839.480 14.950 ;
        RECT 2736.180 14.290 2736.440 14.610 ;
        RECT 2839.280 2.400 2839.420 14.630 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2648.290 17.240 2648.610 17.300 ;
        RECT 2857.130 17.240 2857.450 17.300 ;
        RECT 2648.290 17.100 2857.450 17.240 ;
        RECT 2648.290 17.040 2648.610 17.100 ;
        RECT 2857.130 17.040 2857.450 17.100 ;
      LAYER via ;
        RECT 2648.320 17.040 2648.580 17.300 ;
        RECT 2857.160 17.040 2857.420 17.300 ;
      LAYER met2 ;
        RECT 2649.300 25.570 2649.440 54.000 ;
        RECT 2648.380 25.430 2649.440 25.570 ;
        RECT 2648.380 17.330 2648.520 25.430 ;
        RECT 2648.320 17.010 2648.580 17.330 ;
        RECT 2857.160 17.010 2857.420 17.330 ;
        RECT 2857.220 2.400 2857.360 17.010 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2735.690 20.300 2736.010 20.360 ;
        RECT 2875.070 20.300 2875.390 20.360 ;
        RECT 2735.690 20.160 2875.390 20.300 ;
        RECT 2735.690 20.100 2736.010 20.160 ;
        RECT 2875.070 20.100 2875.390 20.160 ;
      LAYER via ;
        RECT 2735.720 20.100 2735.980 20.360 ;
        RECT 2875.100 20.100 2875.360 20.360 ;
      LAYER met2 ;
        RECT 2735.780 20.390 2735.920 54.000 ;
        RECT 2735.720 20.070 2735.980 20.390 ;
        RECT 2875.100 20.070 2875.360 20.390 ;
        RECT 2875.160 2.400 2875.300 20.070 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2683.710 17.580 2684.030 17.640 ;
        RECT 2893.010 17.580 2893.330 17.640 ;
        RECT 2683.710 17.440 2893.330 17.580 ;
        RECT 2683.710 17.380 2684.030 17.440 ;
        RECT 2893.010 17.380 2893.330 17.440 ;
      LAYER via ;
        RECT 2683.740 17.380 2684.000 17.640 ;
        RECT 2893.040 17.380 2893.300 17.640 ;
      LAYER met2 ;
        RECT 2683.800 17.670 2683.940 54.000 ;
        RECT 2683.740 17.350 2684.000 17.670 ;
        RECT 2893.040 17.350 2893.300 17.670 ;
        RECT 2893.100 2.400 2893.240 17.350 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2742.590 19.960 2742.910 20.020 ;
        RECT 2910.950 19.960 2911.270 20.020 ;
        RECT 2742.590 19.820 2911.270 19.960 ;
        RECT 2742.590 19.760 2742.910 19.820 ;
        RECT 2910.950 19.760 2911.270 19.820 ;
      LAYER via ;
        RECT 2742.620 19.760 2742.880 20.020 ;
        RECT 2910.980 19.760 2911.240 20.020 ;
      LAYER met2 ;
        RECT 2742.680 20.050 2742.820 54.000 ;
        RECT 2742.620 19.730 2742.880 20.050 ;
        RECT 2910.980 19.730 2911.240 20.050 ;
        RECT 2911.040 2.400 2911.180 19.730 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 858.890 17.580 859.210 17.640 ;
        RECT 862.110 17.580 862.430 17.640 ;
        RECT 858.890 17.440 862.430 17.580 ;
        RECT 858.890 17.380 859.210 17.440 ;
        RECT 862.110 17.380 862.430 17.440 ;
      LAYER via ;
        RECT 858.920 17.380 859.180 17.640 ;
        RECT 862.140 17.380 862.400 17.640 ;
      LAYER met2 ;
        RECT 862.200 17.670 862.340 54.000 ;
        RECT 858.920 17.350 859.180 17.670 ;
        RECT 862.140 17.350 862.400 17.670 ;
        RECT 858.980 2.400 859.120 17.350 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 876.830 15.200 877.150 15.260 ;
        RECT 882.350 15.200 882.670 15.260 ;
        RECT 876.830 15.060 882.670 15.200 ;
        RECT 876.830 15.000 877.150 15.060 ;
        RECT 882.350 15.000 882.670 15.060 ;
      LAYER via ;
        RECT 876.860 15.000 877.120 15.260 ;
        RECT 882.380 15.000 882.640 15.260 ;
      LAYER met2 ;
        RECT 882.440 15.290 882.580 54.000 ;
        RECT 876.860 14.970 877.120 15.290 ;
        RECT 882.380 14.970 882.640 15.290 ;
        RECT 876.920 2.400 877.060 14.970 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 896.700 17.410 896.840 54.000 ;
        RECT 894.860 17.270 896.840 17.410 ;
        RECT 894.860 2.400 895.000 17.270 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 912.710 17.580 913.030 17.640 ;
        RECT 917.310 17.580 917.630 17.640 ;
        RECT 912.710 17.440 917.630 17.580 ;
        RECT 912.710 17.380 913.030 17.440 ;
        RECT 917.310 17.380 917.630 17.440 ;
      LAYER via ;
        RECT 912.740 17.380 913.000 17.640 ;
        RECT 917.340 17.380 917.600 17.640 ;
      LAYER met2 ;
        RECT 917.400 17.670 917.540 54.000 ;
        RECT 912.740 17.350 913.000 17.670 ;
        RECT 917.340 17.350 917.600 17.670 ;
        RECT 912.800 2.400 912.940 17.350 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 931.200 17.410 931.340 54.000 ;
        RECT 930.280 17.270 931.340 17.410 ;
        RECT 930.280 2.400 930.420 17.270 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 948.130 17.580 948.450 17.640 ;
        RECT 951.810 17.580 952.130 17.640 ;
        RECT 948.130 17.440 952.130 17.580 ;
        RECT 948.130 17.380 948.450 17.440 ;
        RECT 951.810 17.380 952.130 17.440 ;
      LAYER via ;
        RECT 948.160 17.380 948.420 17.640 ;
        RECT 951.840 17.380 952.100 17.640 ;
      LAYER met2 ;
        RECT 951.900 17.670 952.040 54.000 ;
        RECT 948.160 17.350 948.420 17.670 ;
        RECT 951.840 17.350 952.100 17.670 ;
        RECT 948.220 2.400 948.360 17.350 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 966.070 17.580 966.390 17.640 ;
        RECT 972.510 17.580 972.830 17.640 ;
        RECT 966.070 17.440 972.830 17.580 ;
        RECT 966.070 17.380 966.390 17.440 ;
        RECT 972.510 17.380 972.830 17.440 ;
      LAYER via ;
        RECT 966.100 17.380 966.360 17.640 ;
        RECT 972.540 17.380 972.800 17.640 ;
      LAYER met2 ;
        RECT 972.600 17.670 972.740 54.000 ;
        RECT 966.100 17.350 966.360 17.670 ;
        RECT 972.540 17.350 972.800 17.670 ;
        RECT 966.160 2.400 966.300 17.350 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 984.010 17.580 984.330 17.640 ;
        RECT 986.310 17.580 986.630 17.640 ;
        RECT 984.010 17.440 986.630 17.580 ;
        RECT 984.010 17.380 984.330 17.440 ;
        RECT 986.310 17.380 986.630 17.440 ;
      LAYER via ;
        RECT 984.040 17.380 984.300 17.640 ;
        RECT 986.340 17.380 986.600 17.640 ;
      LAYER met2 ;
        RECT 986.400 17.670 986.540 54.000 ;
        RECT 984.040 17.350 984.300 17.670 ;
        RECT 986.340 17.350 986.600 17.670 ;
        RECT 984.100 2.400 984.240 17.350 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 662.930 17.240 663.250 17.300 ;
        RECT 668.450 17.240 668.770 17.300 ;
        RECT 662.930 17.100 668.770 17.240 ;
        RECT 662.930 17.040 663.250 17.100 ;
        RECT 668.450 17.040 668.770 17.100 ;
      LAYER via ;
        RECT 662.960 17.040 663.220 17.300 ;
        RECT 668.480 17.040 668.740 17.300 ;
      LAYER met2 ;
        RECT 668.540 17.330 668.680 54.000 ;
        RECT 662.960 17.010 663.220 17.330 ;
        RECT 668.480 17.010 668.740 17.330 ;
        RECT 663.020 2.400 663.160 17.010 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1001.950 17.580 1002.270 17.640 ;
        RECT 1007.010 17.580 1007.330 17.640 ;
        RECT 1001.950 17.440 1007.330 17.580 ;
        RECT 1001.950 17.380 1002.270 17.440 ;
        RECT 1007.010 17.380 1007.330 17.440 ;
      LAYER via ;
        RECT 1001.980 17.380 1002.240 17.640 ;
        RECT 1007.040 17.380 1007.300 17.640 ;
      LAYER met2 ;
        RECT 1007.100 17.670 1007.240 54.000 ;
        RECT 1001.980 17.350 1002.240 17.670 ;
        RECT 1007.040 17.350 1007.300 17.670 ;
        RECT 1002.040 2.400 1002.180 17.350 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1020.900 17.410 1021.040 54.000 ;
        RECT 1019.520 17.270 1021.040 17.410 ;
        RECT 1019.520 2.400 1019.660 17.270 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1037.370 17.580 1037.690 17.640 ;
        RECT 1041.510 17.580 1041.830 17.640 ;
        RECT 1037.370 17.440 1041.830 17.580 ;
        RECT 1037.370 17.380 1037.690 17.440 ;
        RECT 1041.510 17.380 1041.830 17.440 ;
      LAYER via ;
        RECT 1037.400 17.380 1037.660 17.640 ;
        RECT 1041.540 17.380 1041.800 17.640 ;
      LAYER met2 ;
        RECT 1041.600 17.670 1041.740 54.000 ;
        RECT 1037.400 17.350 1037.660 17.670 ;
        RECT 1041.540 17.350 1041.800 17.670 ;
        RECT 1037.460 2.400 1037.600 17.350 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1054.940 7.890 1055.080 54.000 ;
        RECT 1054.940 7.750 1055.540 7.890 ;
        RECT 1055.400 2.400 1055.540 7.750 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1073.250 17.580 1073.570 17.640 ;
        RECT 1076.010 17.580 1076.330 17.640 ;
        RECT 1073.250 17.440 1076.330 17.580 ;
        RECT 1073.250 17.380 1073.570 17.440 ;
        RECT 1076.010 17.380 1076.330 17.440 ;
      LAYER via ;
        RECT 1073.280 17.380 1073.540 17.640 ;
        RECT 1076.040 17.380 1076.300 17.640 ;
      LAYER met2 ;
        RECT 1076.100 17.670 1076.240 54.000 ;
        RECT 1073.280 17.350 1073.540 17.670 ;
        RECT 1076.040 17.350 1076.300 17.670 ;
        RECT 1073.340 2.400 1073.480 17.350 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1090.730 17.580 1091.050 17.640 ;
        RECT 1096.250 17.580 1096.570 17.640 ;
        RECT 1090.730 17.440 1096.570 17.580 ;
        RECT 1090.730 17.380 1091.050 17.440 ;
        RECT 1096.250 17.380 1096.570 17.440 ;
      LAYER via ;
        RECT 1090.760 17.380 1091.020 17.640 ;
        RECT 1096.280 17.380 1096.540 17.640 ;
      LAYER met2 ;
        RECT 1096.340 17.670 1096.480 54.000 ;
        RECT 1090.760 17.350 1091.020 17.670 ;
        RECT 1096.280 17.350 1096.540 17.670 ;
        RECT 1090.820 2.400 1090.960 17.350 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.600 17.410 1110.740 54.000 ;
        RECT 1108.760 17.270 1110.740 17.410 ;
        RECT 1108.760 2.400 1108.900 17.270 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1126.610 17.580 1126.930 17.640 ;
        RECT 1131.210 17.580 1131.530 17.640 ;
        RECT 1126.610 17.440 1131.530 17.580 ;
        RECT 1126.610 17.380 1126.930 17.440 ;
        RECT 1131.210 17.380 1131.530 17.440 ;
      LAYER via ;
        RECT 1126.640 17.380 1126.900 17.640 ;
        RECT 1131.240 17.380 1131.500 17.640 ;
      LAYER met2 ;
        RECT 1131.300 17.670 1131.440 54.000 ;
        RECT 1126.640 17.350 1126.900 17.670 ;
        RECT 1131.240 17.350 1131.500 17.670 ;
        RECT 1126.700 2.400 1126.840 17.350 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1145.100 17.410 1145.240 54.000 ;
        RECT 1144.640 17.270 1145.240 17.410 ;
        RECT 1144.640 2.400 1144.780 17.270 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1162.490 17.580 1162.810 17.640 ;
        RECT 1165.710 17.580 1166.030 17.640 ;
        RECT 1162.490 17.440 1166.030 17.580 ;
        RECT 1162.490 17.380 1162.810 17.440 ;
        RECT 1165.710 17.380 1166.030 17.440 ;
      LAYER via ;
        RECT 1162.520 17.380 1162.780 17.640 ;
        RECT 1165.740 17.380 1166.000 17.640 ;
      LAYER met2 ;
        RECT 1165.800 17.670 1165.940 54.000 ;
        RECT 1162.520 17.350 1162.780 17.670 ;
        RECT 1165.740 17.350 1166.000 17.670 ;
        RECT 1162.580 2.400 1162.720 17.350 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 680.410 17.240 680.730 17.300 ;
        RECT 682.710 17.240 683.030 17.300 ;
        RECT 680.410 17.100 683.030 17.240 ;
        RECT 680.410 17.040 680.730 17.100 ;
        RECT 682.710 17.040 683.030 17.100 ;
      LAYER via ;
        RECT 680.440 17.040 680.700 17.300 ;
        RECT 682.740 17.040 683.000 17.300 ;
      LAYER met2 ;
        RECT 682.800 17.330 682.940 54.000 ;
        RECT 680.440 17.010 680.700 17.330 ;
        RECT 682.740 17.010 683.000 17.330 ;
        RECT 680.500 2.400 680.640 17.010 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1179.970 16.220 1180.290 16.280 ;
        RECT 1186.410 16.220 1186.730 16.280 ;
        RECT 1179.970 16.080 1186.730 16.220 ;
        RECT 1179.970 16.020 1180.290 16.080 ;
        RECT 1186.410 16.020 1186.730 16.080 ;
      LAYER via ;
        RECT 1180.000 16.020 1180.260 16.280 ;
        RECT 1186.440 16.020 1186.700 16.280 ;
      LAYER met2 ;
        RECT 1186.500 16.310 1186.640 54.000 ;
        RECT 1180.000 15.990 1180.260 16.310 ;
        RECT 1186.440 15.990 1186.700 16.310 ;
        RECT 1180.060 2.400 1180.200 15.990 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1197.910 17.580 1198.230 17.640 ;
        RECT 1200.210 17.580 1200.530 17.640 ;
        RECT 1197.910 17.440 1200.530 17.580 ;
        RECT 1197.910 17.380 1198.230 17.440 ;
        RECT 1200.210 17.380 1200.530 17.440 ;
      LAYER via ;
        RECT 1197.940 17.380 1198.200 17.640 ;
        RECT 1200.240 17.380 1200.500 17.640 ;
      LAYER met2 ;
        RECT 1200.300 17.670 1200.440 54.000 ;
        RECT 1197.940 17.350 1198.200 17.670 ;
        RECT 1200.240 17.350 1200.500 17.670 ;
        RECT 1198.000 2.400 1198.140 17.350 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1215.850 17.580 1216.170 17.640 ;
        RECT 1220.910 17.580 1221.230 17.640 ;
        RECT 1215.850 17.440 1221.230 17.580 ;
        RECT 1215.850 17.380 1216.170 17.440 ;
        RECT 1220.910 17.380 1221.230 17.440 ;
      LAYER via ;
        RECT 1215.880 17.380 1216.140 17.640 ;
        RECT 1220.940 17.380 1221.200 17.640 ;
      LAYER met2 ;
        RECT 1221.000 17.670 1221.140 54.000 ;
        RECT 1215.880 17.350 1216.140 17.670 ;
        RECT 1220.940 17.350 1221.200 17.670 ;
        RECT 1215.940 2.400 1216.080 17.350 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1234.800 17.410 1234.940 54.000 ;
        RECT 1233.880 17.270 1234.940 17.410 ;
        RECT 1233.880 2.400 1234.020 17.270 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1251.730 17.240 1252.050 17.300 ;
        RECT 1255.410 17.240 1255.730 17.300 ;
        RECT 1251.730 17.100 1255.730 17.240 ;
        RECT 1251.730 17.040 1252.050 17.100 ;
        RECT 1255.410 17.040 1255.730 17.100 ;
      LAYER via ;
        RECT 1251.760 17.040 1252.020 17.300 ;
        RECT 1255.440 17.040 1255.700 17.300 ;
      LAYER met2 ;
        RECT 1255.500 17.330 1255.640 54.000 ;
        RECT 1251.760 17.010 1252.020 17.330 ;
        RECT 1255.440 17.010 1255.700 17.330 ;
        RECT 1251.820 2.400 1251.960 17.010 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1268.840 17.410 1268.980 54.000 ;
        RECT 1268.840 17.270 1269.440 17.410 ;
        RECT 1269.300 2.400 1269.440 17.270 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1287.150 17.580 1287.470 17.640 ;
        RECT 1289.910 17.580 1290.230 17.640 ;
        RECT 1287.150 17.440 1290.230 17.580 ;
        RECT 1287.150 17.380 1287.470 17.440 ;
        RECT 1289.910 17.380 1290.230 17.440 ;
      LAYER via ;
        RECT 1287.180 17.380 1287.440 17.640 ;
        RECT 1289.940 17.380 1290.200 17.640 ;
      LAYER met2 ;
        RECT 1290.000 17.670 1290.140 54.000 ;
        RECT 1287.180 17.350 1287.440 17.670 ;
        RECT 1289.940 17.350 1290.200 17.670 ;
        RECT 1287.240 2.400 1287.380 17.350 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1305.090 15.200 1305.410 15.260 ;
        RECT 1310.610 15.200 1310.930 15.260 ;
        RECT 1305.090 15.060 1310.930 15.200 ;
        RECT 1305.090 15.000 1305.410 15.060 ;
        RECT 1310.610 15.000 1310.930 15.060 ;
      LAYER via ;
        RECT 1305.120 15.000 1305.380 15.260 ;
        RECT 1310.640 15.000 1310.900 15.260 ;
      LAYER met2 ;
        RECT 1310.700 15.290 1310.840 54.000 ;
        RECT 1305.120 14.970 1305.380 15.290 ;
        RECT 1310.640 14.970 1310.900 15.290 ;
        RECT 1305.180 2.400 1305.320 14.970 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1324.500 17.410 1324.640 54.000 ;
        RECT 1323.120 17.270 1324.640 17.410 ;
        RECT 1323.120 2.400 1323.260 17.270 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1340.510 17.580 1340.830 17.640 ;
        RECT 1345.110 17.580 1345.430 17.640 ;
        RECT 1340.510 17.440 1345.430 17.580 ;
        RECT 1340.510 17.380 1340.830 17.440 ;
        RECT 1345.110 17.380 1345.430 17.440 ;
      LAYER via ;
        RECT 1340.540 17.380 1340.800 17.640 ;
        RECT 1345.140 17.380 1345.400 17.640 ;
      LAYER met2 ;
        RECT 1345.200 17.670 1345.340 54.000 ;
        RECT 1340.540 17.350 1340.800 17.670 ;
        RECT 1345.140 17.350 1345.400 17.670 ;
        RECT 1340.600 2.400 1340.740 17.350 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 698.350 17.240 698.670 17.300 ;
        RECT 703.410 17.240 703.730 17.300 ;
        RECT 698.350 17.100 703.730 17.240 ;
        RECT 698.350 17.040 698.670 17.100 ;
        RECT 703.410 17.040 703.730 17.100 ;
      LAYER via ;
        RECT 698.380 17.040 698.640 17.300 ;
        RECT 703.440 17.040 703.700 17.300 ;
      LAYER met2 ;
        RECT 703.500 17.330 703.640 54.000 ;
        RECT 698.380 17.010 698.640 17.330 ;
        RECT 703.440 17.010 703.700 17.330 ;
        RECT 698.440 2.400 698.580 17.010 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1359.460 17.410 1359.600 54.000 ;
        RECT 1358.540 17.270 1359.600 17.410 ;
        RECT 1358.540 2.400 1358.680 17.270 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1374.090 16.220 1374.410 16.280 ;
        RECT 1376.390 16.220 1376.710 16.280 ;
        RECT 1374.090 16.080 1376.710 16.220 ;
        RECT 1374.090 16.020 1374.410 16.080 ;
        RECT 1376.390 16.020 1376.710 16.080 ;
      LAYER via ;
        RECT 1374.120 16.020 1374.380 16.280 ;
        RECT 1376.420 16.020 1376.680 16.280 ;
      LAYER met2 ;
        RECT 1374.180 16.310 1374.320 54.000 ;
        RECT 1374.120 15.990 1374.380 16.310 ;
        RECT 1376.420 15.990 1376.680 16.310 ;
        RECT 1376.480 2.400 1376.620 15.990 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1393.960 17.410 1394.100 54.000 ;
        RECT 1393.960 17.270 1394.560 17.410 ;
        RECT 1394.420 2.400 1394.560 17.270 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1407.670 17.580 1407.990 17.640 ;
        RECT 1412.270 17.580 1412.590 17.640 ;
        RECT 1407.670 17.440 1412.590 17.580 ;
        RECT 1407.670 17.380 1407.990 17.440 ;
        RECT 1412.270 17.380 1412.590 17.440 ;
      LAYER via ;
        RECT 1407.700 17.380 1407.960 17.640 ;
        RECT 1412.300 17.380 1412.560 17.640 ;
      LAYER met2 ;
        RECT 1407.760 17.670 1407.900 54.000 ;
        RECT 1407.700 17.350 1407.960 17.670 ;
        RECT 1412.300 17.350 1412.560 17.670 ;
        RECT 1412.360 2.400 1412.500 17.350 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1428.000 17.410 1428.140 54.000 ;
        RECT 1428.000 17.270 1429.980 17.410 ;
        RECT 1429.840 2.400 1429.980 17.270 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1442.260 17.410 1442.400 54.000 ;
        RECT 1442.260 17.270 1447.920 17.410 ;
        RECT 1447.780 2.400 1447.920 17.270 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1455.050 14.860 1455.370 14.920 ;
        RECT 1465.630 14.860 1465.950 14.920 ;
        RECT 1455.050 14.720 1465.950 14.860 ;
        RECT 1455.050 14.660 1455.370 14.720 ;
        RECT 1465.630 14.660 1465.950 14.720 ;
      LAYER via ;
        RECT 1455.080 14.660 1455.340 14.920 ;
        RECT 1465.660 14.660 1465.920 14.920 ;
      LAYER met2 ;
        RECT 1455.140 14.950 1455.280 54.000 ;
        RECT 1455.080 14.630 1455.340 14.950 ;
        RECT 1465.660 14.630 1465.920 14.950 ;
        RECT 1465.720 2.400 1465.860 14.630 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1475.750 20.300 1476.070 20.360 ;
        RECT 1483.570 20.300 1483.890 20.360 ;
        RECT 1475.750 20.160 1483.890 20.300 ;
        RECT 1475.750 20.100 1476.070 20.160 ;
        RECT 1483.570 20.100 1483.890 20.160 ;
      LAYER via ;
        RECT 1475.780 20.100 1476.040 20.360 ;
        RECT 1483.600 20.100 1483.860 20.360 ;
      LAYER met2 ;
        RECT 1475.840 20.390 1475.980 54.000 ;
        RECT 1475.780 20.070 1476.040 20.390 ;
        RECT 1483.600 20.070 1483.860 20.390 ;
        RECT 1483.660 2.400 1483.800 20.070 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1490.010 17.580 1490.330 17.640 ;
        RECT 1501.510 17.580 1501.830 17.640 ;
        RECT 1490.010 17.440 1501.830 17.580 ;
        RECT 1490.010 17.380 1490.330 17.440 ;
        RECT 1501.510 17.380 1501.830 17.440 ;
      LAYER via ;
        RECT 1490.040 17.380 1490.300 17.640 ;
        RECT 1501.540 17.380 1501.800 17.640 ;
      LAYER met2 ;
        RECT 1490.100 17.670 1490.240 54.000 ;
        RECT 1490.040 17.350 1490.300 17.670 ;
        RECT 1501.540 17.350 1501.800 17.670 ;
        RECT 1501.600 2.400 1501.740 17.350 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1503.810 17.240 1504.130 17.300 ;
        RECT 1518.990 17.240 1519.310 17.300 ;
        RECT 1503.810 17.100 1519.310 17.240 ;
        RECT 1503.810 17.040 1504.130 17.100 ;
        RECT 1518.990 17.040 1519.310 17.100 ;
      LAYER via ;
        RECT 1503.840 17.040 1504.100 17.300 ;
        RECT 1519.020 17.040 1519.280 17.300 ;
      LAYER met2 ;
        RECT 1503.900 17.330 1504.040 54.000 ;
        RECT 1503.840 17.010 1504.100 17.330 ;
        RECT 1519.020 17.010 1519.280 17.330 ;
        RECT 1519.080 2.400 1519.220 17.010 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 717.300 16.730 717.440 54.000 ;
        RECT 716.380 16.590 717.440 16.730 ;
        RECT 716.380 2.400 716.520 16.590 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1517.150 17.920 1517.470 17.980 ;
        RECT 1536.930 17.920 1537.250 17.980 ;
        RECT 1517.150 17.780 1537.250 17.920 ;
        RECT 1517.150 17.720 1517.470 17.780 ;
        RECT 1536.930 17.720 1537.250 17.780 ;
      LAYER via ;
        RECT 1517.180 17.720 1517.440 17.980 ;
        RECT 1536.960 17.720 1537.220 17.980 ;
      LAYER met2 ;
        RECT 1517.240 18.010 1517.380 54.000 ;
        RECT 1517.180 17.690 1517.440 18.010 ;
        RECT 1536.960 17.690 1537.220 18.010 ;
        RECT 1537.020 2.400 1537.160 17.690 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1530.950 17.240 1531.270 17.300 ;
        RECT 1554.870 17.240 1555.190 17.300 ;
        RECT 1530.950 17.100 1555.190 17.240 ;
        RECT 1530.950 17.040 1531.270 17.100 ;
        RECT 1554.870 17.040 1555.190 17.100 ;
      LAYER via ;
        RECT 1530.980 17.040 1531.240 17.300 ;
        RECT 1554.900 17.040 1555.160 17.300 ;
      LAYER met2 ;
        RECT 1531.040 17.330 1531.180 54.000 ;
        RECT 1530.980 17.010 1531.240 17.330 ;
        RECT 1554.900 17.010 1555.160 17.330 ;
        RECT 1554.960 2.400 1555.100 17.010 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1552.110 16.560 1552.430 16.620 ;
        RECT 1572.810 16.560 1573.130 16.620 ;
        RECT 1552.110 16.420 1573.130 16.560 ;
        RECT 1552.110 16.360 1552.430 16.420 ;
        RECT 1572.810 16.360 1573.130 16.420 ;
      LAYER via ;
        RECT 1552.140 16.360 1552.400 16.620 ;
        RECT 1572.840 16.360 1573.100 16.620 ;
      LAYER met2 ;
        RECT 1552.200 16.650 1552.340 54.000 ;
        RECT 1552.140 16.330 1552.400 16.650 ;
        RECT 1572.840 16.330 1573.100 16.650 ;
        RECT 1572.900 2.400 1573.040 16.330 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1565.910 19.280 1566.230 19.340 ;
        RECT 1590.290 19.280 1590.610 19.340 ;
        RECT 1565.910 19.140 1590.610 19.280 ;
        RECT 1565.910 19.080 1566.230 19.140 ;
        RECT 1590.290 19.080 1590.610 19.140 ;
      LAYER via ;
        RECT 1565.940 19.080 1566.200 19.340 ;
        RECT 1590.320 19.080 1590.580 19.340 ;
      LAYER met2 ;
        RECT 1566.000 19.370 1566.140 54.000 ;
        RECT 1565.940 19.050 1566.200 19.370 ;
        RECT 1590.320 19.050 1590.580 19.370 ;
        RECT 1590.380 2.400 1590.520 19.050 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1579.710 17.240 1580.030 17.300 ;
        RECT 1608.230 17.240 1608.550 17.300 ;
        RECT 1579.710 17.100 1608.550 17.240 ;
        RECT 1579.710 17.040 1580.030 17.100 ;
        RECT 1608.230 17.040 1608.550 17.100 ;
      LAYER via ;
        RECT 1579.740 17.040 1580.000 17.300 ;
        RECT 1608.260 17.040 1608.520 17.300 ;
      LAYER met2 ;
        RECT 1579.800 17.330 1579.940 54.000 ;
        RECT 1579.740 17.010 1580.000 17.330 ;
        RECT 1608.260 17.010 1608.520 17.330 ;
        RECT 1608.320 2.400 1608.460 17.010 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1593.050 16.900 1593.370 16.960 ;
        RECT 1626.170 16.900 1626.490 16.960 ;
        RECT 1593.050 16.760 1626.490 16.900 ;
        RECT 1593.050 16.700 1593.370 16.760 ;
        RECT 1626.170 16.700 1626.490 16.760 ;
      LAYER via ;
        RECT 1593.080 16.700 1593.340 16.960 ;
        RECT 1626.200 16.700 1626.460 16.960 ;
      LAYER met2 ;
        RECT 1593.140 16.990 1593.280 54.000 ;
        RECT 1593.080 16.670 1593.340 16.990 ;
        RECT 1626.200 16.670 1626.460 16.990 ;
        RECT 1626.260 2.400 1626.400 16.670 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1614.210 18.260 1614.530 18.320 ;
        RECT 1644.110 18.260 1644.430 18.320 ;
        RECT 1614.210 18.120 1644.430 18.260 ;
        RECT 1614.210 18.060 1614.530 18.120 ;
        RECT 1644.110 18.060 1644.430 18.120 ;
      LAYER via ;
        RECT 1614.240 18.060 1614.500 18.320 ;
        RECT 1644.140 18.060 1644.400 18.320 ;
      LAYER met2 ;
        RECT 1614.300 18.350 1614.440 54.000 ;
        RECT 1614.240 18.030 1614.500 18.350 ;
        RECT 1644.140 18.030 1644.400 18.350 ;
        RECT 1644.200 2.400 1644.340 18.030 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1628.010 19.620 1628.330 19.680 ;
        RECT 1662.050 19.620 1662.370 19.680 ;
        RECT 1628.010 19.480 1662.370 19.620 ;
        RECT 1628.010 19.420 1628.330 19.480 ;
        RECT 1662.050 19.420 1662.370 19.480 ;
      LAYER via ;
        RECT 1628.040 19.420 1628.300 19.680 ;
        RECT 1662.080 19.420 1662.340 19.680 ;
      LAYER met2 ;
        RECT 1628.100 19.710 1628.240 54.000 ;
        RECT 1628.040 19.390 1628.300 19.710 ;
        RECT 1662.080 19.390 1662.340 19.710 ;
        RECT 1662.140 2.400 1662.280 19.390 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1641.810 18.940 1642.130 19.000 ;
        RECT 1679.530 18.940 1679.850 19.000 ;
        RECT 1641.810 18.800 1679.850 18.940 ;
        RECT 1641.810 18.740 1642.130 18.800 ;
        RECT 1679.530 18.740 1679.850 18.800 ;
      LAYER via ;
        RECT 1641.840 18.740 1642.100 19.000 ;
        RECT 1679.560 18.740 1679.820 19.000 ;
      LAYER met2 ;
        RECT 1641.900 19.030 1642.040 54.000 ;
        RECT 1641.840 18.710 1642.100 19.030 ;
        RECT 1679.560 18.710 1679.820 19.030 ;
        RECT 1679.620 2.400 1679.760 18.710 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1655.150 17.580 1655.470 17.640 ;
        RECT 1697.470 17.580 1697.790 17.640 ;
        RECT 1655.150 17.440 1697.790 17.580 ;
        RECT 1655.150 17.380 1655.470 17.440 ;
        RECT 1697.470 17.380 1697.790 17.440 ;
      LAYER via ;
        RECT 1655.180 17.380 1655.440 17.640 ;
        RECT 1697.500 17.380 1697.760 17.640 ;
      LAYER met2 ;
        RECT 1655.240 17.670 1655.380 54.000 ;
        RECT 1655.180 17.350 1655.440 17.670 ;
        RECT 1697.500 17.350 1697.760 17.670 ;
        RECT 1697.560 2.400 1697.700 17.350 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 734.230 17.580 734.550 17.640 ;
        RECT 737.910 17.580 738.230 17.640 ;
        RECT 734.230 17.440 738.230 17.580 ;
        RECT 734.230 17.380 734.550 17.440 ;
        RECT 737.910 17.380 738.230 17.440 ;
      LAYER via ;
        RECT 734.260 17.380 734.520 17.640 ;
        RECT 737.940 17.380 738.200 17.640 ;
      LAYER met2 ;
        RECT 738.000 17.670 738.140 54.000 ;
        RECT 734.260 17.350 734.520 17.670 ;
        RECT 737.940 17.350 738.200 17.670 ;
        RECT 734.320 2.400 734.460 17.350 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1668.950 17.920 1669.270 17.980 ;
        RECT 1715.410 17.920 1715.730 17.980 ;
        RECT 1668.950 17.780 1715.730 17.920 ;
        RECT 1668.950 17.720 1669.270 17.780 ;
        RECT 1715.410 17.720 1715.730 17.780 ;
      LAYER via ;
        RECT 1668.980 17.720 1669.240 17.980 ;
        RECT 1715.440 17.720 1715.700 17.980 ;
      LAYER met2 ;
        RECT 1669.040 18.010 1669.180 54.000 ;
        RECT 1668.980 17.690 1669.240 18.010 ;
        RECT 1715.440 17.690 1715.700 18.010 ;
        RECT 1715.500 2.400 1715.640 17.690 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1689.650 18.600 1689.970 18.660 ;
        RECT 1733.350 18.600 1733.670 18.660 ;
        RECT 1689.650 18.460 1733.670 18.600 ;
        RECT 1689.650 18.400 1689.970 18.460 ;
        RECT 1733.350 18.400 1733.670 18.460 ;
      LAYER via ;
        RECT 1689.680 18.400 1689.940 18.660 ;
        RECT 1733.380 18.400 1733.640 18.660 ;
      LAYER met2 ;
        RECT 1689.740 18.690 1689.880 54.000 ;
        RECT 1689.680 18.370 1689.940 18.690 ;
        RECT 1733.380 18.370 1733.640 18.690 ;
        RECT 1733.440 2.400 1733.580 18.370 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.910 20.300 1704.230 20.360 ;
        RECT 1751.290 20.300 1751.610 20.360 ;
        RECT 1703.910 20.160 1751.610 20.300 ;
        RECT 1703.910 20.100 1704.230 20.160 ;
        RECT 1751.290 20.100 1751.610 20.160 ;
      LAYER via ;
        RECT 1703.940 20.100 1704.200 20.360 ;
        RECT 1751.320 20.100 1751.580 20.360 ;
      LAYER met2 ;
        RECT 1704.000 20.390 1704.140 54.000 ;
        RECT 1703.940 20.070 1704.200 20.390 ;
        RECT 1751.320 20.070 1751.580 20.390 ;
        RECT 1751.380 2.400 1751.520 20.070 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1717.710 18.260 1718.030 18.320 ;
        RECT 1768.770 18.260 1769.090 18.320 ;
        RECT 1717.710 18.120 1769.090 18.260 ;
        RECT 1717.710 18.060 1718.030 18.120 ;
        RECT 1768.770 18.060 1769.090 18.120 ;
      LAYER via ;
        RECT 1717.740 18.060 1718.000 18.320 ;
        RECT 1768.800 18.060 1769.060 18.320 ;
      LAYER met2 ;
        RECT 1717.800 18.350 1717.940 54.000 ;
        RECT 1717.740 18.030 1718.000 18.350 ;
        RECT 1768.800 18.030 1769.060 18.350 ;
        RECT 1768.860 2.400 1769.000 18.030 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1731.050 17.580 1731.370 17.640 ;
        RECT 1786.710 17.580 1787.030 17.640 ;
        RECT 1731.050 17.440 1787.030 17.580 ;
        RECT 1731.050 17.380 1731.370 17.440 ;
        RECT 1786.710 17.380 1787.030 17.440 ;
      LAYER via ;
        RECT 1731.080 17.380 1731.340 17.640 ;
        RECT 1786.740 17.380 1787.000 17.640 ;
      LAYER met2 ;
        RECT 1731.140 17.670 1731.280 54.000 ;
        RECT 1731.080 17.350 1731.340 17.670 ;
        RECT 1786.740 17.350 1787.000 17.670 ;
        RECT 1786.800 2.400 1786.940 17.350 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1751.750 18.600 1752.070 18.660 ;
        RECT 1804.650 18.600 1804.970 18.660 ;
        RECT 1751.750 18.460 1804.970 18.600 ;
        RECT 1751.750 18.400 1752.070 18.460 ;
        RECT 1804.650 18.400 1804.970 18.460 ;
      LAYER via ;
        RECT 1751.780 18.400 1752.040 18.660 ;
        RECT 1804.680 18.400 1804.940 18.660 ;
      LAYER met2 ;
        RECT 1751.840 18.690 1751.980 54.000 ;
        RECT 1751.780 18.370 1752.040 18.690 ;
        RECT 1804.680 18.370 1804.940 18.690 ;
        RECT 1804.740 2.400 1804.880 18.370 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1766.010 19.280 1766.330 19.340 ;
        RECT 1822.590 19.280 1822.910 19.340 ;
        RECT 1766.010 19.140 1822.910 19.280 ;
        RECT 1766.010 19.080 1766.330 19.140 ;
        RECT 1822.590 19.080 1822.910 19.140 ;
      LAYER via ;
        RECT 1766.040 19.080 1766.300 19.340 ;
        RECT 1822.620 19.080 1822.880 19.340 ;
      LAYER met2 ;
        RECT 1766.100 19.370 1766.240 54.000 ;
        RECT 1766.040 19.050 1766.300 19.370 ;
        RECT 1822.620 19.050 1822.880 19.370 ;
        RECT 1822.680 2.400 1822.820 19.050 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1779.810 16.900 1780.130 16.960 ;
        RECT 1840.070 16.900 1840.390 16.960 ;
        RECT 1779.810 16.760 1840.390 16.900 ;
        RECT 1779.810 16.700 1780.130 16.760 ;
        RECT 1840.070 16.700 1840.390 16.760 ;
      LAYER via ;
        RECT 1779.840 16.700 1780.100 16.960 ;
        RECT 1840.100 16.700 1840.360 16.960 ;
      LAYER met2 ;
        RECT 1779.900 16.990 1780.040 54.000 ;
        RECT 1779.840 16.670 1780.100 16.990 ;
        RECT 1840.100 16.670 1840.360 16.990 ;
        RECT 1840.160 2.400 1840.300 16.670 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1793.610 17.580 1793.930 17.640 ;
        RECT 1858.010 17.580 1858.330 17.640 ;
        RECT 1793.610 17.440 1858.330 17.580 ;
        RECT 1793.610 17.380 1793.930 17.440 ;
        RECT 1858.010 17.380 1858.330 17.440 ;
      LAYER via ;
        RECT 1793.640 17.380 1793.900 17.640 ;
        RECT 1858.040 17.380 1858.300 17.640 ;
      LAYER met2 ;
        RECT 1793.700 17.670 1793.840 54.000 ;
        RECT 1793.640 17.350 1793.900 17.670 ;
        RECT 1858.040 17.350 1858.300 17.670 ;
        RECT 1858.100 2.400 1858.240 17.350 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1806.950 18.600 1807.270 18.660 ;
        RECT 1875.950 18.600 1876.270 18.660 ;
        RECT 1806.950 18.460 1876.270 18.600 ;
        RECT 1806.950 18.400 1807.270 18.460 ;
        RECT 1875.950 18.400 1876.270 18.460 ;
      LAYER via ;
        RECT 1806.980 18.400 1807.240 18.660 ;
        RECT 1875.980 18.400 1876.240 18.660 ;
      LAYER met2 ;
        RECT 1807.040 18.690 1807.180 54.000 ;
        RECT 1806.980 18.370 1807.240 18.690 ;
        RECT 1875.980 18.370 1876.240 18.690 ;
        RECT 1876.040 2.400 1876.180 18.370 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 752.170 17.580 752.490 17.640 ;
        RECT 758.610 17.580 758.930 17.640 ;
        RECT 752.170 17.440 758.930 17.580 ;
        RECT 752.170 17.380 752.490 17.440 ;
        RECT 758.610 17.380 758.930 17.440 ;
      LAYER via ;
        RECT 752.200 17.380 752.460 17.640 ;
        RECT 758.640 17.380 758.900 17.640 ;
      LAYER met2 ;
        RECT 758.700 17.670 758.840 54.000 ;
        RECT 752.200 17.350 752.460 17.670 ;
        RECT 758.640 17.350 758.900 17.670 ;
        RECT 752.260 2.400 752.400 17.350 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1827.650 19.280 1827.970 19.340 ;
        RECT 1893.890 19.280 1894.210 19.340 ;
        RECT 1827.650 19.140 1894.210 19.280 ;
        RECT 1827.650 19.080 1827.970 19.140 ;
        RECT 1893.890 19.080 1894.210 19.140 ;
      LAYER via ;
        RECT 1827.680 19.080 1827.940 19.340 ;
        RECT 1893.920 19.080 1894.180 19.340 ;
      LAYER met2 ;
        RECT 1827.740 19.370 1827.880 54.000 ;
        RECT 1827.680 19.050 1827.940 19.370 ;
        RECT 1893.920 19.050 1894.180 19.370 ;
        RECT 1893.980 2.400 1894.120 19.050 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1841.910 18.260 1842.230 18.320 ;
        RECT 1911.830 18.260 1912.150 18.320 ;
        RECT 1841.910 18.120 1912.150 18.260 ;
        RECT 1841.910 18.060 1842.230 18.120 ;
        RECT 1911.830 18.060 1912.150 18.120 ;
      LAYER via ;
        RECT 1841.940 18.060 1842.200 18.320 ;
        RECT 1911.860 18.060 1912.120 18.320 ;
      LAYER met2 ;
        RECT 1842.000 18.350 1842.140 54.000 ;
        RECT 1841.940 18.030 1842.200 18.350 ;
        RECT 1911.860 18.030 1912.120 18.350 ;
        RECT 1911.920 2.400 1912.060 18.030 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1855.710 18.940 1856.030 19.000 ;
        RECT 1929.310 18.940 1929.630 19.000 ;
        RECT 1855.710 18.800 1929.630 18.940 ;
        RECT 1855.710 18.740 1856.030 18.800 ;
        RECT 1929.310 18.740 1929.630 18.800 ;
      LAYER via ;
        RECT 1855.740 18.740 1856.000 19.000 ;
        RECT 1929.340 18.740 1929.600 19.000 ;
      LAYER met2 ;
        RECT 1855.800 19.030 1855.940 54.000 ;
        RECT 1855.740 18.710 1856.000 19.030 ;
        RECT 1929.340 18.710 1929.600 19.030 ;
        RECT 1929.400 2.400 1929.540 18.710 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1869.050 17.580 1869.370 17.640 ;
        RECT 1947.250 17.580 1947.570 17.640 ;
        RECT 1869.050 17.440 1947.570 17.580 ;
        RECT 1869.050 17.380 1869.370 17.440 ;
        RECT 1947.250 17.380 1947.570 17.440 ;
      LAYER via ;
        RECT 1869.080 17.380 1869.340 17.640 ;
        RECT 1947.280 17.380 1947.540 17.640 ;
      LAYER met2 ;
        RECT 1869.140 17.670 1869.280 54.000 ;
        RECT 1869.080 17.350 1869.340 17.670 ;
        RECT 1947.280 17.350 1947.540 17.670 ;
        RECT 1947.340 2.400 1947.480 17.350 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1889.750 20.640 1890.070 20.700 ;
        RECT 1965.190 20.640 1965.510 20.700 ;
        RECT 1889.750 20.500 1965.510 20.640 ;
        RECT 1889.750 20.440 1890.070 20.500 ;
        RECT 1965.190 20.440 1965.510 20.500 ;
      LAYER via ;
        RECT 1889.780 20.440 1890.040 20.700 ;
        RECT 1965.220 20.440 1965.480 20.700 ;
      LAYER met2 ;
        RECT 1889.840 20.730 1889.980 54.000 ;
        RECT 1889.780 20.410 1890.040 20.730 ;
        RECT 1965.220 20.410 1965.480 20.730 ;
        RECT 1965.280 2.400 1965.420 20.410 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1904.010 15.880 1904.330 15.940 ;
        RECT 1983.130 15.880 1983.450 15.940 ;
        RECT 1904.010 15.740 1983.450 15.880 ;
        RECT 1904.010 15.680 1904.330 15.740 ;
        RECT 1983.130 15.680 1983.450 15.740 ;
      LAYER via ;
        RECT 1904.040 15.680 1904.300 15.940 ;
        RECT 1983.160 15.680 1983.420 15.940 ;
      LAYER met2 ;
        RECT 1904.100 15.970 1904.240 54.000 ;
        RECT 1904.040 15.650 1904.300 15.970 ;
        RECT 1983.160 15.650 1983.420 15.970 ;
        RECT 1983.220 2.400 1983.360 15.650 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1917.810 18.260 1918.130 18.320 ;
        RECT 2001.070 18.260 2001.390 18.320 ;
        RECT 1917.810 18.120 2001.390 18.260 ;
        RECT 1917.810 18.060 1918.130 18.120 ;
        RECT 2001.070 18.060 2001.390 18.120 ;
      LAYER via ;
        RECT 1917.840 18.060 1918.100 18.320 ;
        RECT 2001.100 18.060 2001.360 18.320 ;
      LAYER met2 ;
        RECT 1917.900 18.350 1918.040 54.000 ;
        RECT 1917.840 18.030 1918.100 18.350 ;
        RECT 2001.100 18.030 2001.360 18.350 ;
        RECT 2001.160 2.400 2001.300 18.030 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1931.610 16.220 1931.930 16.280 ;
        RECT 2018.550 16.220 2018.870 16.280 ;
        RECT 1931.610 16.080 2018.870 16.220 ;
        RECT 1931.610 16.020 1931.930 16.080 ;
        RECT 2018.550 16.020 2018.870 16.080 ;
      LAYER via ;
        RECT 1931.640 16.020 1931.900 16.280 ;
        RECT 2018.580 16.020 2018.840 16.280 ;
      LAYER met2 ;
        RECT 1931.700 16.310 1931.840 54.000 ;
        RECT 1931.640 15.990 1931.900 16.310 ;
        RECT 2018.580 15.990 2018.840 16.310 ;
        RECT 2018.640 2.400 2018.780 15.990 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1944.950 17.920 1945.270 17.980 ;
        RECT 2036.490 17.920 2036.810 17.980 ;
        RECT 1944.950 17.780 2036.810 17.920 ;
        RECT 1944.950 17.720 1945.270 17.780 ;
        RECT 2036.490 17.720 2036.810 17.780 ;
      LAYER via ;
        RECT 1944.980 17.720 1945.240 17.980 ;
        RECT 2036.520 17.720 2036.780 17.980 ;
      LAYER met2 ;
        RECT 1945.040 18.010 1945.180 54.000 ;
        RECT 1944.980 17.690 1945.240 18.010 ;
        RECT 2036.520 17.690 2036.780 18.010 ;
        RECT 2036.580 2.400 2036.720 17.690 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1966.110 15.540 1966.430 15.600 ;
        RECT 2054.430 15.540 2054.750 15.600 ;
        RECT 1966.110 15.400 2054.750 15.540 ;
        RECT 1966.110 15.340 1966.430 15.400 ;
        RECT 2054.430 15.340 2054.750 15.400 ;
      LAYER via ;
        RECT 1966.140 15.340 1966.400 15.600 ;
        RECT 2054.460 15.340 2054.720 15.600 ;
      LAYER met2 ;
        RECT 1966.200 15.630 1966.340 54.000 ;
        RECT 1966.140 15.310 1966.400 15.630 ;
        RECT 2054.460 15.310 2054.720 15.630 ;
        RECT 2054.520 2.400 2054.660 15.310 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 769.650 17.580 769.970 17.640 ;
        RECT 772.410 17.580 772.730 17.640 ;
        RECT 769.650 17.440 772.730 17.580 ;
        RECT 769.650 17.380 769.970 17.440 ;
        RECT 772.410 17.380 772.730 17.440 ;
      LAYER via ;
        RECT 769.680 17.380 769.940 17.640 ;
        RECT 772.440 17.380 772.700 17.640 ;
      LAYER met2 ;
        RECT 772.500 17.670 772.640 54.000 ;
        RECT 769.680 17.350 769.940 17.670 ;
        RECT 772.440 17.350 772.700 17.670 ;
        RECT 769.740 2.400 769.880 17.350 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1979.910 20.640 1980.230 20.700 ;
        RECT 2072.370 20.640 2072.690 20.700 ;
        RECT 1979.910 20.500 2072.690 20.640 ;
        RECT 1979.910 20.440 1980.230 20.500 ;
        RECT 2072.370 20.440 2072.690 20.500 ;
      LAYER via ;
        RECT 1979.940 20.440 1980.200 20.700 ;
        RECT 2072.400 20.440 2072.660 20.700 ;
      LAYER met2 ;
        RECT 1980.000 20.730 1980.140 54.000 ;
        RECT 1979.940 20.410 1980.200 20.730 ;
        RECT 2072.400 20.410 2072.660 20.730 ;
        RECT 2072.460 2.400 2072.600 20.410 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1993.710 15.880 1994.030 15.940 ;
        RECT 2089.850 15.880 2090.170 15.940 ;
        RECT 1993.710 15.740 2090.170 15.880 ;
        RECT 1993.710 15.680 1994.030 15.740 ;
        RECT 2089.850 15.680 2090.170 15.740 ;
      LAYER via ;
        RECT 1993.740 15.680 1994.000 15.940 ;
        RECT 2089.880 15.680 2090.140 15.940 ;
      LAYER met2 ;
        RECT 1993.800 15.970 1993.940 54.000 ;
        RECT 1993.740 15.650 1994.000 15.970 ;
        RECT 2089.880 15.650 2090.140 15.970 ;
        RECT 2089.940 2.400 2090.080 15.650 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2007.510 18.260 2007.830 18.320 ;
        RECT 2107.790 18.260 2108.110 18.320 ;
        RECT 2007.510 18.120 2108.110 18.260 ;
        RECT 2007.510 18.060 2007.830 18.120 ;
        RECT 2107.790 18.060 2108.110 18.120 ;
      LAYER via ;
        RECT 2007.540 18.060 2007.800 18.320 ;
        RECT 2107.820 18.060 2108.080 18.320 ;
      LAYER met2 ;
        RECT 2007.600 18.350 2007.740 54.000 ;
        RECT 2007.540 18.030 2007.800 18.350 ;
        RECT 2107.820 18.030 2108.080 18.350 ;
        RECT 2107.880 2.400 2108.020 18.030 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2020.850 17.240 2021.170 17.300 ;
        RECT 2125.270 17.240 2125.590 17.300 ;
        RECT 2020.850 17.100 2125.590 17.240 ;
        RECT 2020.850 17.040 2021.170 17.100 ;
        RECT 2125.270 17.040 2125.590 17.100 ;
      LAYER via ;
        RECT 2020.880 17.040 2021.140 17.300 ;
        RECT 2125.300 17.040 2125.560 17.300 ;
      LAYER met2 ;
        RECT 2020.940 17.330 2021.080 54.000 ;
        RECT 2020.880 17.010 2021.140 17.330 ;
        RECT 2125.300 17.010 2125.560 17.330 ;
        RECT 2125.360 16.730 2125.500 17.010 ;
        RECT 2125.360 16.590 2125.960 16.730 ;
        RECT 2125.820 2.400 2125.960 16.590 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2042.010 18.940 2042.330 19.000 ;
        RECT 2143.670 18.940 2143.990 19.000 ;
        RECT 2042.010 18.800 2143.990 18.940 ;
        RECT 2042.010 18.740 2042.330 18.800 ;
        RECT 2143.670 18.740 2143.990 18.800 ;
      LAYER via ;
        RECT 2042.040 18.740 2042.300 19.000 ;
        RECT 2143.700 18.740 2143.960 19.000 ;
      LAYER met2 ;
        RECT 2042.100 19.030 2042.240 54.000 ;
        RECT 2042.040 18.710 2042.300 19.030 ;
        RECT 2143.700 18.710 2143.960 19.030 ;
        RECT 2143.760 2.400 2143.900 18.710 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2055.810 19.960 2056.130 20.020 ;
        RECT 2161.610 19.960 2161.930 20.020 ;
        RECT 2055.810 19.820 2161.930 19.960 ;
        RECT 2055.810 19.760 2056.130 19.820 ;
        RECT 2161.610 19.760 2161.930 19.820 ;
      LAYER via ;
        RECT 2055.840 19.760 2056.100 20.020 ;
        RECT 2161.640 19.760 2161.900 20.020 ;
      LAYER met2 ;
        RECT 2055.900 20.050 2056.040 54.000 ;
        RECT 2055.840 19.730 2056.100 20.050 ;
        RECT 2161.640 19.730 2161.900 20.050 ;
        RECT 2161.700 2.400 2161.840 19.730 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2069.610 18.600 2069.930 18.660 ;
        RECT 2179.090 18.600 2179.410 18.660 ;
        RECT 2069.610 18.460 2179.410 18.600 ;
        RECT 2069.610 18.400 2069.930 18.460 ;
        RECT 2179.090 18.400 2179.410 18.460 ;
      LAYER via ;
        RECT 2069.640 18.400 2069.900 18.660 ;
        RECT 2179.120 18.400 2179.380 18.660 ;
      LAYER met2 ;
        RECT 2069.700 18.690 2069.840 54.000 ;
        RECT 2069.640 18.370 2069.900 18.690 ;
        RECT 2179.120 18.370 2179.380 18.690 ;
        RECT 2179.180 2.400 2179.320 18.370 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2082.950 17.580 2083.270 17.640 ;
        RECT 2197.030 17.580 2197.350 17.640 ;
        RECT 2082.950 17.440 2197.350 17.580 ;
        RECT 2082.950 17.380 2083.270 17.440 ;
        RECT 2197.030 17.380 2197.350 17.440 ;
      LAYER via ;
        RECT 2082.980 17.380 2083.240 17.640 ;
        RECT 2197.060 17.380 2197.320 17.640 ;
      LAYER met2 ;
        RECT 2083.040 17.670 2083.180 54.000 ;
        RECT 2082.980 17.350 2083.240 17.670 ;
        RECT 2197.060 17.350 2197.320 17.670 ;
        RECT 2197.120 2.400 2197.260 17.350 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2104.110 20.640 2104.430 20.700 ;
        RECT 2214.970 20.640 2215.290 20.700 ;
        RECT 2104.110 20.500 2215.290 20.640 ;
        RECT 2104.110 20.440 2104.430 20.500 ;
        RECT 2214.970 20.440 2215.290 20.500 ;
      LAYER via ;
        RECT 2104.140 20.440 2104.400 20.700 ;
        RECT 2215.000 20.440 2215.260 20.700 ;
      LAYER met2 ;
        RECT 2104.200 20.730 2104.340 54.000 ;
        RECT 2104.140 20.410 2104.400 20.730 ;
        RECT 2215.000 20.410 2215.260 20.730 ;
        RECT 2215.060 2.400 2215.200 20.410 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2117.910 20.300 2118.230 20.360 ;
        RECT 2232.910 20.300 2233.230 20.360 ;
        RECT 2117.910 20.160 2233.230 20.300 ;
        RECT 2117.910 20.100 2118.230 20.160 ;
        RECT 2232.910 20.100 2233.230 20.160 ;
      LAYER via ;
        RECT 2117.940 20.100 2118.200 20.360 ;
        RECT 2232.940 20.100 2233.200 20.360 ;
      LAYER met2 ;
        RECT 2118.000 20.390 2118.140 54.000 ;
        RECT 2117.940 20.070 2118.200 20.390 ;
        RECT 2232.940 20.070 2233.200 20.390 ;
        RECT 2233.000 2.400 2233.140 20.070 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 787.590 16.560 787.910 16.620 ;
        RECT 793.110 16.560 793.430 16.620 ;
        RECT 787.590 16.420 793.430 16.560 ;
        RECT 787.590 16.360 787.910 16.420 ;
        RECT 793.110 16.360 793.430 16.420 ;
      LAYER via ;
        RECT 787.620 16.360 787.880 16.620 ;
        RECT 793.140 16.360 793.400 16.620 ;
      LAYER met2 ;
        RECT 793.200 16.650 793.340 54.000 ;
        RECT 787.620 16.330 787.880 16.650 ;
        RECT 793.140 16.330 793.400 16.650 ;
        RECT 787.680 2.400 787.820 16.330 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2132.170 17.240 2132.490 17.300 ;
        RECT 2250.850 17.240 2251.170 17.300 ;
        RECT 2132.170 17.100 2251.170 17.240 ;
        RECT 2132.170 17.040 2132.490 17.100 ;
        RECT 2250.850 17.040 2251.170 17.100 ;
      LAYER via ;
        RECT 2132.200 17.040 2132.460 17.300 ;
        RECT 2250.880 17.040 2251.140 17.300 ;
      LAYER met2 ;
        RECT 2131.800 18.090 2131.940 54.000 ;
        RECT 2131.800 17.950 2132.400 18.090 ;
        RECT 2132.260 17.330 2132.400 17.950 ;
        RECT 2132.200 17.010 2132.460 17.330 ;
        RECT 2250.880 17.010 2251.140 17.330 ;
        RECT 2250.940 2.400 2251.080 17.010 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2145.510 18.260 2145.830 18.320 ;
        RECT 2268.330 18.260 2268.650 18.320 ;
        RECT 2145.510 18.120 2268.650 18.260 ;
        RECT 2145.510 18.060 2145.830 18.120 ;
        RECT 2268.330 18.060 2268.650 18.120 ;
      LAYER via ;
        RECT 2145.540 18.060 2145.800 18.320 ;
        RECT 2268.360 18.060 2268.620 18.320 ;
      LAYER met2 ;
        RECT 2145.600 18.350 2145.740 54.000 ;
        RECT 2145.540 18.030 2145.800 18.350 ;
        RECT 2268.360 18.030 2268.620 18.350 ;
        RECT 2268.420 2.400 2268.560 18.030 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2158.850 17.920 2159.170 17.980 ;
        RECT 2286.270 17.920 2286.590 17.980 ;
        RECT 2158.850 17.780 2286.590 17.920 ;
        RECT 2158.850 17.720 2159.170 17.780 ;
        RECT 2286.270 17.720 2286.590 17.780 ;
      LAYER via ;
        RECT 2158.880 17.720 2159.140 17.980 ;
        RECT 2286.300 17.720 2286.560 17.980 ;
      LAYER met2 ;
        RECT 2158.940 18.010 2159.080 54.000 ;
        RECT 2158.880 17.690 2159.140 18.010 ;
        RECT 2286.300 17.690 2286.560 18.010 ;
        RECT 2286.360 2.400 2286.500 17.690 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.010 15.880 2180.330 15.940 ;
        RECT 2304.210 15.880 2304.530 15.940 ;
        RECT 2180.010 15.740 2304.530 15.880 ;
        RECT 2180.010 15.680 2180.330 15.740 ;
        RECT 2304.210 15.680 2304.530 15.740 ;
      LAYER via ;
        RECT 2180.040 15.680 2180.300 15.940 ;
        RECT 2304.240 15.680 2304.500 15.940 ;
      LAYER met2 ;
        RECT 2180.100 15.970 2180.240 54.000 ;
        RECT 2180.040 15.650 2180.300 15.970 ;
        RECT 2304.240 15.650 2304.500 15.970 ;
        RECT 2304.300 2.400 2304.440 15.650 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2193.810 19.960 2194.130 20.020 ;
        RECT 2322.150 19.960 2322.470 20.020 ;
        RECT 2193.810 19.820 2322.470 19.960 ;
        RECT 2193.810 19.760 2194.130 19.820 ;
        RECT 2322.150 19.760 2322.470 19.820 ;
      LAYER via ;
        RECT 2193.840 19.760 2194.100 20.020 ;
        RECT 2322.180 19.760 2322.440 20.020 ;
      LAYER met2 ;
        RECT 2193.900 20.050 2194.040 54.000 ;
        RECT 2193.840 19.730 2194.100 20.050 ;
        RECT 2322.180 19.730 2322.440 20.050 ;
        RECT 2322.240 2.400 2322.380 19.730 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2207.610 18.600 2207.930 18.660 ;
        RECT 2339.170 18.600 2339.490 18.660 ;
        RECT 2207.610 18.460 2339.490 18.600 ;
        RECT 2207.610 18.400 2207.930 18.460 ;
        RECT 2339.170 18.400 2339.490 18.460 ;
      LAYER via ;
        RECT 2207.640 18.400 2207.900 18.660 ;
        RECT 2339.200 18.400 2339.460 18.660 ;
      LAYER met2 ;
        RECT 2207.700 18.690 2207.840 54.000 ;
        RECT 2207.640 18.370 2207.900 18.690 ;
        RECT 2339.200 18.370 2339.460 18.690 ;
        RECT 2339.260 16.730 2339.400 18.370 ;
        RECT 2339.260 16.590 2339.860 16.730 ;
        RECT 2339.720 2.400 2339.860 16.590 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2220.950 19.620 2221.270 19.680 ;
        RECT 2357.570 19.620 2357.890 19.680 ;
        RECT 2220.950 19.480 2357.890 19.620 ;
        RECT 2220.950 19.420 2221.270 19.480 ;
        RECT 2357.570 19.420 2357.890 19.480 ;
      LAYER via ;
        RECT 2220.980 19.420 2221.240 19.680 ;
        RECT 2357.600 19.420 2357.860 19.680 ;
      LAYER met2 ;
        RECT 2221.040 19.710 2221.180 54.000 ;
        RECT 2220.980 19.390 2221.240 19.710 ;
        RECT 2357.600 19.390 2357.860 19.710 ;
        RECT 2357.660 2.400 2357.800 19.390 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2242.110 14.520 2242.430 14.580 ;
        RECT 2375.510 14.520 2375.830 14.580 ;
        RECT 2242.110 14.380 2375.830 14.520 ;
        RECT 2242.110 14.320 2242.430 14.380 ;
        RECT 2375.510 14.320 2375.830 14.380 ;
      LAYER via ;
        RECT 2242.140 14.320 2242.400 14.580 ;
        RECT 2375.540 14.320 2375.800 14.580 ;
      LAYER met2 ;
        RECT 2242.200 14.610 2242.340 54.000 ;
        RECT 2242.140 14.290 2242.400 14.610 ;
        RECT 2375.540 14.290 2375.800 14.610 ;
        RECT 2375.600 2.400 2375.740 14.290 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2255.910 14.860 2256.230 14.920 ;
        RECT 2393.450 14.860 2393.770 14.920 ;
        RECT 2255.910 14.720 2393.770 14.860 ;
        RECT 2255.910 14.660 2256.230 14.720 ;
        RECT 2393.450 14.660 2393.770 14.720 ;
      LAYER via ;
        RECT 2255.940 14.660 2256.200 14.920 ;
        RECT 2393.480 14.660 2393.740 14.920 ;
      LAYER met2 ;
        RECT 2256.000 14.950 2256.140 54.000 ;
        RECT 2255.940 14.630 2256.200 14.950 ;
        RECT 2393.480 14.630 2393.740 14.950 ;
        RECT 2393.540 2.400 2393.680 14.630 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 18.260 2270.030 18.320 ;
        RECT 2411.390 18.260 2411.710 18.320 ;
        RECT 2269.710 18.120 2411.710 18.260 ;
        RECT 2269.710 18.060 2270.030 18.120 ;
        RECT 2411.390 18.060 2411.710 18.120 ;
      LAYER via ;
        RECT 2269.740 18.060 2270.000 18.320 ;
        RECT 2411.420 18.060 2411.680 18.320 ;
      LAYER met2 ;
        RECT 2269.800 18.350 2269.940 54.000 ;
        RECT 2269.740 18.030 2270.000 18.350 ;
        RECT 2411.420 18.030 2411.680 18.350 ;
        RECT 2411.480 2.400 2411.620 18.030 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 807.000 17.410 807.140 54.000 ;
        RECT 805.620 17.270 807.140 17.410 ;
        RECT 805.620 2.400 805.760 17.270 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 17.240 3.150 17.300 ;
        RECT 201.090 17.240 201.410 17.300 ;
        RECT 2.830 17.100 201.410 17.240 ;
        RECT 2.830 17.040 3.150 17.100 ;
        RECT 201.090 17.040 201.410 17.100 ;
      LAYER via ;
        RECT 2.860 17.040 3.120 17.300 ;
        RECT 201.120 17.040 201.380 17.300 ;
      LAYER met2 ;
        RECT 201.180 17.330 201.320 54.000 ;
        RECT 2.860 17.010 3.120 17.330 ;
        RECT 201.120 17.010 201.380 17.330 ;
        RECT 2.920 2.400 3.060 17.010 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 200.630 17.580 200.950 17.640 ;
        RECT 8.350 17.440 200.950 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 200.630 17.380 200.950 17.440 ;
      LAYER via ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 200.660 17.380 200.920 17.640 ;
      LAYER met2 ;
        RECT 200.720 17.670 200.860 54.000 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 200.660 17.350 200.920 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 17.920 14.650 17.980 ;
        RECT 207.070 17.920 207.390 17.980 ;
        RECT 14.330 17.780 207.390 17.920 ;
        RECT 14.330 17.720 14.650 17.780 ;
        RECT 207.070 17.720 207.390 17.780 ;
      LAYER via ;
        RECT 14.360 17.720 14.620 17.980 ;
        RECT 207.100 17.720 207.360 17.980 ;
      LAYER met2 ;
        RECT 207.160 18.010 207.300 54.000 ;
        RECT 14.360 17.690 14.620 18.010 ;
        RECT 207.100 17.690 207.360 18.010 ;
        RECT 14.420 2.400 14.560 17.690 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 24.040 38.570 24.100 ;
        RECT 227.770 24.040 228.090 24.100 ;
        RECT 38.250 23.900 228.090 24.040 ;
        RECT 38.250 23.840 38.570 23.900 ;
        RECT 227.770 23.840 228.090 23.900 ;
      LAYER via ;
        RECT 38.280 23.840 38.540 24.100 ;
        RECT 227.800 23.840 228.060 24.100 ;
      LAYER met2 ;
        RECT 227.860 24.130 228.000 54.000 ;
        RECT 38.280 23.810 38.540 24.130 ;
        RECT 227.800 23.810 228.060 24.130 ;
        RECT 38.340 2.400 38.480 23.810 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 269.260 17.100 353.120 17.240 ;
        RECT 240.650 16.900 240.970 16.960 ;
        RECT 269.260 16.900 269.400 17.100 ;
        RECT 240.650 16.760 269.400 16.900 ;
        RECT 240.650 16.700 240.970 16.760 ;
        RECT 352.980 16.560 353.120 17.100 ;
        RECT 400.270 16.560 400.590 16.620 ;
        RECT 352.980 16.420 400.590 16.560 ;
        RECT 400.270 16.360 400.590 16.420 ;
      LAYER via ;
        RECT 240.680 16.700 240.940 16.960 ;
        RECT 400.300 16.360 400.560 16.620 ;
      LAYER met2 ;
        RECT 240.680 16.670 240.940 16.990 ;
        RECT 240.740 2.400 240.880 16.670 ;
        RECT 400.360 16.650 400.500 54.000 ;
        RECT 400.300 16.330 400.560 16.650 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 375.890 19.620 376.210 19.680 ;
        RECT 414.990 19.620 415.310 19.680 ;
        RECT 375.890 19.480 415.310 19.620 ;
        RECT 375.890 19.420 376.210 19.480 ;
        RECT 414.990 19.420 415.310 19.480 ;
        RECT 258.130 18.260 258.450 18.320 ;
        RECT 375.890 18.260 376.210 18.320 ;
        RECT 258.130 18.120 376.210 18.260 ;
        RECT 258.130 18.060 258.450 18.120 ;
        RECT 375.890 18.060 376.210 18.120 ;
      LAYER via ;
        RECT 375.920 19.420 376.180 19.680 ;
        RECT 415.020 19.420 415.280 19.680 ;
        RECT 258.160 18.060 258.420 18.320 ;
        RECT 375.920 18.060 376.180 18.320 ;
      LAYER met2 ;
        RECT 415.080 19.710 415.220 54.000 ;
        RECT 375.920 19.390 376.180 19.710 ;
        RECT 415.020 19.390 415.280 19.710 ;
        RECT 375.980 18.350 376.120 19.390 ;
        RECT 258.160 18.030 258.420 18.350 ;
        RECT 375.920 18.030 376.180 18.350 ;
        RECT 258.220 2.400 258.360 18.030 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 424.190 19.620 424.510 19.680 ;
        RECT 434.770 19.620 435.090 19.680 ;
        RECT 424.190 19.480 435.090 19.620 ;
        RECT 424.190 19.420 424.510 19.480 ;
        RECT 434.770 19.420 435.090 19.480 ;
        RECT 310.570 17.920 310.890 17.980 ;
        RECT 424.190 17.920 424.510 17.980 ;
        RECT 310.570 17.780 424.510 17.920 ;
        RECT 310.570 17.720 310.890 17.780 ;
        RECT 424.190 17.720 424.510 17.780 ;
        RECT 276.070 16.900 276.390 16.960 ;
        RECT 310.570 16.900 310.890 16.960 ;
        RECT 276.070 16.760 310.890 16.900 ;
        RECT 276.070 16.700 276.390 16.760 ;
        RECT 310.570 16.700 310.890 16.760 ;
      LAYER via ;
        RECT 424.220 19.420 424.480 19.680 ;
        RECT 434.800 19.420 435.060 19.680 ;
        RECT 310.600 17.720 310.860 17.980 ;
        RECT 424.220 17.720 424.480 17.980 ;
        RECT 276.100 16.700 276.360 16.960 ;
        RECT 310.600 16.700 310.860 16.960 ;
      LAYER met2 ;
        RECT 434.860 19.710 435.000 54.000 ;
        RECT 424.220 19.390 424.480 19.710 ;
        RECT 434.800 19.390 435.060 19.710 ;
        RECT 424.280 18.010 424.420 19.390 ;
        RECT 310.600 17.690 310.860 18.010 ;
        RECT 424.220 17.690 424.480 18.010 ;
        RECT 310.660 16.990 310.800 17.690 ;
        RECT 276.100 16.670 276.360 16.990 ;
        RECT 310.600 16.670 310.860 16.990 ;
        RECT 276.160 2.400 276.300 16.670 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 18.600 294.330 18.660 ;
        RECT 449.030 18.600 449.350 18.660 ;
        RECT 294.010 18.460 449.350 18.600 ;
        RECT 294.010 18.400 294.330 18.460 ;
        RECT 449.030 18.400 449.350 18.460 ;
      LAYER via ;
        RECT 294.040 18.400 294.300 18.660 ;
        RECT 449.060 18.400 449.320 18.660 ;
      LAYER met2 ;
        RECT 449.120 18.690 449.260 54.000 ;
        RECT 294.040 18.370 294.300 18.690 ;
        RECT 449.060 18.370 449.320 18.690 ;
        RECT 294.100 2.400 294.240 18.370 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 18.940 312.270 19.000 ;
        RECT 462.370 18.940 462.690 19.000 ;
        RECT 311.950 18.800 462.690 18.940 ;
        RECT 311.950 18.740 312.270 18.800 ;
        RECT 462.370 18.740 462.690 18.800 ;
      LAYER via ;
        RECT 311.980 18.740 312.240 19.000 ;
        RECT 462.400 18.740 462.660 19.000 ;
      LAYER met2 ;
        RECT 462.460 19.030 462.600 54.000 ;
        RECT 311.980 18.710 312.240 19.030 ;
        RECT 462.400 18.710 462.660 19.030 ;
        RECT 312.040 2.400 312.180 18.710 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 24.380 330.210 24.440 ;
        RECT 476.170 24.380 476.490 24.440 ;
        RECT 329.890 24.240 476.490 24.380 ;
        RECT 329.890 24.180 330.210 24.240 ;
        RECT 476.170 24.180 476.490 24.240 ;
      LAYER via ;
        RECT 329.920 24.180 330.180 24.440 ;
        RECT 476.200 24.180 476.460 24.440 ;
      LAYER met2 ;
        RECT 476.260 24.470 476.400 54.000 ;
        RECT 329.920 24.150 330.180 24.470 ;
        RECT 476.200 24.150 476.460 24.470 ;
        RECT 329.980 2.400 330.120 24.150 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 24.720 347.690 24.780 ;
        RECT 491.350 24.720 491.670 24.780 ;
        RECT 347.370 24.580 491.670 24.720 ;
        RECT 347.370 24.520 347.690 24.580 ;
        RECT 491.350 24.520 491.670 24.580 ;
      LAYER via ;
        RECT 347.400 24.520 347.660 24.780 ;
        RECT 491.380 24.520 491.640 24.780 ;
      LAYER met2 ;
        RECT 491.440 24.810 491.580 54.000 ;
        RECT 347.400 24.490 347.660 24.810 ;
        RECT 491.380 24.490 491.640 24.810 ;
        RECT 347.460 2.400 347.600 24.490 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 364.850 19.280 365.170 19.340 ;
        RECT 510.670 19.280 510.990 19.340 ;
        RECT 364.850 19.140 510.990 19.280 ;
        RECT 364.850 19.080 365.170 19.140 ;
        RECT 510.670 19.080 510.990 19.140 ;
      LAYER via ;
        RECT 364.880 19.080 365.140 19.340 ;
        RECT 510.700 19.080 510.960 19.340 ;
      LAYER met2 ;
        RECT 510.760 19.370 510.900 54.000 ;
        RECT 364.880 19.050 365.140 19.370 ;
        RECT 510.700 19.050 510.960 19.370 ;
        RECT 364.940 9.930 365.080 19.050 ;
        RECT 364.940 9.790 365.540 9.930 ;
        RECT 365.400 2.400 365.540 9.790 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 400.360 17.440 519.640 17.580 ;
        RECT 383.250 17.240 383.570 17.300 ;
        RECT 400.360 17.240 400.500 17.440 ;
        RECT 383.250 17.100 400.500 17.240 ;
        RECT 519.500 17.240 519.640 17.440 ;
        RECT 524.470 17.240 524.790 17.300 ;
        RECT 519.500 17.100 524.790 17.240 ;
        RECT 383.250 17.040 383.570 17.100 ;
        RECT 524.470 17.040 524.790 17.100 ;
      LAYER via ;
        RECT 383.280 17.040 383.540 17.300 ;
        RECT 524.500 17.040 524.760 17.300 ;
      LAYER met2 ;
        RECT 524.560 17.330 524.700 54.000 ;
        RECT 383.280 17.010 383.540 17.330 ;
        RECT 524.500 17.010 524.760 17.330 ;
        RECT 383.340 2.400 383.480 17.010 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 17.240 401.510 17.300 ;
        RECT 538.270 17.240 538.590 17.300 ;
        RECT 401.190 17.100 519.180 17.240 ;
        RECT 401.190 17.040 401.510 17.100 ;
        RECT 519.040 16.900 519.180 17.100 ;
        RECT 525.020 17.100 538.590 17.240 ;
        RECT 525.020 16.900 525.160 17.100 ;
        RECT 538.270 17.040 538.590 17.100 ;
        RECT 519.040 16.760 525.160 16.900 ;
      LAYER via ;
        RECT 401.220 17.040 401.480 17.300 ;
        RECT 538.300 17.040 538.560 17.300 ;
      LAYER met2 ;
        RECT 538.360 17.330 538.500 54.000 ;
        RECT 401.220 17.010 401.480 17.330 ;
        RECT 538.300 17.010 538.560 17.330 ;
        RECT 401.280 2.400 401.420 17.010 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 62.170 24.720 62.490 24.780 ;
        RECT 248.470 24.720 248.790 24.780 ;
        RECT 62.170 24.580 248.790 24.720 ;
        RECT 62.170 24.520 62.490 24.580 ;
        RECT 248.470 24.520 248.790 24.580 ;
      LAYER via ;
        RECT 62.200 24.520 62.460 24.780 ;
        RECT 248.500 24.520 248.760 24.780 ;
      LAYER met2 ;
        RECT 248.560 24.810 248.700 54.000 ;
        RECT 62.200 24.490 62.460 24.810 ;
        RECT 248.500 24.490 248.760 24.810 ;
        RECT 62.260 2.400 62.400 24.490 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 20.300 419.450 20.360 ;
        RECT 552.530 20.300 552.850 20.360 ;
        RECT 419.130 20.160 552.850 20.300 ;
        RECT 419.130 20.100 419.450 20.160 ;
        RECT 552.530 20.100 552.850 20.160 ;
      LAYER via ;
        RECT 419.160 20.100 419.420 20.360 ;
        RECT 552.560 20.100 552.820 20.360 ;
      LAYER met2 ;
        RECT 552.620 20.390 552.760 54.000 ;
        RECT 419.160 20.070 419.420 20.390 ;
        RECT 552.560 20.070 552.820 20.390 ;
        RECT 419.220 2.400 419.360 20.070 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 19.620 436.930 19.680 ;
        RECT 566.790 19.620 567.110 19.680 ;
        RECT 436.610 19.480 567.110 19.620 ;
        RECT 436.610 19.420 436.930 19.480 ;
        RECT 566.790 19.420 567.110 19.480 ;
      LAYER via ;
        RECT 436.640 19.420 436.900 19.680 ;
        RECT 566.820 19.420 567.080 19.680 ;
      LAYER met2 ;
        RECT 566.880 19.710 567.020 54.000 ;
        RECT 436.640 19.390 436.900 19.710 ;
        RECT 566.820 19.390 567.080 19.710 ;
        RECT 436.700 2.400 436.840 19.390 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 454.550 18.600 454.870 18.660 ;
        RECT 454.550 18.460 455.700 18.600 ;
        RECT 454.550 18.400 454.870 18.460 ;
        RECT 455.560 17.920 455.700 18.460 ;
        RECT 587.030 17.920 587.350 17.980 ;
        RECT 455.560 17.780 587.350 17.920 ;
        RECT 587.030 17.720 587.350 17.780 ;
      LAYER via ;
        RECT 454.580 18.400 454.840 18.660 ;
        RECT 587.060 17.720 587.320 17.980 ;
      LAYER met2 ;
        RECT 454.580 18.370 454.840 18.690 ;
        RECT 454.640 2.400 454.780 18.370 ;
        RECT 587.120 18.010 587.260 54.000 ;
        RECT 587.060 17.690 587.320 18.010 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.490 18.600 472.810 18.660 ;
        RECT 600.370 18.600 600.690 18.660 ;
        RECT 472.490 18.460 600.690 18.600 ;
        RECT 472.490 18.400 472.810 18.460 ;
        RECT 600.370 18.400 600.690 18.460 ;
      LAYER via ;
        RECT 472.520 18.400 472.780 18.660 ;
        RECT 600.400 18.400 600.660 18.660 ;
      LAYER met2 ;
        RECT 600.460 18.690 600.600 54.000 ;
        RECT 472.520 18.370 472.780 18.690 ;
        RECT 600.400 18.370 600.660 18.690 ;
        RECT 472.580 2.400 472.720 18.370 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 490.430 19.960 490.750 20.020 ;
        RECT 614.170 19.960 614.490 20.020 ;
        RECT 490.430 19.820 614.490 19.960 ;
        RECT 490.430 19.760 490.750 19.820 ;
        RECT 614.170 19.760 614.490 19.820 ;
      LAYER via ;
        RECT 490.460 19.760 490.720 20.020 ;
        RECT 614.200 19.760 614.460 20.020 ;
      LAYER met2 ;
        RECT 614.260 20.050 614.400 54.000 ;
        RECT 490.460 19.730 490.720 20.050 ;
        RECT 614.200 19.730 614.460 20.050 ;
        RECT 490.520 2.400 490.660 19.730 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 18.940 508.230 19.000 ;
        RECT 628.890 18.940 629.210 19.000 ;
        RECT 507.910 18.800 629.210 18.940 ;
        RECT 507.910 18.740 508.230 18.800 ;
        RECT 628.890 18.740 629.210 18.800 ;
      LAYER via ;
        RECT 507.940 18.740 508.200 19.000 ;
        RECT 628.920 18.740 629.180 19.000 ;
      LAYER met2 ;
        RECT 628.980 19.030 629.120 54.000 ;
        RECT 507.940 18.710 508.200 19.030 ;
        RECT 628.920 18.710 629.180 19.030 ;
        RECT 508.000 2.400 508.140 18.710 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.670 18.600 648.990 18.660 ;
        RECT 614.720 18.460 648.990 18.600 ;
        RECT 614.720 17.580 614.860 18.460 ;
        RECT 648.670 18.400 648.990 18.460 ;
        RECT 579.760 17.440 614.860 17.580 ;
        RECT 525.850 16.900 526.170 16.960 ;
        RECT 579.760 16.900 579.900 17.440 ;
        RECT 525.850 16.760 579.900 16.900 ;
        RECT 525.850 16.700 526.170 16.760 ;
      LAYER via ;
        RECT 648.700 18.400 648.960 18.660 ;
        RECT 525.880 16.700 526.140 16.960 ;
      LAYER met2 ;
        RECT 648.760 18.690 648.900 54.000 ;
        RECT 648.700 18.370 648.960 18.690 ;
        RECT 525.880 16.670 526.140 16.990 ;
        RECT 525.940 2.400 526.080 16.670 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 580.220 17.100 662.700 17.240 ;
        RECT 543.790 16.560 544.110 16.620 ;
        RECT 580.220 16.560 580.360 17.100 ;
        RECT 543.790 16.420 580.360 16.560 ;
        RECT 662.560 16.560 662.700 17.100 ;
        RECT 663.390 16.560 663.710 16.620 ;
        RECT 662.560 16.420 663.710 16.560 ;
        RECT 543.790 16.360 544.110 16.420 ;
        RECT 663.390 16.360 663.710 16.420 ;
      LAYER via ;
        RECT 543.820 16.360 544.080 16.620 ;
        RECT 663.420 16.360 663.680 16.620 ;
      LAYER met2 ;
        RECT 663.480 16.650 663.620 54.000 ;
        RECT 543.820 16.330 544.080 16.650 ;
        RECT 663.420 16.330 663.680 16.650 ;
        RECT 543.880 2.400 544.020 16.330 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 20.640 562.050 20.700 ;
        RECT 565.410 20.640 565.730 20.700 ;
        RECT 561.730 20.500 565.730 20.640 ;
        RECT 561.730 20.440 562.050 20.500 ;
        RECT 565.410 20.440 565.730 20.500 ;
      LAYER via ;
        RECT 561.760 20.440 562.020 20.700 ;
        RECT 565.440 20.440 565.700 20.700 ;
      LAYER met2 ;
        RECT 565.500 20.730 565.640 54.000 ;
        RECT 561.760 20.410 562.020 20.730 ;
        RECT 565.440 20.410 565.700 20.730 ;
        RECT 561.820 2.400 561.960 20.410 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.670 20.640 579.990 20.700 ;
        RECT 585.650 20.640 585.970 20.700 ;
        RECT 579.670 20.500 585.970 20.640 ;
        RECT 579.670 20.440 579.990 20.500 ;
        RECT 585.650 20.440 585.970 20.500 ;
      LAYER via ;
        RECT 579.700 20.440 579.960 20.700 ;
        RECT 585.680 20.440 585.940 20.700 ;
      LAYER met2 ;
        RECT 585.740 20.730 585.880 54.000 ;
        RECT 579.700 20.410 579.960 20.730 ;
        RECT 585.680 20.410 585.940 20.730 ;
        RECT 579.760 2.400 579.900 20.410 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 24.380 86.410 24.440 ;
        RECT 269.170 24.380 269.490 24.440 ;
        RECT 86.090 24.240 269.490 24.380 ;
        RECT 86.090 24.180 86.410 24.240 ;
        RECT 269.170 24.180 269.490 24.240 ;
      LAYER via ;
        RECT 86.120 24.180 86.380 24.440 ;
        RECT 269.200 24.180 269.460 24.440 ;
      LAYER met2 ;
        RECT 269.260 24.470 269.400 54.000 ;
        RECT 86.120 24.150 86.380 24.470 ;
        RECT 269.200 24.150 269.460 24.470 ;
        RECT 86.180 2.400 86.320 24.150 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 597.150 17.920 597.470 17.980 ;
        RECT 599.910 17.920 600.230 17.980 ;
        RECT 597.150 17.780 600.230 17.920 ;
        RECT 597.150 17.720 597.470 17.780 ;
        RECT 599.910 17.720 600.230 17.780 ;
      LAYER via ;
        RECT 597.180 17.720 597.440 17.980 ;
        RECT 599.940 17.720 600.200 17.980 ;
      LAYER met2 ;
        RECT 600.000 18.010 600.140 54.000 ;
        RECT 597.180 17.690 597.440 18.010 ;
        RECT 599.940 17.690 600.200 18.010 ;
        RECT 597.240 2.400 597.380 17.690 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 615.090 17.580 615.410 17.640 ;
        RECT 620.610 17.580 620.930 17.640 ;
        RECT 615.090 17.440 620.930 17.580 ;
        RECT 615.090 17.380 615.410 17.440 ;
        RECT 620.610 17.380 620.930 17.440 ;
      LAYER via ;
        RECT 615.120 17.380 615.380 17.640 ;
        RECT 620.640 17.380 620.900 17.640 ;
      LAYER met2 ;
        RECT 620.700 17.670 620.840 54.000 ;
        RECT 615.120 17.350 615.380 17.670 ;
        RECT 620.640 17.350 620.900 17.670 ;
        RECT 615.180 2.400 615.320 17.350 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 25.060 109.870 25.120 ;
        RECT 289.870 25.060 290.190 25.120 ;
        RECT 109.550 24.920 290.190 25.060 ;
        RECT 109.550 24.860 109.870 24.920 ;
        RECT 289.870 24.860 290.190 24.920 ;
      LAYER via ;
        RECT 109.580 24.860 109.840 25.120 ;
        RECT 289.900 24.860 290.160 25.120 ;
      LAYER met2 ;
        RECT 289.960 25.150 290.100 54.000 ;
        RECT 109.580 24.830 109.840 25.150 ;
        RECT 289.900 24.830 290.160 25.150 ;
        RECT 109.640 2.400 109.780 24.830 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 133.470 25.400 133.790 25.460 ;
        RECT 310.570 25.400 310.890 25.460 ;
        RECT 133.470 25.260 310.890 25.400 ;
        RECT 133.470 25.200 133.790 25.260 ;
        RECT 310.570 25.200 310.890 25.260 ;
      LAYER via ;
        RECT 133.500 25.200 133.760 25.460 ;
        RECT 310.600 25.200 310.860 25.460 ;
      LAYER met2 ;
        RECT 310.660 25.490 310.800 54.000 ;
        RECT 133.500 25.170 133.760 25.490 ;
        RECT 310.600 25.170 310.860 25.490 ;
        RECT 133.560 2.400 133.700 25.170 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 25.740 151.730 25.800 ;
        RECT 324.370 25.740 324.690 25.800 ;
        RECT 151.410 25.600 324.690 25.740 ;
        RECT 151.410 25.540 151.730 25.600 ;
        RECT 324.370 25.540 324.690 25.600 ;
      LAYER via ;
        RECT 151.440 25.540 151.700 25.800 ;
        RECT 324.400 25.540 324.660 25.800 ;
      LAYER met2 ;
        RECT 324.460 25.830 324.600 54.000 ;
        RECT 151.440 25.510 151.700 25.830 ;
        RECT 324.400 25.510 324.660 25.830 ;
        RECT 151.500 2.400 151.640 25.510 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 169.350 26.420 169.670 26.480 ;
        RECT 338.170 26.420 338.490 26.480 ;
        RECT 169.350 26.280 338.490 26.420 ;
        RECT 169.350 26.220 169.670 26.280 ;
        RECT 338.170 26.220 338.490 26.280 ;
      LAYER via ;
        RECT 169.380 26.220 169.640 26.480 ;
        RECT 338.200 26.220 338.460 26.480 ;
      LAYER met2 ;
        RECT 338.260 26.510 338.400 54.000 ;
        RECT 169.380 26.190 169.640 26.510 ;
        RECT 338.200 26.190 338.460 26.510 ;
        RECT 169.440 2.400 169.580 26.190 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 26.760 187.150 26.820 ;
        RECT 353.350 26.760 353.670 26.820 ;
        RECT 186.830 26.620 353.670 26.760 ;
        RECT 186.830 26.560 187.150 26.620 ;
        RECT 353.350 26.560 353.670 26.620 ;
      LAYER via ;
        RECT 186.860 26.560 187.120 26.820 ;
        RECT 353.380 26.560 353.640 26.820 ;
      LAYER met2 ;
        RECT 353.440 26.850 353.580 54.000 ;
        RECT 186.860 26.530 187.120 26.850 ;
        RECT 353.380 26.530 353.640 26.850 ;
        RECT 186.920 2.400 187.060 26.530 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 204.770 26.080 205.090 26.140 ;
        RECT 373.130 26.080 373.450 26.140 ;
        RECT 204.770 25.940 373.450 26.080 ;
        RECT 204.770 25.880 205.090 25.940 ;
        RECT 373.130 25.880 373.450 25.940 ;
      LAYER via ;
        RECT 204.800 25.880 205.060 26.140 ;
        RECT 373.160 25.880 373.420 26.140 ;
      LAYER met2 ;
        RECT 373.220 26.170 373.360 54.000 ;
        RECT 204.800 25.850 205.060 26.170 ;
        RECT 373.160 25.850 373.420 26.170 ;
        RECT 204.860 2.400 205.000 25.850 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 236.970 24.040 237.290 24.100 ;
        RECT 386.470 24.040 386.790 24.100 ;
        RECT 236.970 23.900 386.790 24.040 ;
        RECT 236.970 23.840 237.290 23.900 ;
        RECT 386.470 23.840 386.790 23.900 ;
        RECT 222.710 18.600 223.030 18.660 ;
        RECT 236.970 18.600 237.290 18.660 ;
        RECT 222.710 18.460 237.290 18.600 ;
        RECT 222.710 18.400 223.030 18.460 ;
        RECT 236.970 18.400 237.290 18.460 ;
      LAYER via ;
        RECT 237.000 23.840 237.260 24.100 ;
        RECT 386.500 23.840 386.760 24.100 ;
        RECT 222.740 18.400 223.000 18.660 ;
        RECT 237.000 18.400 237.260 18.660 ;
      LAYER met2 ;
        RECT 386.560 24.130 386.700 54.000 ;
        RECT 237.000 23.810 237.260 24.130 ;
        RECT 386.500 23.810 386.760 24.130 ;
        RECT 237.060 18.690 237.200 23.810 ;
        RECT 222.740 18.370 223.000 18.690 ;
        RECT 237.000 18.370 237.260 18.690 ;
        RECT 222.800 2.400 222.940 18.370 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 306.920 20.630 306.980 ;
        RECT 20.310 306.780 54.000 306.920 ;
        RECT 20.310 306.720 20.630 306.780 ;
      LAYER via ;
        RECT 20.340 306.720 20.600 306.980 ;
      LAYER met2 ;
        RECT 20.340 306.690 20.600 307.010 ;
        RECT 20.400 2.400 20.540 306.690 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.910 307.940 48.230 308.000 ;
        RECT 47.910 307.800 54.000 307.940 ;
        RECT 47.910 307.740 48.230 307.800 ;
        RECT 44.230 16.900 44.550 16.960 ;
        RECT 47.910 16.900 48.230 16.960 ;
        RECT 44.230 16.760 48.230 16.900 ;
        RECT 44.230 16.700 44.550 16.760 ;
        RECT 47.910 16.700 48.230 16.760 ;
      LAYER via ;
        RECT 47.940 307.740 48.200 308.000 ;
        RECT 44.260 16.700 44.520 16.960 ;
        RECT 47.940 16.700 48.200 16.960 ;
      LAYER met2 ;
        RECT 47.940 307.710 48.200 308.030 ;
        RECT 48.000 16.990 48.140 307.710 ;
        RECT 44.260 16.670 44.520 16.990 ;
        RECT 47.940 16.670 48.200 16.990 ;
        RECT 44.320 2.400 44.460 16.670 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 248.100 3.130 248.240 54.000 ;
        RECT 246.720 2.990 248.240 3.130 ;
        RECT 246.720 2.400 246.860 2.990 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 264.110 17.240 264.430 17.300 ;
        RECT 268.710 17.240 269.030 17.300 ;
        RECT 264.110 17.100 269.030 17.240 ;
        RECT 264.110 17.040 264.430 17.100 ;
        RECT 268.710 17.040 269.030 17.100 ;
      LAYER via ;
        RECT 264.140 17.040 264.400 17.300 ;
        RECT 268.740 17.040 269.000 17.300 ;
      LAYER met2 ;
        RECT 268.800 17.330 268.940 54.000 ;
        RECT 264.140 17.010 264.400 17.330 ;
        RECT 268.740 17.010 269.000 17.330 ;
        RECT 264.200 2.400 264.340 17.010 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.600 17.410 282.740 54.000 ;
        RECT 282.140 17.270 282.740 17.410 ;
        RECT 282.140 2.400 282.280 17.270 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 299.990 17.920 300.310 17.980 ;
        RECT 303.210 17.920 303.530 17.980 ;
        RECT 299.990 17.780 303.530 17.920 ;
        RECT 299.990 17.720 300.310 17.780 ;
        RECT 303.210 17.720 303.530 17.780 ;
      LAYER via ;
        RECT 300.020 17.720 300.280 17.980 ;
        RECT 303.240 17.720 303.500 17.980 ;
      LAYER met2 ;
        RECT 303.300 18.010 303.440 54.000 ;
        RECT 300.020 17.690 300.280 18.010 ;
        RECT 303.240 17.690 303.500 18.010 ;
        RECT 300.080 2.400 300.220 17.690 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.930 16.900 318.250 16.960 ;
        RECT 323.910 16.900 324.230 16.960 ;
        RECT 317.930 16.760 324.230 16.900 ;
        RECT 317.930 16.700 318.250 16.760 ;
        RECT 323.910 16.700 324.230 16.760 ;
      LAYER via ;
        RECT 317.960 16.700 318.220 16.960 ;
        RECT 323.940 16.700 324.200 16.960 ;
      LAYER met2 ;
        RECT 324.000 16.990 324.140 54.000 ;
        RECT 317.960 16.670 318.220 16.990 ;
        RECT 323.940 16.670 324.200 16.990 ;
        RECT 318.020 2.400 318.160 16.670 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 337.800 16.900 337.940 54.000 ;
        RECT 335.960 16.760 337.940 16.900 ;
        RECT 335.960 2.400 336.100 16.760 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 353.350 17.240 353.670 17.300 ;
        RECT 358.410 17.240 358.730 17.300 ;
        RECT 353.350 17.100 358.730 17.240 ;
        RECT 353.350 17.040 353.670 17.100 ;
        RECT 358.410 17.040 358.730 17.100 ;
      LAYER via ;
        RECT 353.380 17.040 353.640 17.300 ;
        RECT 358.440 17.040 358.700 17.300 ;
      LAYER met2 ;
        RECT 358.500 17.330 358.640 54.000 ;
        RECT 353.380 17.010 353.640 17.330 ;
        RECT 358.440 17.010 358.700 17.330 ;
        RECT 353.440 2.400 353.580 17.010 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 370.370 48.520 370.690 48.580 ;
        RECT 371.290 48.520 371.610 48.580 ;
        RECT 370.370 48.380 371.610 48.520 ;
        RECT 370.370 48.320 370.690 48.380 ;
        RECT 371.290 48.320 371.610 48.380 ;
      LAYER via ;
        RECT 370.400 48.320 370.660 48.580 ;
        RECT 371.320 48.320 371.580 48.580 ;
      LAYER met2 ;
        RECT 370.460 48.610 370.600 54.000 ;
        RECT 370.400 48.290 370.660 48.610 ;
        RECT 371.320 48.290 371.580 48.610 ;
        RECT 371.380 2.400 371.520 48.290 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 389.230 20.640 389.550 20.700 ;
        RECT 392.910 20.640 393.230 20.700 ;
        RECT 389.230 20.500 393.230 20.640 ;
        RECT 389.230 20.440 389.550 20.500 ;
        RECT 392.910 20.440 393.230 20.500 ;
      LAYER via ;
        RECT 389.260 20.440 389.520 20.700 ;
        RECT 392.940 20.440 393.200 20.700 ;
      LAYER met2 ;
        RECT 393.000 20.730 393.140 54.000 ;
        RECT 389.260 20.410 389.520 20.730 ;
        RECT 392.940 20.410 393.200 20.730 ;
        RECT 389.320 2.400 389.460 20.410 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 407.170 18.260 407.490 18.320 ;
        RECT 413.150 18.260 413.470 18.320 ;
        RECT 407.170 18.120 413.470 18.260 ;
        RECT 407.170 18.060 407.490 18.120 ;
        RECT 413.150 18.060 413.470 18.120 ;
      LAYER via ;
        RECT 407.200 18.060 407.460 18.320 ;
        RECT 413.180 18.060 413.440 18.320 ;
      LAYER met2 ;
        RECT 413.240 18.350 413.380 54.000 ;
        RECT 407.200 18.030 407.460 18.350 ;
        RECT 413.180 18.030 413.440 18.350 ;
        RECT 407.260 2.400 407.400 18.030 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.240 2.400 68.380 54.000 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 424.650 17.920 424.970 17.980 ;
        RECT 427.410 17.920 427.730 17.980 ;
        RECT 424.650 17.780 427.730 17.920 ;
        RECT 424.650 17.720 424.970 17.780 ;
        RECT 427.410 17.720 427.730 17.780 ;
      LAYER via ;
        RECT 424.680 17.720 424.940 17.980 ;
        RECT 427.440 17.720 427.700 17.980 ;
      LAYER met2 ;
        RECT 427.500 18.010 427.640 54.000 ;
        RECT 424.680 17.690 424.940 18.010 ;
        RECT 427.440 17.690 427.700 18.010 ;
        RECT 424.740 2.400 424.880 17.690 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 442.590 17.920 442.910 17.980 ;
        RECT 448.110 17.920 448.430 17.980 ;
        RECT 442.590 17.780 448.430 17.920 ;
        RECT 442.590 17.720 442.910 17.780 ;
        RECT 448.110 17.720 448.430 17.780 ;
      LAYER via ;
        RECT 442.620 17.720 442.880 17.980 ;
        RECT 448.140 17.720 448.400 17.980 ;
      LAYER met2 ;
        RECT 448.200 18.010 448.340 54.000 ;
        RECT 442.620 17.690 442.880 18.010 ;
        RECT 448.140 17.690 448.400 18.010 ;
        RECT 442.680 2.400 442.820 17.690 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 462.000 16.730 462.140 54.000 ;
        RECT 460.620 16.590 462.140 16.730 ;
        RECT 460.620 2.400 460.760 16.590 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 478.470 16.900 478.790 16.960 ;
        RECT 482.610 16.900 482.930 16.960 ;
        RECT 478.470 16.760 482.930 16.900 ;
        RECT 478.470 16.700 478.790 16.760 ;
        RECT 482.610 16.700 482.930 16.760 ;
      LAYER via ;
        RECT 478.500 16.700 478.760 16.960 ;
        RECT 482.640 16.700 482.900 16.960 ;
      LAYER met2 ;
        RECT 482.700 16.990 482.840 54.000 ;
        RECT 478.500 16.670 478.760 16.990 ;
        RECT 482.640 16.670 482.900 16.990 ;
        RECT 478.560 2.400 478.700 16.670 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.500 2.400 496.640 54.000 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 513.890 16.900 514.210 16.960 ;
        RECT 517.110 16.900 517.430 16.960 ;
        RECT 513.890 16.760 517.430 16.900 ;
        RECT 513.890 16.700 514.210 16.760 ;
        RECT 517.110 16.700 517.430 16.760 ;
      LAYER via ;
        RECT 513.920 16.700 514.180 16.960 ;
        RECT 517.140 16.700 517.400 16.960 ;
      LAYER met2 ;
        RECT 517.200 16.990 517.340 54.000 ;
        RECT 513.920 16.670 514.180 16.990 ;
        RECT 517.140 16.670 517.400 16.990 ;
        RECT 513.980 2.400 514.120 16.670 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 531.830 18.260 532.150 18.320 ;
        RECT 537.810 18.260 538.130 18.320 ;
        RECT 531.830 18.120 538.130 18.260 ;
        RECT 531.830 18.060 532.150 18.120 ;
        RECT 537.810 18.060 538.130 18.120 ;
      LAYER via ;
        RECT 531.860 18.060 532.120 18.320 ;
        RECT 537.840 18.060 538.100 18.320 ;
      LAYER met2 ;
        RECT 537.900 18.350 538.040 54.000 ;
        RECT 531.860 18.030 532.120 18.350 ;
        RECT 537.840 18.030 538.100 18.350 ;
        RECT 531.920 2.400 532.060 18.030 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 549.770 2.960 550.090 3.020 ;
        RECT 551.610 2.960 551.930 3.020 ;
        RECT 549.770 2.820 551.930 2.960 ;
        RECT 549.770 2.760 550.090 2.820 ;
        RECT 551.610 2.760 551.930 2.820 ;
      LAYER via ;
        RECT 549.800 2.760 550.060 3.020 ;
        RECT 551.640 2.760 551.900 3.020 ;
      LAYER met2 ;
        RECT 551.700 3.050 551.840 54.000 ;
        RECT 549.800 2.730 550.060 3.050 ;
        RECT 551.640 2.730 551.900 3.050 ;
        RECT 549.860 2.400 550.000 2.730 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 567.710 20.640 568.030 20.700 ;
        RECT 572.310 20.640 572.630 20.700 ;
        RECT 567.710 20.500 572.630 20.640 ;
        RECT 567.710 20.440 568.030 20.500 ;
        RECT 572.310 20.440 572.630 20.500 ;
      LAYER via ;
        RECT 567.740 20.440 568.000 20.700 ;
        RECT 572.340 20.440 572.600 20.700 ;
      LAYER met2 ;
        RECT 572.400 20.730 572.540 54.000 ;
        RECT 567.740 20.410 568.000 20.730 ;
        RECT 572.340 20.410 572.600 20.730 ;
        RECT 567.800 2.400 567.940 20.410 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 586.200 20.130 586.340 54.000 ;
        RECT 585.740 19.990 586.340 20.130 ;
        RECT 585.740 2.400 585.880 19.990 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 91.610 15.200 91.930 15.260 ;
        RECT 96.210 15.200 96.530 15.260 ;
        RECT 91.610 15.060 96.530 15.200 ;
        RECT 91.610 15.000 91.930 15.060 ;
        RECT 96.210 15.000 96.530 15.060 ;
      LAYER via ;
        RECT 91.640 15.000 91.900 15.260 ;
        RECT 96.240 15.000 96.500 15.260 ;
      LAYER met2 ;
        RECT 96.300 15.290 96.440 54.000 ;
        RECT 91.640 14.970 91.900 15.290 ;
        RECT 96.240 14.970 96.500 15.290 ;
        RECT 91.700 2.400 91.840 14.970 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 603.130 17.920 603.450 17.980 ;
        RECT 606.810 17.920 607.130 17.980 ;
        RECT 603.130 17.780 607.130 17.920 ;
        RECT 603.130 17.720 603.450 17.780 ;
        RECT 606.810 17.720 607.130 17.780 ;
      LAYER via ;
        RECT 603.160 17.720 603.420 17.980 ;
        RECT 606.840 17.720 607.100 17.980 ;
      LAYER met2 ;
        RECT 606.900 18.010 607.040 54.000 ;
        RECT 603.160 17.690 603.420 18.010 ;
        RECT 606.840 17.690 607.100 18.010 ;
        RECT 603.220 2.400 603.360 17.690 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 621.070 16.560 621.390 16.620 ;
        RECT 627.510 16.560 627.830 16.620 ;
        RECT 621.070 16.420 627.830 16.560 ;
        RECT 621.070 16.360 621.390 16.420 ;
        RECT 627.510 16.360 627.830 16.420 ;
      LAYER via ;
        RECT 621.100 16.360 621.360 16.620 ;
        RECT 627.540 16.360 627.800 16.620 ;
      LAYER met2 ;
        RECT 627.600 16.650 627.740 54.000 ;
        RECT 621.100 16.330 621.360 16.650 ;
        RECT 627.540 16.330 627.800 16.650 ;
        RECT 621.160 2.400 621.300 16.330 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.000 17.410 117.140 54.000 ;
        RECT 115.620 17.270 117.140 17.410 ;
        RECT 115.620 2.400 115.760 17.270 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 139.450 16.900 139.770 16.960 ;
        RECT 144.510 16.900 144.830 16.960 ;
        RECT 139.450 16.760 144.830 16.900 ;
        RECT 139.450 16.700 139.770 16.760 ;
        RECT 144.510 16.700 144.830 16.760 ;
      LAYER via ;
        RECT 139.480 16.700 139.740 16.960 ;
        RECT 144.540 16.700 144.800 16.960 ;
      LAYER met2 ;
        RECT 144.600 16.990 144.740 54.000 ;
        RECT 139.480 16.670 139.740 16.990 ;
        RECT 144.540 16.670 144.800 16.990 ;
        RECT 139.540 2.400 139.680 16.670 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 158.400 17.410 158.540 54.000 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 174.870 16.900 175.190 16.960 ;
        RECT 179.010 16.900 179.330 16.960 ;
        RECT 174.870 16.760 179.330 16.900 ;
        RECT 174.870 16.700 175.190 16.760 ;
        RECT 179.010 16.700 179.330 16.760 ;
      LAYER via ;
        RECT 174.900 16.700 175.160 16.960 ;
        RECT 179.040 16.700 179.300 16.960 ;
      LAYER met2 ;
        RECT 179.100 16.990 179.240 54.000 ;
        RECT 174.900 16.670 175.160 16.990 ;
        RECT 179.040 16.670 179.300 16.990 ;
        RECT 174.960 2.400 175.100 16.670 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.440 3.130 192.580 54.000 ;
        RECT 192.440 2.990 193.040 3.130 ;
        RECT 192.900 2.400 193.040 2.990 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 210.750 20.640 211.070 20.700 ;
        RECT 213.510 20.640 213.830 20.700 ;
        RECT 210.750 20.500 213.830 20.640 ;
        RECT 210.750 20.440 211.070 20.500 ;
        RECT 213.510 20.440 213.830 20.500 ;
      LAYER via ;
        RECT 210.780 20.440 211.040 20.700 ;
        RECT 213.540 20.440 213.800 20.700 ;
      LAYER met2 ;
        RECT 213.600 20.730 213.740 54.000 ;
        RECT 210.780 20.410 211.040 20.730 ;
        RECT 213.540 20.410 213.800 20.730 ;
        RECT 210.840 2.400 210.980 20.410 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 228.690 17.580 229.010 17.640 ;
        RECT 234.210 17.580 234.530 17.640 ;
        RECT 228.690 17.440 234.530 17.580 ;
        RECT 228.690 17.380 229.010 17.440 ;
        RECT 234.210 17.380 234.530 17.440 ;
      LAYER via ;
        RECT 228.720 17.380 228.980 17.640 ;
        RECT 234.240 17.380 234.500 17.640 ;
      LAYER met2 ;
        RECT 234.300 17.670 234.440 54.000 ;
        RECT 228.720 17.350 228.980 17.670 ;
        RECT 234.240 17.350 234.500 17.670 ;
        RECT 228.780 2.400 228.920 17.350 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 50.210 16.900 50.530 16.960 ;
        RECT 54.810 16.900 55.130 16.960 ;
        RECT 50.210 16.760 55.130 16.900 ;
        RECT 50.210 16.700 50.530 16.760 ;
        RECT 54.810 16.700 55.130 16.760 ;
      LAYER via ;
        RECT 50.240 16.700 50.500 16.960 ;
        RECT 54.840 16.700 55.100 16.960 ;
      LAYER met2 ;
        RECT 54.900 16.990 55.040 54.000 ;
        RECT 50.240 16.670 50.500 16.990 ;
        RECT 54.840 16.670 55.100 16.990 ;
        RECT 50.300 2.400 50.440 16.670 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 252.610 20.640 252.930 20.700 ;
        RECT 254.910 20.640 255.230 20.700 ;
        RECT 252.610 20.500 255.230 20.640 ;
        RECT 252.610 20.440 252.930 20.500 ;
        RECT 254.910 20.440 255.230 20.500 ;
      LAYER via ;
        RECT 252.640 20.440 252.900 20.700 ;
        RECT 254.940 20.440 255.200 20.700 ;
      LAYER met2 ;
        RECT 255.000 20.730 255.140 54.000 ;
        RECT 252.640 20.410 252.900 20.730 ;
        RECT 254.940 20.410 255.200 20.730 ;
        RECT 252.700 2.400 252.840 20.410 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 270.090 17.920 270.410 17.980 ;
        RECT 275.610 17.920 275.930 17.980 ;
        RECT 270.090 17.780 275.930 17.920 ;
        RECT 270.090 17.720 270.410 17.780 ;
        RECT 275.610 17.720 275.930 17.780 ;
      LAYER via ;
        RECT 270.120 17.720 270.380 17.980 ;
        RECT 275.640 17.720 275.900 17.980 ;
      LAYER met2 ;
        RECT 275.700 18.010 275.840 54.000 ;
        RECT 270.120 17.690 270.380 18.010 ;
        RECT 275.640 17.690 275.900 18.010 ;
        RECT 270.180 2.400 270.320 17.690 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 289.500 3.130 289.640 54.000 ;
        RECT 288.120 2.990 289.640 3.130 ;
        RECT 288.120 2.400 288.260 2.990 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 305.970 17.920 306.290 17.980 ;
        RECT 310.110 17.920 310.430 17.980 ;
        RECT 305.970 17.780 310.430 17.920 ;
        RECT 305.970 17.720 306.290 17.780 ;
        RECT 310.110 17.720 310.430 17.780 ;
      LAYER via ;
        RECT 306.000 17.720 306.260 17.980 ;
        RECT 310.140 17.720 310.400 17.980 ;
      LAYER met2 ;
        RECT 310.200 18.010 310.340 54.000 ;
        RECT 306.000 17.690 306.260 18.010 ;
        RECT 310.140 17.690 310.400 18.010 ;
        RECT 306.060 2.400 306.200 17.690 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.450 19.960 323.770 20.020 ;
        RECT 341.390 19.960 341.710 20.020 ;
        RECT 323.450 19.820 341.710 19.960 ;
        RECT 323.450 19.760 323.770 19.820 ;
        RECT 341.390 19.760 341.710 19.820 ;
      LAYER via ;
        RECT 323.480 19.760 323.740 20.020 ;
        RECT 341.420 19.760 341.680 20.020 ;
      LAYER met2 ;
        RECT 341.480 20.050 341.620 54.000 ;
        RECT 323.480 19.730 323.740 20.050 ;
        RECT 341.420 19.730 341.680 20.050 ;
        RECT 323.540 9.930 323.680 19.730 ;
        RECT 323.540 9.790 324.140 9.930 ;
        RECT 324.000 2.400 324.140 9.790 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 341.390 16.900 341.710 16.960 ;
        RECT 344.610 16.900 344.930 16.960 ;
        RECT 341.390 16.760 344.930 16.900 ;
        RECT 341.390 16.700 341.710 16.760 ;
        RECT 344.610 16.700 344.930 16.760 ;
      LAYER via ;
        RECT 341.420 16.700 341.680 16.960 ;
        RECT 344.640 16.700 344.900 16.960 ;
      LAYER met2 ;
        RECT 344.700 16.990 344.840 54.000 ;
        RECT 341.420 16.670 341.680 16.990 ;
        RECT 344.640 16.670 344.900 16.990 ;
        RECT 341.480 2.400 341.620 16.670 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 359.330 20.640 359.650 20.700 ;
        RECT 365.310 20.640 365.630 20.700 ;
        RECT 359.330 20.500 365.630 20.640 ;
        RECT 359.330 20.440 359.650 20.500 ;
        RECT 365.310 20.440 365.630 20.500 ;
      LAYER via ;
        RECT 359.360 20.440 359.620 20.700 ;
        RECT 365.340 20.440 365.600 20.700 ;
      LAYER met2 ;
        RECT 365.400 20.730 365.540 54.000 ;
        RECT 359.360 20.410 359.620 20.730 ;
        RECT 365.340 20.410 365.600 20.730 ;
        RECT 359.420 2.400 359.560 20.410 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 379.200 3.130 379.340 54.000 ;
        RECT 377.360 2.990 379.340 3.130 ;
        RECT 377.360 2.400 377.500 2.990 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 395.210 20.640 395.530 20.700 ;
        RECT 399.810 20.640 400.130 20.700 ;
        RECT 395.210 20.500 400.130 20.640 ;
        RECT 395.210 20.440 395.530 20.500 ;
        RECT 399.810 20.440 400.130 20.500 ;
      LAYER via ;
        RECT 395.240 20.440 395.500 20.700 ;
        RECT 399.840 20.440 400.100 20.700 ;
      LAYER met2 ;
        RECT 399.900 20.730 400.040 54.000 ;
        RECT 395.240 20.410 395.500 20.730 ;
        RECT 399.840 20.410 400.100 20.730 ;
        RECT 395.300 2.400 395.440 20.410 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.700 17.410 413.840 54.000 ;
        RECT 413.240 17.270 413.840 17.410 ;
        RECT 413.240 2.400 413.380 17.270 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.600 17.410 75.740 54.000 ;
        RECT 74.220 17.270 75.740 17.410 ;
        RECT 74.220 2.400 74.360 17.270 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 430.630 17.920 430.950 17.980 ;
        RECT 434.310 17.920 434.630 17.980 ;
        RECT 430.630 17.780 434.630 17.920 ;
        RECT 430.630 17.720 430.950 17.780 ;
        RECT 434.310 17.720 434.630 17.780 ;
      LAYER via ;
        RECT 430.660 17.720 430.920 17.980 ;
        RECT 434.340 17.720 434.600 17.980 ;
      LAYER met2 ;
        RECT 434.400 18.010 434.540 54.000 ;
        RECT 430.660 17.690 430.920 18.010 ;
        RECT 434.340 17.690 434.600 18.010 ;
        RECT 430.720 2.400 430.860 17.690 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 448.570 17.920 448.890 17.980 ;
        RECT 455.010 17.920 455.330 17.980 ;
        RECT 448.570 17.780 455.330 17.920 ;
        RECT 448.570 17.720 448.890 17.780 ;
        RECT 455.010 17.720 455.330 17.780 ;
      LAYER via ;
        RECT 448.600 17.720 448.860 17.980 ;
        RECT 455.040 17.720 455.300 17.980 ;
      LAYER met2 ;
        RECT 455.100 18.010 455.240 54.000 ;
        RECT 448.600 17.690 448.860 18.010 ;
        RECT 455.040 17.690 455.300 18.010 ;
        RECT 448.660 2.400 448.800 17.690 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 466.510 16.900 466.830 16.960 ;
        RECT 468.810 16.900 469.130 16.960 ;
        RECT 466.510 16.760 469.130 16.900 ;
        RECT 466.510 16.700 466.830 16.760 ;
        RECT 468.810 16.700 469.130 16.760 ;
      LAYER via ;
        RECT 466.540 16.700 466.800 16.960 ;
        RECT 468.840 16.700 469.100 16.960 ;
      LAYER met2 ;
        RECT 468.900 16.990 469.040 54.000 ;
        RECT 466.540 16.670 466.800 16.990 ;
        RECT 468.840 16.670 469.100 16.990 ;
        RECT 466.600 2.400 466.740 16.670 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 484.450 16.900 484.770 16.960 ;
        RECT 489.510 16.900 489.830 16.960 ;
        RECT 484.450 16.760 489.830 16.900 ;
        RECT 484.450 16.700 484.770 16.760 ;
        RECT 489.510 16.700 489.830 16.760 ;
      LAYER via ;
        RECT 484.480 16.700 484.740 16.960 ;
        RECT 489.540 16.700 489.800 16.960 ;
      LAYER met2 ;
        RECT 489.600 16.990 489.740 54.000 ;
        RECT 484.480 16.670 484.740 16.990 ;
        RECT 489.540 16.670 489.800 16.990 ;
        RECT 484.540 2.400 484.680 16.670 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 503.400 16.730 503.540 54.000 ;
        RECT 502.480 16.590 503.540 16.730 ;
        RECT 502.480 2.400 502.620 16.590 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 519.870 17.580 520.190 17.640 ;
        RECT 524.010 17.580 524.330 17.640 ;
        RECT 519.870 17.440 524.330 17.580 ;
        RECT 519.870 17.380 520.190 17.440 ;
        RECT 524.010 17.380 524.330 17.440 ;
      LAYER via ;
        RECT 519.900 17.380 520.160 17.640 ;
        RECT 524.040 17.380 524.300 17.640 ;
      LAYER met2 ;
        RECT 524.100 17.670 524.240 54.000 ;
        RECT 519.900 17.350 520.160 17.670 ;
        RECT 524.040 17.350 524.300 17.670 ;
        RECT 519.960 2.400 520.100 17.350 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.440 17.410 537.580 54.000 ;
        RECT 537.440 17.270 538.040 17.410 ;
        RECT 537.900 2.400 538.040 17.270 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 555.750 20.640 556.070 20.700 ;
        RECT 558.510 20.640 558.830 20.700 ;
        RECT 555.750 20.500 558.830 20.640 ;
        RECT 555.750 20.440 556.070 20.500 ;
        RECT 558.510 20.440 558.830 20.500 ;
      LAYER via ;
        RECT 555.780 20.440 556.040 20.700 ;
        RECT 558.540 20.440 558.800 20.700 ;
      LAYER met2 ;
        RECT 558.600 20.730 558.740 54.000 ;
        RECT 555.780 20.410 556.040 20.730 ;
        RECT 558.540 20.410 558.800 20.730 ;
        RECT 555.840 2.400 555.980 20.410 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 573.690 17.580 574.010 17.640 ;
        RECT 579.210 17.580 579.530 17.640 ;
        RECT 573.690 17.440 579.530 17.580 ;
        RECT 573.690 17.380 574.010 17.440 ;
        RECT 579.210 17.380 579.530 17.440 ;
      LAYER via ;
        RECT 573.720 17.380 573.980 17.640 ;
        RECT 579.240 17.380 579.500 17.640 ;
      LAYER met2 ;
        RECT 579.300 17.670 579.440 54.000 ;
        RECT 573.720 17.350 573.980 17.670 ;
        RECT 579.240 17.350 579.500 17.670 ;
        RECT 573.780 2.400 573.920 17.350 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 591.170 14.180 591.490 14.240 ;
        RECT 593.010 14.180 593.330 14.240 ;
        RECT 591.170 14.040 593.330 14.180 ;
        RECT 591.170 13.980 591.490 14.040 ;
        RECT 593.010 13.980 593.330 14.040 ;
      LAYER via ;
        RECT 591.200 13.980 591.460 14.240 ;
        RECT 593.040 13.980 593.300 14.240 ;
      LAYER met2 ;
        RECT 593.100 14.270 593.240 54.000 ;
        RECT 591.200 13.950 591.460 14.270 ;
        RECT 593.040 13.950 593.300 14.270 ;
        RECT 591.260 2.400 591.400 13.950 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 97.590 19.620 97.910 19.680 ;
        RECT 203.390 19.620 203.710 19.680 ;
        RECT 97.590 19.480 203.710 19.620 ;
        RECT 97.590 19.420 97.910 19.480 ;
        RECT 203.390 19.420 203.710 19.480 ;
      LAYER via ;
        RECT 97.620 19.420 97.880 19.680 ;
        RECT 203.420 19.420 203.680 19.680 ;
      LAYER met2 ;
        RECT 203.480 19.710 203.620 54.000 ;
        RECT 97.620 19.390 97.880 19.710 ;
        RECT 203.420 19.390 203.680 19.710 ;
        RECT 97.680 2.400 97.820 19.390 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 609.110 17.920 609.430 17.980 ;
        RECT 613.710 17.920 614.030 17.980 ;
        RECT 609.110 17.780 614.030 17.920 ;
        RECT 609.110 17.720 609.430 17.780 ;
        RECT 613.710 17.720 614.030 17.780 ;
      LAYER via ;
        RECT 609.140 17.720 609.400 17.980 ;
        RECT 613.740 17.720 614.000 17.980 ;
      LAYER met2 ;
        RECT 613.800 18.010 613.940 54.000 ;
        RECT 609.140 17.690 609.400 18.010 ;
        RECT 613.740 17.690 614.000 18.010 ;
        RECT 609.200 2.400 609.340 17.690 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 627.140 2.400 627.280 54.000 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 16.900 121.830 16.960 ;
        RECT 123.810 16.900 124.130 16.960 ;
        RECT 121.510 16.760 124.130 16.900 ;
        RECT 121.510 16.700 121.830 16.760 ;
        RECT 123.810 16.700 124.130 16.760 ;
      LAYER via ;
        RECT 121.540 16.700 121.800 16.960 ;
        RECT 123.840 16.700 124.100 16.960 ;
      LAYER met2 ;
        RECT 123.900 16.990 124.040 54.000 ;
        RECT 121.540 16.670 121.800 16.990 ;
        RECT 123.840 16.670 124.100 16.990 ;
        RECT 121.600 2.400 121.740 16.670 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 145.430 18.940 145.750 19.000 ;
        RECT 299.990 18.940 300.310 19.000 ;
        RECT 145.430 18.800 300.310 18.940 ;
        RECT 145.430 18.740 145.750 18.800 ;
        RECT 299.990 18.740 300.310 18.800 ;
      LAYER via ;
        RECT 145.460 18.740 145.720 19.000 ;
        RECT 300.020 18.740 300.280 19.000 ;
      LAYER met2 ;
        RECT 300.080 19.030 300.220 54.000 ;
        RECT 145.460 18.710 145.720 19.030 ;
        RECT 300.020 18.710 300.280 19.030 ;
        RECT 145.520 2.400 145.660 18.710 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 165.300 17.410 165.440 54.000 ;
        RECT 163.460 17.270 165.440 17.410 ;
        RECT 163.460 2.400 163.600 17.270 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 180.850 19.280 181.170 19.340 ;
        RECT 320.690 19.280 321.010 19.340 ;
        RECT 180.850 19.140 321.010 19.280 ;
        RECT 180.850 19.080 181.170 19.140 ;
        RECT 320.690 19.080 321.010 19.140 ;
      LAYER via ;
        RECT 180.880 19.080 181.140 19.340 ;
        RECT 320.720 19.080 320.980 19.340 ;
      LAYER met2 ;
        RECT 320.780 19.370 320.920 54.000 ;
        RECT 180.880 19.050 181.140 19.370 ;
        RECT 320.720 19.050 320.980 19.370 ;
        RECT 180.940 2.400 181.080 19.050 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 199.800 3.130 199.940 54.000 ;
        RECT 198.880 2.990 199.940 3.130 ;
        RECT 198.880 2.400 199.020 2.990 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 375.430 17.580 375.750 17.640 ;
        RECT 234.760 17.440 375.750 17.580 ;
        RECT 216.730 17.240 217.050 17.300 ;
        RECT 234.760 17.240 234.900 17.440 ;
        RECT 375.430 17.380 375.750 17.440 ;
        RECT 216.730 17.100 234.900 17.240 ;
        RECT 216.730 17.040 217.050 17.100 ;
      LAYER via ;
        RECT 216.760 17.040 217.020 17.300 ;
        RECT 375.460 17.380 375.720 17.640 ;
      LAYER met2 ;
        RECT 375.980 20.130 376.120 54.000 ;
        RECT 375.520 19.990 376.120 20.130 ;
        RECT 375.520 17.670 375.660 19.990 ;
        RECT 375.460 17.350 375.720 17.670 ;
        RECT 216.760 17.010 217.020 17.330 ;
        RECT 216.820 2.400 216.960 17.010 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 383.250 19.960 383.570 20.020 ;
        RECT 367.700 19.820 383.570 19.960 ;
        RECT 234.670 19.620 234.990 19.680 ;
        RECT 367.700 19.620 367.840 19.820 ;
        RECT 383.250 19.760 383.570 19.820 ;
        RECT 234.670 19.480 367.840 19.620 ;
        RECT 234.670 19.420 234.990 19.480 ;
      LAYER via ;
        RECT 234.700 19.420 234.960 19.680 ;
        RECT 383.280 19.760 383.540 20.020 ;
      LAYER met2 ;
        RECT 383.340 20.050 383.480 54.000 ;
        RECT 383.280 19.730 383.540 20.050 ;
        RECT 234.700 19.390 234.960 19.710 ;
        RECT 234.760 2.400 234.900 19.390 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 56.190 18.600 56.510 18.660 ;
        RECT 217.190 18.600 217.510 18.660 ;
        RECT 56.190 18.460 217.510 18.600 ;
        RECT 56.190 18.400 56.510 18.460 ;
        RECT 217.190 18.400 217.510 18.460 ;
      LAYER via ;
        RECT 56.220 18.400 56.480 18.660 ;
        RECT 217.220 18.400 217.480 18.660 ;
      LAYER met2 ;
        RECT 217.280 18.690 217.420 54.000 ;
        RECT 56.220 18.370 56.480 18.690 ;
        RECT 217.220 18.370 217.480 18.690 ;
        RECT 56.280 2.400 56.420 18.370 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 80.110 16.900 80.430 16.960 ;
        RECT 82.410 16.900 82.730 16.960 ;
        RECT 80.110 16.760 82.730 16.900 ;
        RECT 80.110 16.700 80.430 16.760 ;
        RECT 82.410 16.700 82.730 16.760 ;
      LAYER via ;
        RECT 80.140 16.700 80.400 16.960 ;
        RECT 82.440 16.700 82.700 16.960 ;
      LAYER met2 ;
        RECT 82.500 16.990 82.640 54.000 ;
        RECT 80.140 16.670 80.400 16.990 ;
        RECT 82.440 16.670 82.700 16.990 ;
        RECT 80.200 2.400 80.340 16.670 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 103.570 19.960 103.890 20.020 ;
        RECT 237.890 19.960 238.210 20.020 ;
        RECT 103.570 19.820 238.210 19.960 ;
        RECT 103.570 19.760 103.890 19.820 ;
        RECT 237.890 19.760 238.210 19.820 ;
      LAYER via ;
        RECT 103.600 19.760 103.860 20.020 ;
        RECT 237.920 19.760 238.180 20.020 ;
      LAYER met2 ;
        RECT 237.980 20.050 238.120 54.000 ;
        RECT 103.600 19.730 103.860 20.050 ;
        RECT 237.920 19.730 238.180 20.050 ;
        RECT 103.660 2.400 103.800 19.730 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 127.490 16.900 127.810 16.960 ;
        RECT 130.710 16.900 131.030 16.960 ;
        RECT 127.490 16.760 131.030 16.900 ;
        RECT 127.490 16.700 127.810 16.760 ;
        RECT 130.710 16.700 131.030 16.760 ;
      LAYER via ;
        RECT 127.520 16.700 127.780 16.960 ;
        RECT 130.740 16.700 131.000 16.960 ;
      LAYER met2 ;
        RECT 130.800 16.990 130.940 54.000 ;
        RECT 127.520 16.670 127.780 16.990 ;
        RECT 130.740 16.670 131.000 16.990 ;
        RECT 127.580 2.400 127.720 16.670 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.290 18.260 26.610 18.320 ;
        RECT 214.890 18.260 215.210 18.320 ;
        RECT 26.290 18.120 215.210 18.260 ;
        RECT 26.290 18.060 26.610 18.120 ;
        RECT 214.890 18.060 215.210 18.120 ;
      LAYER via ;
        RECT 26.320 18.060 26.580 18.320 ;
        RECT 214.920 18.060 215.180 18.320 ;
      LAYER met2 ;
        RECT 214.980 18.350 215.120 54.000 ;
        RECT 26.320 18.030 26.580 18.350 ;
        RECT 214.920 18.030 215.180 18.350 ;
        RECT 26.380 2.400 26.520 18.030 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 34.110 307.260 34.430 307.320 ;
        RECT 34.110 307.120 54.000 307.260 ;
        RECT 34.110 307.060 34.430 307.120 ;
      LAYER via ;
        RECT 34.140 307.060 34.400 307.320 ;
      LAYER met2 ;
        RECT 34.140 307.030 34.400 307.350 ;
        RECT 34.200 3.130 34.340 307.030 ;
        RECT 32.360 2.990 34.340 3.130 ;
        RECT 32.360 2.400 32.500 2.990 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 184.020 3466.000 187.020 3529.000 ;
        RECT 364.020 3466.000 367.020 3529.000 ;
        RECT 544.020 3466.000 547.020 3529.000 ;
        RECT 724.020 3466.000 727.020 3529.000 ;
        RECT 904.020 3466.000 907.020 3529.000 ;
        RECT 1084.020 3466.000 1087.020 3529.000 ;
        RECT 1264.020 3466.000 1267.020 3529.000 ;
        RECT 1444.020 3466.000 1447.020 3529.000 ;
        RECT 1624.020 3466.000 1627.020 3529.000 ;
        RECT 1804.020 3466.000 1807.020 3529.000 ;
        RECT 1984.020 3466.000 1987.020 3529.000 ;
        RECT 2164.020 3466.000 2167.020 3529.000 ;
        RECT 2344.020 3466.000 2347.020 3529.000 ;
        RECT 2524.020 3466.000 2527.020 3529.000 ;
        RECT 2704.020 3466.000 2707.020 3529.000 ;
        RECT 184.020 -9.320 187.020 54.000 ;
        RECT 364.020 -9.320 367.020 54.000 ;
        RECT 544.020 -9.320 547.020 54.000 ;
        RECT 724.020 -9.320 727.020 54.000 ;
        RECT 904.020 -9.320 907.020 54.000 ;
        RECT 1084.020 -9.320 1087.020 54.000 ;
        RECT 1264.020 -9.320 1267.020 54.000 ;
        RECT 1444.020 -9.320 1447.020 54.000 ;
        RECT 1624.020 -9.320 1627.020 54.000 ;
        RECT 1804.020 -9.320 1807.020 54.000 ;
        RECT 1984.020 -9.320 1987.020 54.000 ;
        RECT 2164.020 -9.320 2167.020 54.000 ;
        RECT 2344.020 -9.320 2347.020 54.000 ;
        RECT 2524.020 -9.320 2527.020 54.000 ;
        RECT 2704.020 -9.320 2707.020 54.000 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 54.000 3432.380 ;
        RECT 2866.000 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 54.000 3252.380 ;
        RECT 2866.000 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 54.000 3072.380 ;
        RECT 2866.000 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 54.000 2892.380 ;
        RECT 2866.000 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 54.000 2712.380 ;
        RECT 2866.000 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 54.000 2532.380 ;
        RECT 2866.000 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 54.000 2352.380 ;
        RECT 2866.000 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 54.000 2172.380 ;
        RECT 2866.000 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 54.000 1992.380 ;
        RECT 2866.000 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 54.000 1812.380 ;
        RECT 2866.000 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 54.000 1632.380 ;
        RECT 2866.000 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 54.000 1452.380 ;
        RECT 2866.000 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 54.000 1272.380 ;
        RECT 2866.000 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 54.000 1092.380 ;
        RECT 2866.000 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 54.000 912.380 ;
        RECT 2866.000 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 54.000 732.380 ;
        RECT 2866.000 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 54.000 552.380 ;
        RECT 2866.000 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 54.000 372.380 ;
        RECT 2866.000 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 54.000 192.380 ;
        RECT 2866.000 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 3466.000 97.020 3529.000 ;
        RECT 274.020 3466.000 277.020 3529.000 ;
        RECT 454.020 3466.000 457.020 3529.000 ;
        RECT 634.020 3466.000 637.020 3529.000 ;
        RECT 814.020 3466.000 817.020 3529.000 ;
        RECT 994.020 3466.000 997.020 3529.000 ;
        RECT 1174.020 3466.000 1177.020 3529.000 ;
        RECT 1354.020 3466.000 1357.020 3529.000 ;
        RECT 1534.020 3466.000 1537.020 3529.000 ;
        RECT 1714.020 3466.000 1717.020 3529.000 ;
        RECT 1894.020 3466.000 1897.020 3529.000 ;
        RECT 2074.020 3466.000 2077.020 3529.000 ;
        RECT 2254.020 3466.000 2257.020 3529.000 ;
        RECT 2434.020 3466.000 2437.020 3529.000 ;
        RECT 2614.020 3466.000 2617.020 3529.000 ;
        RECT 2794.020 3466.000 2797.020 3529.000 ;
        RECT 94.020 -9.320 97.020 54.000 ;
        RECT 274.020 -9.320 277.020 54.000 ;
        RECT 454.020 -9.320 457.020 54.000 ;
        RECT 634.020 -9.320 637.020 54.000 ;
        RECT 814.020 -9.320 817.020 54.000 ;
        RECT 994.020 -9.320 997.020 54.000 ;
        RECT 1174.020 -9.320 1177.020 54.000 ;
        RECT 1354.020 -9.320 1357.020 54.000 ;
        RECT 1534.020 -9.320 1537.020 54.000 ;
        RECT 1714.020 -9.320 1717.020 54.000 ;
        RECT 1894.020 -9.320 1897.020 54.000 ;
        RECT 2074.020 -9.320 2077.020 54.000 ;
        RECT 2254.020 -9.320 2257.020 54.000 ;
        RECT 2434.020 -9.320 2437.020 54.000 ;
        RECT 2614.020 -9.320 2617.020 54.000 ;
        RECT 2794.020 -9.320 2797.020 54.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 54.000 3342.380 ;
        RECT 2866.000 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 54.000 3162.380 ;
        RECT 2866.000 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 54.000 2982.380 ;
        RECT 2866.000 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 54.000 2802.380 ;
        RECT 2866.000 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 54.000 2622.380 ;
        RECT 2866.000 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 54.000 2442.380 ;
        RECT 2866.000 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 54.000 2262.380 ;
        RECT 2866.000 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 54.000 2082.380 ;
        RECT 2866.000 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 54.000 1902.380 ;
        RECT 2866.000 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 54.000 1722.380 ;
        RECT 2866.000 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 54.000 1542.380 ;
        RECT 2866.000 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 54.000 1362.380 ;
        RECT 2866.000 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 54.000 1182.380 ;
        RECT 2866.000 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 54.000 1002.380 ;
        RECT 2866.000 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 54.000 822.380 ;
        RECT 2866.000 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 54.000 642.380 ;
        RECT 2866.000 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 54.000 462.380 ;
        RECT 2866.000 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 54.000 282.380 ;
        RECT 2866.000 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 54.000 102.380 ;
        RECT 2866.000 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 202.020 3466.000 205.020 3538.400 ;
        RECT 382.020 3466.000 385.020 3538.400 ;
        RECT 562.020 3466.000 565.020 3538.400 ;
        RECT 742.020 3466.000 745.020 3538.400 ;
        RECT 922.020 3466.000 925.020 3538.400 ;
        RECT 1102.020 3466.000 1105.020 3538.400 ;
        RECT 1282.020 3466.000 1285.020 3538.400 ;
        RECT 1462.020 3466.000 1465.020 3538.400 ;
        RECT 1642.020 3466.000 1645.020 3538.400 ;
        RECT 1822.020 3466.000 1825.020 3538.400 ;
        RECT 2002.020 3466.000 2005.020 3538.400 ;
        RECT 2182.020 3466.000 2185.020 3538.400 ;
        RECT 2362.020 3466.000 2365.020 3538.400 ;
        RECT 2542.020 3466.000 2545.020 3538.400 ;
        RECT 2722.020 3466.000 2725.020 3538.400 ;
        RECT 202.020 -18.720 205.020 54.000 ;
        RECT 382.020 -18.720 385.020 54.000 ;
        RECT 562.020 -18.720 565.020 54.000 ;
        RECT 742.020 -18.720 745.020 54.000 ;
        RECT 922.020 -18.720 925.020 54.000 ;
        RECT 1102.020 -18.720 1105.020 54.000 ;
        RECT 1282.020 -18.720 1285.020 54.000 ;
        RECT 1462.020 -18.720 1465.020 54.000 ;
        RECT 1642.020 -18.720 1645.020 54.000 ;
        RECT 1822.020 -18.720 1825.020 54.000 ;
        RECT 2002.020 -18.720 2005.020 54.000 ;
        RECT 2182.020 -18.720 2185.020 54.000 ;
        RECT 2362.020 -18.720 2365.020 54.000 ;
        RECT 2542.020 -18.720 2545.020 54.000 ;
        RECT 2722.020 -18.720 2725.020 54.000 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 54.000 3450.380 ;
        RECT 2866.000 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 54.000 3270.380 ;
        RECT 2866.000 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 54.000 3090.380 ;
        RECT 2866.000 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 54.000 2910.380 ;
        RECT 2866.000 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 54.000 2730.380 ;
        RECT 2866.000 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 54.000 2550.380 ;
        RECT 2866.000 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 54.000 2370.380 ;
        RECT 2866.000 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 54.000 2190.380 ;
        RECT 2866.000 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 54.000 2010.380 ;
        RECT 2866.000 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 54.000 1830.380 ;
        RECT 2866.000 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 54.000 1650.380 ;
        RECT 2866.000 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 54.000 1470.380 ;
        RECT 2866.000 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 54.000 1290.380 ;
        RECT 2866.000 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 54.000 1110.380 ;
        RECT 2866.000 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 54.000 930.380 ;
        RECT 2866.000 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 54.000 750.380 ;
        RECT 2866.000 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 54.000 570.380 ;
        RECT 2866.000 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 54.000 390.380 ;
        RECT 2866.000 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 54.000 210.380 ;
        RECT 2866.000 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 112.020 3466.000 115.020 3538.400 ;
        RECT 292.020 3466.000 295.020 3538.400 ;
        RECT 472.020 3466.000 475.020 3538.400 ;
        RECT 652.020 3466.000 655.020 3538.400 ;
        RECT 832.020 3466.000 835.020 3538.400 ;
        RECT 1012.020 3466.000 1015.020 3538.400 ;
        RECT 1192.020 3466.000 1195.020 3538.400 ;
        RECT 1372.020 3466.000 1375.020 3538.400 ;
        RECT 1552.020 3466.000 1555.020 3538.400 ;
        RECT 1732.020 3466.000 1735.020 3538.400 ;
        RECT 1912.020 3466.000 1915.020 3538.400 ;
        RECT 2092.020 3466.000 2095.020 3538.400 ;
        RECT 2272.020 3466.000 2275.020 3538.400 ;
        RECT 2452.020 3466.000 2455.020 3538.400 ;
        RECT 2632.020 3466.000 2635.020 3538.400 ;
        RECT 2812.020 3466.000 2815.020 3538.400 ;
        RECT 112.020 -18.720 115.020 54.000 ;
        RECT 292.020 -18.720 295.020 54.000 ;
        RECT 472.020 -18.720 475.020 54.000 ;
        RECT 652.020 -18.720 655.020 54.000 ;
        RECT 832.020 -18.720 835.020 54.000 ;
        RECT 1012.020 -18.720 1015.020 54.000 ;
        RECT 1192.020 -18.720 1195.020 54.000 ;
        RECT 1372.020 -18.720 1375.020 54.000 ;
        RECT 1552.020 -18.720 1555.020 54.000 ;
        RECT 1732.020 -18.720 1735.020 54.000 ;
        RECT 1912.020 -18.720 1915.020 54.000 ;
        RECT 2092.020 -18.720 2095.020 54.000 ;
        RECT 2272.020 -18.720 2275.020 54.000 ;
        RECT 2452.020 -18.720 2455.020 54.000 ;
        RECT 2632.020 -18.720 2635.020 54.000 ;
        RECT 2812.020 -18.720 2815.020 54.000 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 54.000 3360.380 ;
        RECT 2866.000 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 54.000 3180.380 ;
        RECT 2866.000 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 54.000 3000.380 ;
        RECT 2866.000 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 54.000 2820.380 ;
        RECT 2866.000 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 54.000 2640.380 ;
        RECT 2866.000 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 54.000 2460.380 ;
        RECT 2866.000 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 54.000 2280.380 ;
        RECT 2866.000 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 54.000 2100.380 ;
        RECT 2866.000 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 54.000 1920.380 ;
        RECT 2866.000 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 54.000 1740.380 ;
        RECT 2866.000 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 54.000 1560.380 ;
        RECT 2866.000 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 54.000 1380.380 ;
        RECT 2866.000 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 54.000 1200.380 ;
        RECT 2866.000 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 54.000 1020.380 ;
        RECT 2866.000 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 54.000 840.380 ;
        RECT 2866.000 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 54.000 660.380 ;
        RECT 2866.000 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 54.000 480.380 ;
        RECT 2866.000 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 54.000 300.380 ;
        RECT 2866.000 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 54.000 120.380 ;
        RECT 2866.000 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 220.020 3466.000 223.020 3547.800 ;
        RECT 400.020 3466.000 403.020 3547.800 ;
        RECT 580.020 3466.000 583.020 3547.800 ;
        RECT 760.020 3466.000 763.020 3547.800 ;
        RECT 940.020 3466.000 943.020 3547.800 ;
        RECT 1120.020 3466.000 1123.020 3547.800 ;
        RECT 1300.020 3466.000 1303.020 3547.800 ;
        RECT 1480.020 3466.000 1483.020 3547.800 ;
        RECT 1660.020 3466.000 1663.020 3547.800 ;
        RECT 1840.020 3466.000 1843.020 3547.800 ;
        RECT 2020.020 3466.000 2023.020 3547.800 ;
        RECT 2200.020 3466.000 2203.020 3547.800 ;
        RECT 2380.020 3466.000 2383.020 3547.800 ;
        RECT 2560.020 3466.000 2563.020 3547.800 ;
        RECT 2740.020 3466.000 2743.020 3547.800 ;
        RECT 220.020 -28.120 223.020 54.000 ;
        RECT 400.020 -28.120 403.020 54.000 ;
        RECT 580.020 -28.120 583.020 54.000 ;
        RECT 760.020 -28.120 763.020 54.000 ;
        RECT 940.020 -28.120 943.020 54.000 ;
        RECT 1120.020 -28.120 1123.020 54.000 ;
        RECT 1300.020 -28.120 1303.020 54.000 ;
        RECT 1480.020 -28.120 1483.020 54.000 ;
        RECT 1660.020 -28.120 1663.020 54.000 ;
        RECT 1840.020 -28.120 1843.020 54.000 ;
        RECT 2020.020 -28.120 2023.020 54.000 ;
        RECT 2200.020 -28.120 2203.020 54.000 ;
        RECT 2380.020 -28.120 2383.020 54.000 ;
        RECT 2560.020 -28.120 2563.020 54.000 ;
        RECT 2740.020 -28.120 2743.020 54.000 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3466.000 222.110 3466.670 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3466.000 402.110 3466.670 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3466.000 582.110 3466.670 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3466.000 762.110 3466.670 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3466.000 942.110 3466.670 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3466.000 1122.110 3466.670 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3466.000 1302.110 3466.670 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3466.000 1482.110 3466.670 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3466.000 1662.110 3466.670 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3466.000 1842.110 3466.670 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3466.000 2022.110 3466.670 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3466.000 2202.110 3466.670 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3466.000 2382.110 3466.670 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3466.000 2562.110 3466.670 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3466.000 2742.110 3466.670 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3466.000 2953.100 3468.380 ;
        RECT -33.480 3465.380 54.000 3466.000 ;
        RECT 2866.000 3465.380 2953.100 3466.000 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 54.000 3288.380 ;
        RECT 2866.000 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 54.000 3108.380 ;
        RECT 2866.000 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 54.000 2928.380 ;
        RECT 2866.000 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 54.000 2748.380 ;
        RECT 2866.000 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 54.000 2568.380 ;
        RECT 2866.000 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 54.000 2388.380 ;
        RECT 2866.000 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 54.000 2208.380 ;
        RECT 2866.000 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 54.000 2028.380 ;
        RECT 2866.000 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 54.000 1848.380 ;
        RECT 2866.000 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 54.000 1668.380 ;
        RECT 2866.000 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 54.000 1488.380 ;
        RECT 2866.000 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 54.000 1308.380 ;
        RECT 2866.000 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 54.000 1128.380 ;
        RECT 2866.000 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 54.000 948.380 ;
        RECT 2866.000 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 54.000 768.380 ;
        RECT 2866.000 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 54.000 588.380 ;
        RECT 2866.000 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 54.000 408.380 ;
        RECT 2866.000 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 54.000 228.380 ;
        RECT 2866.000 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 130.020 3466.000 133.020 3547.800 ;
        RECT 310.020 3466.000 313.020 3547.800 ;
        RECT 490.020 3466.000 493.020 3547.800 ;
        RECT 670.020 3466.000 673.020 3547.800 ;
        RECT 850.020 3466.000 853.020 3547.800 ;
        RECT 1030.020 3466.000 1033.020 3547.800 ;
        RECT 1210.020 3466.000 1213.020 3547.800 ;
        RECT 1390.020 3466.000 1393.020 3547.800 ;
        RECT 1570.020 3466.000 1573.020 3547.800 ;
        RECT 1750.020 3466.000 1753.020 3547.800 ;
        RECT 1930.020 3466.000 1933.020 3547.800 ;
        RECT 2110.020 3466.000 2113.020 3547.800 ;
        RECT 2290.020 3466.000 2293.020 3547.800 ;
        RECT 2470.020 3466.000 2473.020 3547.800 ;
        RECT 2650.020 3466.000 2653.020 3547.800 ;
        RECT 2830.020 3466.000 2833.020 3547.800 ;
        RECT 130.020 -28.120 133.020 54.000 ;
        RECT 310.020 -28.120 313.020 54.000 ;
        RECT 490.020 -28.120 493.020 54.000 ;
        RECT 670.020 -28.120 673.020 54.000 ;
        RECT 850.020 -28.120 853.020 54.000 ;
        RECT 1030.020 -28.120 1033.020 54.000 ;
        RECT 1210.020 -28.120 1213.020 54.000 ;
        RECT 1390.020 -28.120 1393.020 54.000 ;
        RECT 1570.020 -28.120 1573.020 54.000 ;
        RECT 1750.020 -28.120 1753.020 54.000 ;
        RECT 1930.020 -28.120 1933.020 54.000 ;
        RECT 2110.020 -28.120 2113.020 54.000 ;
        RECT 2290.020 -28.120 2293.020 54.000 ;
        RECT 2470.020 -28.120 2473.020 54.000 ;
        RECT 2650.020 -28.120 2653.020 54.000 ;
        RECT 2830.020 -28.120 2833.020 54.000 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 54.000 3378.380 ;
        RECT 2866.000 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 54.000 3198.380 ;
        RECT 2866.000 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 54.000 3018.380 ;
        RECT 2866.000 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 54.000 2838.380 ;
        RECT 2866.000 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 54.000 2658.380 ;
        RECT 2866.000 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 54.000 2478.380 ;
        RECT 2866.000 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 54.000 2298.380 ;
        RECT 2866.000 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 54.000 2118.380 ;
        RECT 2866.000 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 54.000 1938.380 ;
        RECT 2866.000 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 54.000 1758.380 ;
        RECT 2866.000 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 54.000 1578.380 ;
        RECT 2866.000 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 54.000 1398.380 ;
        RECT 2866.000 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 54.000 1218.380 ;
        RECT 2866.000 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 54.000 1038.380 ;
        RECT 2866.000 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 54.000 858.380 ;
        RECT 2866.000 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 54.000 678.380 ;
        RECT 2866.000 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 54.000 498.380 ;
        RECT 2866.000 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 54.000 318.380 ;
        RECT 2866.000 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 54.000 138.380 ;
        RECT 2866.000 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 58.020 3466.000 61.020 3557.200 ;
        RECT 238.020 3466.000 241.020 3557.200 ;
        RECT 418.020 3466.000 421.020 3557.200 ;
        RECT 598.020 3466.000 601.020 3557.200 ;
        RECT 778.020 3466.000 781.020 3557.200 ;
        RECT 958.020 3466.000 961.020 3557.200 ;
        RECT 1138.020 3466.000 1141.020 3557.200 ;
        RECT 1318.020 3466.000 1321.020 3557.200 ;
        RECT 1498.020 3466.000 1501.020 3557.200 ;
        RECT 1678.020 3466.000 1681.020 3557.200 ;
        RECT 1858.020 3466.000 1861.020 3557.200 ;
        RECT 2038.020 3466.000 2041.020 3557.200 ;
        RECT 2218.020 3466.000 2221.020 3557.200 ;
        RECT 2398.020 3466.000 2401.020 3557.200 ;
        RECT 2578.020 3466.000 2581.020 3557.200 ;
        RECT 2758.020 3466.000 2761.020 3557.200 ;
        RECT 58.020 -37.520 61.020 54.000 ;
        RECT 238.020 -37.520 241.020 54.000 ;
        RECT 418.020 -37.520 421.020 54.000 ;
        RECT 598.020 -37.520 601.020 54.000 ;
        RECT 778.020 -37.520 781.020 54.000 ;
        RECT 958.020 -37.520 961.020 54.000 ;
        RECT 1138.020 -37.520 1141.020 54.000 ;
        RECT 1318.020 -37.520 1321.020 54.000 ;
        RECT 1498.020 -37.520 1501.020 54.000 ;
        RECT 1678.020 -37.520 1681.020 54.000 ;
        RECT 1858.020 -37.520 1861.020 54.000 ;
        RECT 2038.020 -37.520 2041.020 54.000 ;
        RECT 2218.020 -37.520 2221.020 54.000 ;
        RECT 2398.020 -37.520 2401.020 54.000 ;
        RECT 2578.020 -37.520 2581.020 54.000 ;
        RECT 2758.020 -37.520 2761.020 54.000 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 54.000 3306.380 ;
        RECT 2866.000 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 54.000 3126.380 ;
        RECT 2866.000 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 54.000 2946.380 ;
        RECT 2866.000 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 54.000 2766.380 ;
        RECT 2866.000 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 54.000 2586.380 ;
        RECT 2866.000 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 54.000 2406.380 ;
        RECT 2866.000 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 54.000 2226.380 ;
        RECT 2866.000 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 54.000 2046.380 ;
        RECT 2866.000 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 54.000 1866.380 ;
        RECT 2866.000 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 54.000 1686.380 ;
        RECT 2866.000 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 54.000 1506.380 ;
        RECT 2866.000 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 54.000 1326.380 ;
        RECT 2866.000 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 54.000 1146.380 ;
        RECT 2866.000 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 54.000 966.380 ;
        RECT 2866.000 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 54.000 786.380 ;
        RECT 2866.000 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 54.000 606.380 ;
        RECT 2866.000 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 54.000 426.380 ;
        RECT 2866.000 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 54.000 246.380 ;
        RECT 2866.000 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 54.000 66.380 ;
        RECT 2866.000 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 148.020 3466.000 151.020 3557.200 ;
        RECT 328.020 3466.000 331.020 3557.200 ;
        RECT 508.020 3466.000 511.020 3557.200 ;
        RECT 688.020 3466.000 691.020 3557.200 ;
        RECT 868.020 3466.000 871.020 3557.200 ;
        RECT 1048.020 3466.000 1051.020 3557.200 ;
        RECT 1228.020 3466.000 1231.020 3557.200 ;
        RECT 1408.020 3466.000 1411.020 3557.200 ;
        RECT 1588.020 3466.000 1591.020 3557.200 ;
        RECT 1768.020 3466.000 1771.020 3557.200 ;
        RECT 1948.020 3466.000 1951.020 3557.200 ;
        RECT 2128.020 3466.000 2131.020 3557.200 ;
        RECT 2308.020 3466.000 2311.020 3557.200 ;
        RECT 2488.020 3466.000 2491.020 3557.200 ;
        RECT 2668.020 3466.000 2671.020 3557.200 ;
        RECT 2848.020 3466.000 2851.020 3557.200 ;
        RECT 148.020 -37.520 151.020 54.000 ;
        RECT 328.020 -37.520 331.020 54.000 ;
        RECT 508.020 -37.520 511.020 54.000 ;
        RECT 688.020 -37.520 691.020 54.000 ;
        RECT 868.020 -37.520 871.020 54.000 ;
        RECT 1048.020 -37.520 1051.020 54.000 ;
        RECT 1228.020 -37.520 1231.020 54.000 ;
        RECT 1408.020 -37.520 1411.020 54.000 ;
        RECT 1588.020 -37.520 1591.020 54.000 ;
        RECT 1768.020 -37.520 1771.020 54.000 ;
        RECT 1948.020 -37.520 1951.020 54.000 ;
        RECT 2128.020 -37.520 2131.020 54.000 ;
        RECT 2308.020 -37.520 2311.020 54.000 ;
        RECT 2488.020 -37.520 2491.020 54.000 ;
        RECT 2668.020 -37.520 2671.020 54.000 ;
        RECT 2848.020 -37.520 2851.020 54.000 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 54.000 3396.380 ;
        RECT 2866.000 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 54.000 3216.380 ;
        RECT 2866.000 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 54.000 3036.380 ;
        RECT 2866.000 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 54.000 2856.380 ;
        RECT 2866.000 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 54.000 2676.380 ;
        RECT 2866.000 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 54.000 2496.380 ;
        RECT 2866.000 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 54.000 2316.380 ;
        RECT 2866.000 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 54.000 2136.380 ;
        RECT 2866.000 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 54.000 1956.380 ;
        RECT 2866.000 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 54.000 1776.380 ;
        RECT 2866.000 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 54.000 1596.380 ;
        RECT 2866.000 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 54.000 1416.380 ;
        RECT 2866.000 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 54.000 1236.380 ;
        RECT 2866.000 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 54.000 1056.380 ;
        RECT 2866.000 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 54.000 876.380 ;
        RECT 2866.000 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 54.000 696.380 ;
        RECT 2866.000 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 54.000 516.380 ;
        RECT 2866.000 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 54.000 336.380 ;
        RECT 2866.000 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 54.000 156.380 ;
        RECT 2866.000 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 203.155 330.795 2691.755 3407.285 ;
      LAYER met1 ;
        RECT 54.000 89.800 2866.000 3464.220 ;
      LAYER met2 ;
        RECT 54.840 54.000 2839.480 3466.000 ;
      LAYER met3 ;
        RECT 54.000 138.215 2866.000 3435.865 ;
      LAYER met4 ;
        RECT 58.020 54.000 2851.020 3466.000 ;
      LAYER met5 ;
        RECT 54.000 63.370 2866.000 3466.000 ;
  END
END user_project_wrapper
END LIBRARY

