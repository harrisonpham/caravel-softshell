VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN -0.005 0.000 ;
  SIZE 2494.885 BY 3100.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.310 3096.000 8.590 3100.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 666.110 3096.000 666.390 3100.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 731.890 3096.000 732.170 3100.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 797.670 3096.000 797.950 3100.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 863.450 3096.000 863.730 3100.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.230 3096.000 929.510 3100.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 995.010 3096.000 995.290 3100.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1060.790 3096.000 1061.070 3100.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.570 3096.000 1126.850 3100.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1192.350 3096.000 1192.630 3100.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1258.130 3096.000 1258.410 3100.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.090 3096.000 74.370 3100.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1323.910 3096.000 1324.190 3100.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1389.690 3096.000 1389.970 3100.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1455.470 3096.000 1455.750 3100.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1521.250 3096.000 1521.530 3100.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1587.030 3096.000 1587.310 3100.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1652.810 3096.000 1653.090 3100.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1718.590 3096.000 1718.870 3100.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1784.370 3096.000 1784.650 3100.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1850.150 3096.000 1850.430 3100.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1915.930 3096.000 1916.210 3100.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.870 3096.000 140.150 3100.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1981.710 3096.000 1981.990 3100.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2047.490 3096.000 2047.770 3100.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.270 3096.000 2113.550 3100.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2179.050 3096.000 2179.330 3100.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2244.830 3096.000 2245.110 3100.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.610 3096.000 2310.890 3100.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2376.390 3096.000 2376.670 3100.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2442.170 3096.000 2442.450 3100.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 205.650 3096.000 205.930 3100.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 271.430 3096.000 271.710 3100.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 337.210 3096.000 337.490 3100.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 402.990 3096.000 403.270 3100.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 468.770 3096.000 469.050 3100.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 534.550 3096.000 534.830 3100.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 600.330 3096.000 600.610 3100.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.930 3096.000 30.210 3100.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 687.730 3096.000 688.010 3100.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 753.510 3096.000 753.790 3100.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 819.290 3096.000 819.570 3100.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 885.530 3096.000 885.810 3100.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 951.310 3096.000 951.590 3100.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1017.090 3096.000 1017.370 3100.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1082.870 3096.000 1083.150 3100.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1148.650 3096.000 1148.930 3100.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1214.430 3096.000 1214.710 3100.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1280.210 3096.000 1280.490 3100.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.710 3096.000 95.990 3100.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1345.990 3096.000 1346.270 3100.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1411.770 3096.000 1412.050 3100.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.550 3096.000 1477.830 3100.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1543.330 3096.000 1543.610 3100.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1609.110 3096.000 1609.390 3100.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1674.890 3096.000 1675.170 3100.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1740.670 3096.000 1740.950 3100.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1806.450 3096.000 1806.730 3100.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1872.230 3096.000 1872.510 3100.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1938.010 3096.000 1938.290 3100.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 161.490 3096.000 161.770 3100.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2003.790 3096.000 2004.070 3100.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2069.570 3096.000 2069.850 3100.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2135.350 3096.000 2135.630 3100.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2201.130 3096.000 2201.410 3100.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2266.910 3096.000 2267.190 3100.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2332.690 3096.000 2332.970 3100.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2398.470 3096.000 2398.750 3100.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2464.250 3096.000 2464.530 3100.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 227.270 3096.000 227.550 3100.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 293.050 3096.000 293.330 3100.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 358.830 3096.000 359.110 3100.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 424.610 3096.000 424.890 3100.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 490.390 3096.000 490.670 3100.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 556.170 3096.000 556.450 3100.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 621.950 3096.000 622.230 3100.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.010 3096.000 52.290 3100.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 709.810 3096.000 710.090 3100.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 775.590 3096.000 775.870 3100.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 841.370 3096.000 841.650 3100.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 907.150 3096.000 907.430 3100.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 972.930 3096.000 973.210 3100.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1038.710 3096.000 1038.990 3100.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1104.490 3096.000 1104.770 3100.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1170.270 3096.000 1170.550 3100.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1236.050 3096.000 1236.330 3100.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1301.830 3096.000 1302.110 3100.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.790 3096.000 118.070 3100.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1367.610 3096.000 1367.890 3100.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1433.390 3096.000 1433.670 3100.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1499.170 3096.000 1499.450 3100.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1564.950 3096.000 1565.230 3100.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1630.730 3096.000 1631.010 3100.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1696.970 3096.000 1697.250 3100.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.750 3096.000 1763.030 3100.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1828.530 3096.000 1828.810 3100.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1894.310 3096.000 1894.590 3100.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1960.090 3096.000 1960.370 3100.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.570 3096.000 183.850 3100.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2025.870 3096.000 2026.150 3100.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2091.650 3096.000 2091.930 3100.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2157.430 3096.000 2157.710 3100.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2223.210 3096.000 2223.490 3100.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2288.990 3096.000 2289.270 3100.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2354.770 3096.000 2355.050 3100.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2420.550 3096.000 2420.830 3100.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2486.330 3096.000 2486.610 3100.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 249.350 3096.000 249.630 3100.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 315.130 3096.000 315.410 3100.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 380.910 3096.000 381.190 3100.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 446.690 3096.000 446.970 3100.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 512.470 3096.000 512.750 3100.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 578.250 3096.000 578.530 3100.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 644.030 3096.000 644.310 3100.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 540.530 0.000 540.810 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2071.410 0.000 2071.690 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2086.590 0.000 2086.870 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2101.770 0.000 2102.050 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2117.410 0.000 2117.690 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2132.590 0.000 2132.870 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2147.770 0.000 2148.050 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2162.950 0.000 2163.230 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.590 0.000 2178.870 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2193.770 0.000 2194.050 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2208.950 0.000 2209.230 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 693.710 0.000 693.990 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2224.590 0.000 2224.870 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2239.770 0.000 2240.050 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2254.950 0.000 2255.230 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2270.130 0.000 2270.410 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2285.770 0.000 2286.050 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2300.950 0.000 2301.230 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2316.130 0.000 2316.410 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2331.310 0.000 2331.590 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2346.950 0.000 2347.230 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2362.130 0.000 2362.410 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 708.890 0.000 709.170 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2377.310 0.000 2377.590 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2392.950 0.000 2393.230 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2408.130 0.000 2408.410 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2423.310 0.000 2423.590 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2438.490 0.000 2438.770 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2454.130 0.000 2454.410 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2469.310 0.000 2469.590 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2484.490 0.000 2484.770 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 724.530 0.000 724.810 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 739.710 0.000 739.990 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 754.890 0.000 755.170 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 770.070 0.000 770.350 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 785.710 0.000 785.990 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 800.890 0.000 801.170 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 816.070 0.000 816.350 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 831.250 0.000 831.530 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 556.170 0.000 556.450 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.890 0.000 847.170 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 862.070 0.000 862.350 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 877.250 0.000 877.530 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 892.890 0.000 893.170 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 908.070 0.000 908.350 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 923.250 0.000 923.530 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 938.430 0.000 938.710 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 954.070 0.000 954.350 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 969.250 0.000 969.530 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 984.430 0.000 984.710 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 571.350 0.000 571.630 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1000.070 0.000 1000.350 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1015.250 0.000 1015.530 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1030.430 0.000 1030.710 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1045.610 0.000 1045.890 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.250 0.000 1061.530 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1076.430 0.000 1076.710 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1091.610 0.000 1091.890 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1106.790 0.000 1107.070 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1122.430 0.000 1122.710 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1137.610 0.000 1137.890 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 586.530 0.000 586.810 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1152.790 0.000 1153.070 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.430 0.000 1168.710 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1183.610 0.000 1183.890 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1198.790 0.000 1199.070 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1213.970 0.000 1214.250 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1229.610 0.000 1229.890 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1244.790 0.000 1245.070 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1259.970 0.000 1260.250 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.150 0.000 1275.430 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1290.790 0.000 1291.070 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 601.710 0.000 601.990 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1305.970 0.000 1306.250 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1321.150 0.000 1321.430 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1336.790 0.000 1337.070 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1351.970 0.000 1352.250 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1367.150 0.000 1367.430 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.330 0.000 1382.610 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1397.970 0.000 1398.250 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1413.150 0.000 1413.430 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1428.330 0.000 1428.610 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1443.510 0.000 1443.790 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 617.350 0.000 617.630 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1459.150 0.000 1459.430 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1474.330 0.000 1474.610 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.510 0.000 1489.790 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1505.150 0.000 1505.430 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1520.330 0.000 1520.610 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1535.510 0.000 1535.790 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1550.690 0.000 1550.970 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1566.330 0.000 1566.610 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1581.510 0.000 1581.790 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.690 0.000 1596.970 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 632.530 0.000 632.810 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1612.330 0.000 1612.610 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1627.510 0.000 1627.790 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1642.690 0.000 1642.970 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1657.870 0.000 1658.150 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1673.510 0.000 1673.790 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1688.690 0.000 1688.970 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.870 0.000 1704.150 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1719.050 0.000 1719.330 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1734.690 0.000 1734.970 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1749.870 0.000 1750.150 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 647.710 0.000 647.990 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1765.050 0.000 1765.330 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1780.690 0.000 1780.970 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1795.870 0.000 1796.150 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1811.050 0.000 1811.330 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1826.230 0.000 1826.510 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1841.870 0.000 1842.150 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.050 0.000 1857.330 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1872.230 0.000 1872.510 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1887.410 0.000 1887.690 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1903.050 0.000 1903.330 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.890 0.000 663.170 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1918.230 0.000 1918.510 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1933.410 0.000 1933.690 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1949.050 0.000 1949.330 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1964.230 0.000 1964.510 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1979.410 0.000 1979.690 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1994.590 0.000 1994.870 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2010.230 0.000 2010.510 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2025.410 0.000 2025.690 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2040.590 0.000 2040.870 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2056.230 0.000 2056.510 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 678.530 0.000 678.810 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 545.590 0.000 545.870 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2076.470 0.000 2076.750 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2091.650 0.000 2091.930 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2106.830 0.000 2107.110 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2122.470 0.000 2122.750 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.650 0.000 2137.930 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2152.830 0.000 2153.110 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2168.470 0.000 2168.750 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2183.650 0.000 2183.930 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2198.830 0.000 2199.110 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2214.010 0.000 2214.290 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 698.770 0.000 699.050 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2229.650 0.000 2229.930 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.830 0.000 2245.110 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2260.010 0.000 2260.290 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2275.190 0.000 2275.470 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2290.830 0.000 2291.110 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2306.010 0.000 2306.290 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2321.190 0.000 2321.470 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2336.830 0.000 2337.110 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2352.010 0.000 2352.290 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2367.190 0.000 2367.470 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 713.950 0.000 714.230 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2382.370 0.000 2382.650 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2398.010 0.000 2398.290 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2413.190 0.000 2413.470 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2428.370 0.000 2428.650 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2443.550 0.000 2443.830 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2459.190 0.000 2459.470 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2474.370 0.000 2474.650 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2489.550 0.000 2489.830 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 729.590 0.000 729.870 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 744.770 0.000 745.050 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 759.950 0.000 760.230 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 775.130 0.000 775.410 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 790.770 0.000 791.050 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 805.950 0.000 806.230 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 821.130 0.000 821.410 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 836.770 0.000 837.050 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 561.230 0.000 561.510 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 851.950 0.000 852.230 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 867.130 0.000 867.410 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 882.310 0.000 882.590 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 897.950 0.000 898.230 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 913.130 0.000 913.410 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 928.310 0.000 928.590 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 943.490 0.000 943.770 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.130 0.000 959.410 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 974.310 0.000 974.590 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 989.490 0.000 989.770 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 576.410 0.000 576.690 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1005.130 0.000 1005.410 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1020.310 0.000 1020.590 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1035.490 0.000 1035.770 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1050.670 0.000 1050.950 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1066.310 0.000 1066.590 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1081.490 0.000 1081.770 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1096.670 0.000 1096.950 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1112.310 0.000 1112.590 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1127.490 0.000 1127.770 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1142.670 0.000 1142.950 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 591.590 0.000 591.870 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1157.850 0.000 1158.130 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.490 0.000 1173.770 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1188.670 0.000 1188.950 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1203.850 0.000 1204.130 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1219.030 0.000 1219.310 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1234.670 0.000 1234.950 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1249.850 0.000 1250.130 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1265.030 0.000 1265.310 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1280.670 0.000 1280.950 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1295.850 0.000 1296.130 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 606.770 0.000 607.050 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1311.030 0.000 1311.310 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1326.210 0.000 1326.490 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1341.850 0.000 1342.130 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1357.030 0.000 1357.310 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1372.210 0.000 1372.490 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1387.390 0.000 1387.670 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1403.030 0.000 1403.310 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1418.210 0.000 1418.490 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1433.390 0.000 1433.670 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1449.030 0.000 1449.310 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 622.410 0.000 622.690 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1464.210 0.000 1464.490 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1479.390 0.000 1479.670 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1494.570 0.000 1494.850 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1510.210 0.000 1510.490 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1525.390 0.000 1525.670 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1540.570 0.000 1540.850 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1556.210 0.000 1556.490 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1571.390 0.000 1571.670 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1586.570 0.000 1586.850 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1601.750 0.000 1602.030 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 637.590 0.000 637.870 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1617.390 0.000 1617.670 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1632.570 0.000 1632.850 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1647.750 0.000 1648.030 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.930 0.000 1663.210 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1678.570 0.000 1678.850 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1693.750 0.000 1694.030 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1708.930 0.000 1709.210 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1724.570 0.000 1724.850 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1739.750 0.000 1740.030 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1754.930 0.000 1755.210 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 652.770 0.000 653.050 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1770.110 0.000 1770.390 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1785.750 0.000 1786.030 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1800.930 0.000 1801.210 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.110 0.000 1816.390 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1831.290 0.000 1831.570 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1846.930 0.000 1847.210 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1862.110 0.000 1862.390 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1877.290 0.000 1877.570 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1892.930 0.000 1893.210 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1908.110 0.000 1908.390 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 668.410 0.000 668.690 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.290 0.000 1923.570 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1938.470 0.000 1938.750 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1954.110 0.000 1954.390 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1969.290 0.000 1969.570 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1984.470 0.000 1984.750 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2000.110 0.000 2000.390 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2015.290 0.000 2015.570 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.470 0.000 2030.750 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2045.650 0.000 2045.930 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2061.290 0.000 2061.570 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 683.590 0.000 683.870 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 550.650 0.000 550.930 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2081.530 0.000 2081.810 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2096.710 0.000 2096.990 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2112.350 0.000 2112.630 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2127.530 0.000 2127.810 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2142.710 0.000 2142.990 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2157.890 0.000 2158.170 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2173.530 0.000 2173.810 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2188.710 0.000 2188.990 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2203.890 0.000 2204.170 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2219.070 0.000 2219.350 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 703.830 0.000 704.110 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2234.710 0.000 2234.990 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2249.890 0.000 2250.170 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2265.070 0.000 2265.350 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2280.710 0.000 2280.990 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2295.890 0.000 2296.170 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2311.070 0.000 2311.350 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2326.250 0.000 2326.530 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2341.890 0.000 2342.170 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.070 0.000 2357.350 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2372.250 0.000 2372.530 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 719.010 0.000 719.290 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2387.430 0.000 2387.710 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2403.070 0.000 2403.350 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2418.250 0.000 2418.530 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2433.430 0.000 2433.710 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2449.070 0.000 2449.350 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.250 0.000 2464.530 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2479.430 0.000 2479.710 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2494.610 0.000 2494.890 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.650 0.000 734.930 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 749.830 0.000 750.110 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 765.010 0.000 765.290 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 780.650 0.000 780.930 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 795.830 0.000 796.110 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.010 0.000 811.290 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 826.190 0.000 826.470 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 841.830 0.000 842.110 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 566.290 0.000 566.570 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 857.010 0.000 857.290 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 872.190 0.000 872.470 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 887.370 0.000 887.650 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 903.010 0.000 903.290 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.190 0.000 918.470 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 933.370 0.000 933.650 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.010 0.000 949.290 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 964.190 0.000 964.470 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 979.370 0.000 979.650 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 994.550 0.000 994.830 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 581.470 0.000 581.750 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1010.190 0.000 1010.470 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.370 0.000 1025.650 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1040.550 0.000 1040.830 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1056.190 0.000 1056.470 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1071.370 0.000 1071.650 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1086.550 0.000 1086.830 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1101.730 0.000 1102.010 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1117.370 0.000 1117.650 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.550 0.000 1132.830 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1147.730 0.000 1148.010 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 596.650 0.000 596.930 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.910 0.000 1163.190 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1178.550 0.000 1178.830 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1193.730 0.000 1194.010 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1208.910 0.000 1209.190 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1224.550 0.000 1224.830 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.730 0.000 1240.010 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1254.910 0.000 1255.190 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1270.090 0.000 1270.370 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1285.730 0.000 1286.010 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1300.910 0.000 1301.190 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 612.290 0.000 612.570 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1316.090 0.000 1316.370 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1331.270 0.000 1331.550 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.910 0.000 1347.190 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1362.090 0.000 1362.370 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1377.270 0.000 1377.550 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1392.910 0.000 1393.190 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1408.090 0.000 1408.370 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1423.270 0.000 1423.550 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1438.450 0.000 1438.730 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1454.090 0.000 1454.370 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 627.470 0.000 627.750 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1469.270 0.000 1469.550 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1484.450 0.000 1484.730 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1500.090 0.000 1500.370 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1515.270 0.000 1515.550 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1530.450 0.000 1530.730 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1545.630 0.000 1545.910 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1561.270 0.000 1561.550 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1576.450 0.000 1576.730 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1591.630 0.000 1591.910 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1606.810 0.000 1607.090 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 642.650 0.000 642.930 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1622.450 0.000 1622.730 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1637.630 0.000 1637.910 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1652.810 0.000 1653.090 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1668.450 0.000 1668.730 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1683.630 0.000 1683.910 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1698.810 0.000 1699.090 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1713.990 0.000 1714.270 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1729.630 0.000 1729.910 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1744.810 0.000 1745.090 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1759.990 0.000 1760.270 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 657.830 0.000 658.110 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1775.170 0.000 1775.450 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1790.810 0.000 1791.090 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1805.990 0.000 1806.270 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1821.170 0.000 1821.450 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1836.810 0.000 1837.090 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1851.990 0.000 1852.270 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1867.170 0.000 1867.450 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1882.350 0.000 1882.630 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1897.990 0.000 1898.270 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1913.170 0.000 1913.450 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 673.470 0.000 673.750 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1928.350 0.000 1928.630 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1943.530 0.000 1943.810 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1959.170 0.000 1959.450 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1974.350 0.000 1974.630 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1989.530 0.000 1989.810 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2005.170 0.000 2005.450 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2020.350 0.000 2020.630 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2035.530 0.000 2035.810 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2050.710 0.000 2050.990 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2066.350 0.000 2066.630 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 688.650 0.000 688.930 4.000 ;
    END
  END la_oen[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.030 0.000 0.310 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.090 0.000 5.370 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.150 0.000 10.430 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.390 0.000 30.670 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 203.810 0.000 204.090 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.990 0.000 219.270 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 234.630 0.000 234.910 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 249.810 0.000 250.090 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.990 0.000 265.270 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 280.630 0.000 280.910 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 295.810 0.000 296.090 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 310.990 0.000 311.270 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 326.170 0.000 326.450 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 341.810 0.000 342.090 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.630 0.000 50.910 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 356.990 0.000 357.270 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 372.170 0.000 372.450 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 387.350 0.000 387.630 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 402.990 0.000 403.270 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 418.170 0.000 418.450 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 433.350 0.000 433.630 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 448.990 0.000 449.270 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 464.170 0.000 464.450 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 479.350 0.000 479.630 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 494.530 0.000 494.810 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.330 0.000 71.610 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 510.170 0.000 510.450 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.350 0.000 525.630 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.570 0.000 91.850 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.270 0.000 112.550 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.450 0.000 127.730 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 142.630 0.000 142.910 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.810 0.000 158.090 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.450 0.000 173.730 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 188.630 0.000 188.910 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.210 0.000 15.490 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.450 0.000 35.730 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.870 0.000 209.150 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.510 0.000 224.790 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 239.690 0.000 239.970 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.870 0.000 255.150 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 270.050 0.000 270.330 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 285.690 0.000 285.970 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.870 0.000 301.150 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.050 0.000 316.330 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 331.230 0.000 331.510 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 346.870 0.000 347.150 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.150 0.000 56.430 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 362.050 0.000 362.330 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 377.230 0.000 377.510 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 392.870 0.000 393.150 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 408.050 0.000 408.330 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 423.230 0.000 423.510 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 438.410 0.000 438.690 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.050 0.000 454.330 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 469.230 0.000 469.510 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 484.410 0.000 484.690 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 500.050 0.000 500.330 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.390 0.000 76.670 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 515.230 0.000 515.510 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 530.410 0.000 530.690 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.630 0.000 96.910 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.330 0.000 117.610 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.510 0.000 132.790 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 147.690 0.000 147.970 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 162.870 0.000 163.150 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.510 0.000 178.790 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 193.690 0.000 193.970 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.510 0.000 40.790 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 213.930 0.000 214.210 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 229.570 0.000 229.850 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 244.750 0.000 245.030 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 259.930 0.000 260.210 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 275.110 0.000 275.390 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 290.750 0.000 291.030 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.930 0.000 306.210 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 321.110 0.000 321.390 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 336.750 0.000 337.030 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 351.930 0.000 352.210 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.210 0.000 61.490 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 367.110 0.000 367.390 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 382.290 0.000 382.570 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 397.930 0.000 398.210 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.110 0.000 413.390 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 428.290 0.000 428.570 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 443.470 0.000 443.750 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 459.110 0.000 459.390 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 474.290 0.000 474.570 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 489.470 0.000 489.750 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 505.110 0.000 505.390 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.450 0.000 81.730 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 520.290 0.000 520.570 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 535.470 0.000 535.750 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.690 0.000 101.970 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 122.390 0.000 122.670 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.570 0.000 137.850 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 152.750 0.000 153.030 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 168.390 0.000 168.670 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.570 0.000 183.850 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.750 0.000 199.030 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.570 0.000 45.850 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.270 0.000 66.550 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.510 0.000 86.790 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 106.750 0.000 107.030 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.270 0.000 20.550 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.330 0.000 25.610 4.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.680 10.640 20.280 3087.440 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.480 10.640 97.080 3087.440 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 3.160 10.795 2491.760 3087.285 ;
      LAYER met1 ;
        RECT 3.160 4.460 2491.760 3091.240 ;
      LAYER met2 ;
        RECT 0.030 3095.720 8.030 3096.000 ;
        RECT 8.870 3095.720 29.650 3096.000 ;
        RECT 30.490 3095.720 51.730 3096.000 ;
        RECT 52.570 3095.720 73.810 3096.000 ;
        RECT 74.650 3095.720 95.430 3096.000 ;
        RECT 96.270 3095.720 117.510 3096.000 ;
        RECT 118.350 3095.720 139.590 3096.000 ;
        RECT 140.430 3095.720 161.210 3096.000 ;
        RECT 162.050 3095.720 183.290 3096.000 ;
        RECT 184.130 3095.720 205.370 3096.000 ;
        RECT 206.210 3095.720 226.990 3096.000 ;
        RECT 227.830 3095.720 249.070 3096.000 ;
        RECT 249.910 3095.720 271.150 3096.000 ;
        RECT 271.990 3095.720 292.770 3096.000 ;
        RECT 293.610 3095.720 314.850 3096.000 ;
        RECT 315.690 3095.720 336.930 3096.000 ;
        RECT 337.770 3095.720 358.550 3096.000 ;
        RECT 359.390 3095.720 380.630 3096.000 ;
        RECT 381.470 3095.720 402.710 3096.000 ;
        RECT 403.550 3095.720 424.330 3096.000 ;
        RECT 425.170 3095.720 446.410 3096.000 ;
        RECT 447.250 3095.720 468.490 3096.000 ;
        RECT 469.330 3095.720 490.110 3096.000 ;
        RECT 490.950 3095.720 512.190 3096.000 ;
        RECT 513.030 3095.720 534.270 3096.000 ;
        RECT 535.110 3095.720 555.890 3096.000 ;
        RECT 556.730 3095.720 577.970 3096.000 ;
        RECT 578.810 3095.720 600.050 3096.000 ;
        RECT 600.890 3095.720 621.670 3096.000 ;
        RECT 622.510 3095.720 643.750 3096.000 ;
        RECT 644.590 3095.720 665.830 3096.000 ;
        RECT 666.670 3095.720 687.450 3096.000 ;
        RECT 688.290 3095.720 709.530 3096.000 ;
        RECT 710.370 3095.720 731.610 3096.000 ;
        RECT 732.450 3095.720 753.230 3096.000 ;
        RECT 754.070 3095.720 775.310 3096.000 ;
        RECT 776.150 3095.720 797.390 3096.000 ;
        RECT 798.230 3095.720 819.010 3096.000 ;
        RECT 819.850 3095.720 841.090 3096.000 ;
        RECT 841.930 3095.720 863.170 3096.000 ;
        RECT 864.010 3095.720 885.250 3096.000 ;
        RECT 886.090 3095.720 906.870 3096.000 ;
        RECT 907.710 3095.720 928.950 3096.000 ;
        RECT 929.790 3095.720 951.030 3096.000 ;
        RECT 951.870 3095.720 972.650 3096.000 ;
        RECT 973.490 3095.720 994.730 3096.000 ;
        RECT 995.570 3095.720 1016.810 3096.000 ;
        RECT 1017.650 3095.720 1038.430 3096.000 ;
        RECT 1039.270 3095.720 1060.510 3096.000 ;
        RECT 1061.350 3095.720 1082.590 3096.000 ;
        RECT 1083.430 3095.720 1104.210 3096.000 ;
        RECT 1105.050 3095.720 1126.290 3096.000 ;
        RECT 1127.130 3095.720 1148.370 3096.000 ;
        RECT 1149.210 3095.720 1169.990 3096.000 ;
        RECT 1170.830 3095.720 1192.070 3096.000 ;
        RECT 1192.910 3095.720 1214.150 3096.000 ;
        RECT 1214.990 3095.720 1235.770 3096.000 ;
        RECT 1236.610 3095.720 1257.850 3096.000 ;
        RECT 1258.690 3095.720 1279.930 3096.000 ;
        RECT 1280.770 3095.720 1301.550 3096.000 ;
        RECT 1302.390 3095.720 1323.630 3096.000 ;
        RECT 1324.470 3095.720 1345.710 3096.000 ;
        RECT 1346.550 3095.720 1367.330 3096.000 ;
        RECT 1368.170 3095.720 1389.410 3096.000 ;
        RECT 1390.250 3095.720 1411.490 3096.000 ;
        RECT 1412.330 3095.720 1433.110 3096.000 ;
        RECT 1433.950 3095.720 1455.190 3096.000 ;
        RECT 1456.030 3095.720 1477.270 3096.000 ;
        RECT 1478.110 3095.720 1498.890 3096.000 ;
        RECT 1499.730 3095.720 1520.970 3096.000 ;
        RECT 1521.810 3095.720 1543.050 3096.000 ;
        RECT 1543.890 3095.720 1564.670 3096.000 ;
        RECT 1565.510 3095.720 1586.750 3096.000 ;
        RECT 1587.590 3095.720 1608.830 3096.000 ;
        RECT 1609.670 3095.720 1630.450 3096.000 ;
        RECT 1631.290 3095.720 1652.530 3096.000 ;
        RECT 1653.370 3095.720 1674.610 3096.000 ;
        RECT 1675.450 3095.720 1696.690 3096.000 ;
        RECT 1697.530 3095.720 1718.310 3096.000 ;
        RECT 1719.150 3095.720 1740.390 3096.000 ;
        RECT 1741.230 3095.720 1762.470 3096.000 ;
        RECT 1763.310 3095.720 1784.090 3096.000 ;
        RECT 1784.930 3095.720 1806.170 3096.000 ;
        RECT 1807.010 3095.720 1828.250 3096.000 ;
        RECT 1829.090 3095.720 1849.870 3096.000 ;
        RECT 1850.710 3095.720 1871.950 3096.000 ;
        RECT 1872.790 3095.720 1894.030 3096.000 ;
        RECT 1894.870 3095.720 1915.650 3096.000 ;
        RECT 1916.490 3095.720 1937.730 3096.000 ;
        RECT 1938.570 3095.720 1959.810 3096.000 ;
        RECT 1960.650 3095.720 1981.430 3096.000 ;
        RECT 1982.270 3095.720 2003.510 3096.000 ;
        RECT 2004.350 3095.720 2025.590 3096.000 ;
        RECT 2026.430 3095.720 2047.210 3096.000 ;
        RECT 2048.050 3095.720 2069.290 3096.000 ;
        RECT 2070.130 3095.720 2091.370 3096.000 ;
        RECT 2092.210 3095.720 2112.990 3096.000 ;
        RECT 2113.830 3095.720 2135.070 3096.000 ;
        RECT 2135.910 3095.720 2157.150 3096.000 ;
        RECT 2157.990 3095.720 2178.770 3096.000 ;
        RECT 2179.610 3095.720 2200.850 3096.000 ;
        RECT 2201.690 3095.720 2222.930 3096.000 ;
        RECT 2223.770 3095.720 2244.550 3096.000 ;
        RECT 2245.390 3095.720 2266.630 3096.000 ;
        RECT 2267.470 3095.720 2288.710 3096.000 ;
        RECT 2289.550 3095.720 2310.330 3096.000 ;
        RECT 2311.170 3095.720 2332.410 3096.000 ;
        RECT 2333.250 3095.720 2354.490 3096.000 ;
        RECT 2355.330 3095.720 2376.110 3096.000 ;
        RECT 2376.950 3095.720 2398.190 3096.000 ;
        RECT 2399.030 3095.720 2420.270 3096.000 ;
        RECT 2421.110 3095.720 2441.890 3096.000 ;
        RECT 2442.730 3095.720 2463.970 3096.000 ;
        RECT 2464.810 3095.720 2486.050 3096.000 ;
        RECT 2486.890 3095.720 2489.820 3096.000 ;
        RECT 0.030 4.280 2489.820 3095.720 ;
        RECT 0.590 4.000 4.810 4.280 ;
        RECT 5.650 4.000 9.870 4.280 ;
        RECT 10.710 4.000 14.930 4.280 ;
        RECT 15.770 4.000 19.990 4.280 ;
        RECT 20.830 4.000 25.050 4.280 ;
        RECT 25.890 4.000 30.110 4.280 ;
        RECT 30.950 4.000 35.170 4.280 ;
        RECT 36.010 4.000 40.230 4.280 ;
        RECT 41.070 4.000 45.290 4.280 ;
        RECT 46.130 4.000 50.350 4.280 ;
        RECT 51.190 4.000 55.870 4.280 ;
        RECT 56.710 4.000 60.930 4.280 ;
        RECT 61.770 4.000 65.990 4.280 ;
        RECT 66.830 4.000 71.050 4.280 ;
        RECT 71.890 4.000 76.110 4.280 ;
        RECT 76.950 4.000 81.170 4.280 ;
        RECT 82.010 4.000 86.230 4.280 ;
        RECT 87.070 4.000 91.290 4.280 ;
        RECT 92.130 4.000 96.350 4.280 ;
        RECT 97.190 4.000 101.410 4.280 ;
        RECT 102.250 4.000 106.470 4.280 ;
        RECT 107.310 4.000 111.990 4.280 ;
        RECT 112.830 4.000 117.050 4.280 ;
        RECT 117.890 4.000 122.110 4.280 ;
        RECT 122.950 4.000 127.170 4.280 ;
        RECT 128.010 4.000 132.230 4.280 ;
        RECT 133.070 4.000 137.290 4.280 ;
        RECT 138.130 4.000 142.350 4.280 ;
        RECT 143.190 4.000 147.410 4.280 ;
        RECT 148.250 4.000 152.470 4.280 ;
        RECT 153.310 4.000 157.530 4.280 ;
        RECT 158.370 4.000 162.590 4.280 ;
        RECT 163.430 4.000 168.110 4.280 ;
        RECT 168.950 4.000 173.170 4.280 ;
        RECT 174.010 4.000 178.230 4.280 ;
        RECT 179.070 4.000 183.290 4.280 ;
        RECT 184.130 4.000 188.350 4.280 ;
        RECT 189.190 4.000 193.410 4.280 ;
        RECT 194.250 4.000 198.470 4.280 ;
        RECT 199.310 4.000 203.530 4.280 ;
        RECT 204.370 4.000 208.590 4.280 ;
        RECT 209.430 4.000 213.650 4.280 ;
        RECT 214.490 4.000 218.710 4.280 ;
        RECT 219.550 4.000 224.230 4.280 ;
        RECT 225.070 4.000 229.290 4.280 ;
        RECT 230.130 4.000 234.350 4.280 ;
        RECT 235.190 4.000 239.410 4.280 ;
        RECT 240.250 4.000 244.470 4.280 ;
        RECT 245.310 4.000 249.530 4.280 ;
        RECT 250.370 4.000 254.590 4.280 ;
        RECT 255.430 4.000 259.650 4.280 ;
        RECT 260.490 4.000 264.710 4.280 ;
        RECT 265.550 4.000 269.770 4.280 ;
        RECT 270.610 4.000 274.830 4.280 ;
        RECT 275.670 4.000 280.350 4.280 ;
        RECT 281.190 4.000 285.410 4.280 ;
        RECT 286.250 4.000 290.470 4.280 ;
        RECT 291.310 4.000 295.530 4.280 ;
        RECT 296.370 4.000 300.590 4.280 ;
        RECT 301.430 4.000 305.650 4.280 ;
        RECT 306.490 4.000 310.710 4.280 ;
        RECT 311.550 4.000 315.770 4.280 ;
        RECT 316.610 4.000 320.830 4.280 ;
        RECT 321.670 4.000 325.890 4.280 ;
        RECT 326.730 4.000 330.950 4.280 ;
        RECT 331.790 4.000 336.470 4.280 ;
        RECT 337.310 4.000 341.530 4.280 ;
        RECT 342.370 4.000 346.590 4.280 ;
        RECT 347.430 4.000 351.650 4.280 ;
        RECT 352.490 4.000 356.710 4.280 ;
        RECT 357.550 4.000 361.770 4.280 ;
        RECT 362.610 4.000 366.830 4.280 ;
        RECT 367.670 4.000 371.890 4.280 ;
        RECT 372.730 4.000 376.950 4.280 ;
        RECT 377.790 4.000 382.010 4.280 ;
        RECT 382.850 4.000 387.070 4.280 ;
        RECT 387.910 4.000 392.590 4.280 ;
        RECT 393.430 4.000 397.650 4.280 ;
        RECT 398.490 4.000 402.710 4.280 ;
        RECT 403.550 4.000 407.770 4.280 ;
        RECT 408.610 4.000 412.830 4.280 ;
        RECT 413.670 4.000 417.890 4.280 ;
        RECT 418.730 4.000 422.950 4.280 ;
        RECT 423.790 4.000 428.010 4.280 ;
        RECT 428.850 4.000 433.070 4.280 ;
        RECT 433.910 4.000 438.130 4.280 ;
        RECT 438.970 4.000 443.190 4.280 ;
        RECT 444.030 4.000 448.710 4.280 ;
        RECT 449.550 4.000 453.770 4.280 ;
        RECT 454.610 4.000 458.830 4.280 ;
        RECT 459.670 4.000 463.890 4.280 ;
        RECT 464.730 4.000 468.950 4.280 ;
        RECT 469.790 4.000 474.010 4.280 ;
        RECT 474.850 4.000 479.070 4.280 ;
        RECT 479.910 4.000 484.130 4.280 ;
        RECT 484.970 4.000 489.190 4.280 ;
        RECT 490.030 4.000 494.250 4.280 ;
        RECT 495.090 4.000 499.770 4.280 ;
        RECT 500.610 4.000 504.830 4.280 ;
        RECT 505.670 4.000 509.890 4.280 ;
        RECT 510.730 4.000 514.950 4.280 ;
        RECT 515.790 4.000 520.010 4.280 ;
        RECT 520.850 4.000 525.070 4.280 ;
        RECT 525.910 4.000 530.130 4.280 ;
        RECT 530.970 4.000 535.190 4.280 ;
        RECT 536.030 4.000 540.250 4.280 ;
        RECT 541.090 4.000 545.310 4.280 ;
        RECT 546.150 4.000 550.370 4.280 ;
        RECT 551.210 4.000 555.890 4.280 ;
        RECT 556.730 4.000 560.950 4.280 ;
        RECT 561.790 4.000 566.010 4.280 ;
        RECT 566.850 4.000 571.070 4.280 ;
        RECT 571.910 4.000 576.130 4.280 ;
        RECT 576.970 4.000 581.190 4.280 ;
        RECT 582.030 4.000 586.250 4.280 ;
        RECT 587.090 4.000 591.310 4.280 ;
        RECT 592.150 4.000 596.370 4.280 ;
        RECT 597.210 4.000 601.430 4.280 ;
        RECT 602.270 4.000 606.490 4.280 ;
        RECT 607.330 4.000 612.010 4.280 ;
        RECT 612.850 4.000 617.070 4.280 ;
        RECT 617.910 4.000 622.130 4.280 ;
        RECT 622.970 4.000 627.190 4.280 ;
        RECT 628.030 4.000 632.250 4.280 ;
        RECT 633.090 4.000 637.310 4.280 ;
        RECT 638.150 4.000 642.370 4.280 ;
        RECT 643.210 4.000 647.430 4.280 ;
        RECT 648.270 4.000 652.490 4.280 ;
        RECT 653.330 4.000 657.550 4.280 ;
        RECT 658.390 4.000 662.610 4.280 ;
        RECT 663.450 4.000 668.130 4.280 ;
        RECT 668.970 4.000 673.190 4.280 ;
        RECT 674.030 4.000 678.250 4.280 ;
        RECT 679.090 4.000 683.310 4.280 ;
        RECT 684.150 4.000 688.370 4.280 ;
        RECT 689.210 4.000 693.430 4.280 ;
        RECT 694.270 4.000 698.490 4.280 ;
        RECT 699.330 4.000 703.550 4.280 ;
        RECT 704.390 4.000 708.610 4.280 ;
        RECT 709.450 4.000 713.670 4.280 ;
        RECT 714.510 4.000 718.730 4.280 ;
        RECT 719.570 4.000 724.250 4.280 ;
        RECT 725.090 4.000 729.310 4.280 ;
        RECT 730.150 4.000 734.370 4.280 ;
        RECT 735.210 4.000 739.430 4.280 ;
        RECT 740.270 4.000 744.490 4.280 ;
        RECT 745.330 4.000 749.550 4.280 ;
        RECT 750.390 4.000 754.610 4.280 ;
        RECT 755.450 4.000 759.670 4.280 ;
        RECT 760.510 4.000 764.730 4.280 ;
        RECT 765.570 4.000 769.790 4.280 ;
        RECT 770.630 4.000 774.850 4.280 ;
        RECT 775.690 4.000 780.370 4.280 ;
        RECT 781.210 4.000 785.430 4.280 ;
        RECT 786.270 4.000 790.490 4.280 ;
        RECT 791.330 4.000 795.550 4.280 ;
        RECT 796.390 4.000 800.610 4.280 ;
        RECT 801.450 4.000 805.670 4.280 ;
        RECT 806.510 4.000 810.730 4.280 ;
        RECT 811.570 4.000 815.790 4.280 ;
        RECT 816.630 4.000 820.850 4.280 ;
        RECT 821.690 4.000 825.910 4.280 ;
        RECT 826.750 4.000 830.970 4.280 ;
        RECT 831.810 4.000 836.490 4.280 ;
        RECT 837.330 4.000 841.550 4.280 ;
        RECT 842.390 4.000 846.610 4.280 ;
        RECT 847.450 4.000 851.670 4.280 ;
        RECT 852.510 4.000 856.730 4.280 ;
        RECT 857.570 4.000 861.790 4.280 ;
        RECT 862.630 4.000 866.850 4.280 ;
        RECT 867.690 4.000 871.910 4.280 ;
        RECT 872.750 4.000 876.970 4.280 ;
        RECT 877.810 4.000 882.030 4.280 ;
        RECT 882.870 4.000 887.090 4.280 ;
        RECT 887.930 4.000 892.610 4.280 ;
        RECT 893.450 4.000 897.670 4.280 ;
        RECT 898.510 4.000 902.730 4.280 ;
        RECT 903.570 4.000 907.790 4.280 ;
        RECT 908.630 4.000 912.850 4.280 ;
        RECT 913.690 4.000 917.910 4.280 ;
        RECT 918.750 4.000 922.970 4.280 ;
        RECT 923.810 4.000 928.030 4.280 ;
        RECT 928.870 4.000 933.090 4.280 ;
        RECT 933.930 4.000 938.150 4.280 ;
        RECT 938.990 4.000 943.210 4.280 ;
        RECT 944.050 4.000 948.730 4.280 ;
        RECT 949.570 4.000 953.790 4.280 ;
        RECT 954.630 4.000 958.850 4.280 ;
        RECT 959.690 4.000 963.910 4.280 ;
        RECT 964.750 4.000 968.970 4.280 ;
        RECT 969.810 4.000 974.030 4.280 ;
        RECT 974.870 4.000 979.090 4.280 ;
        RECT 979.930 4.000 984.150 4.280 ;
        RECT 984.990 4.000 989.210 4.280 ;
        RECT 990.050 4.000 994.270 4.280 ;
        RECT 995.110 4.000 999.790 4.280 ;
        RECT 1000.630 4.000 1004.850 4.280 ;
        RECT 1005.690 4.000 1009.910 4.280 ;
        RECT 1010.750 4.000 1014.970 4.280 ;
        RECT 1015.810 4.000 1020.030 4.280 ;
        RECT 1020.870 4.000 1025.090 4.280 ;
        RECT 1025.930 4.000 1030.150 4.280 ;
        RECT 1030.990 4.000 1035.210 4.280 ;
        RECT 1036.050 4.000 1040.270 4.280 ;
        RECT 1041.110 4.000 1045.330 4.280 ;
        RECT 1046.170 4.000 1050.390 4.280 ;
        RECT 1051.230 4.000 1055.910 4.280 ;
        RECT 1056.750 4.000 1060.970 4.280 ;
        RECT 1061.810 4.000 1066.030 4.280 ;
        RECT 1066.870 4.000 1071.090 4.280 ;
        RECT 1071.930 4.000 1076.150 4.280 ;
        RECT 1076.990 4.000 1081.210 4.280 ;
        RECT 1082.050 4.000 1086.270 4.280 ;
        RECT 1087.110 4.000 1091.330 4.280 ;
        RECT 1092.170 4.000 1096.390 4.280 ;
        RECT 1097.230 4.000 1101.450 4.280 ;
        RECT 1102.290 4.000 1106.510 4.280 ;
        RECT 1107.350 4.000 1112.030 4.280 ;
        RECT 1112.870 4.000 1117.090 4.280 ;
        RECT 1117.930 4.000 1122.150 4.280 ;
        RECT 1122.990 4.000 1127.210 4.280 ;
        RECT 1128.050 4.000 1132.270 4.280 ;
        RECT 1133.110 4.000 1137.330 4.280 ;
        RECT 1138.170 4.000 1142.390 4.280 ;
        RECT 1143.230 4.000 1147.450 4.280 ;
        RECT 1148.290 4.000 1152.510 4.280 ;
        RECT 1153.350 4.000 1157.570 4.280 ;
        RECT 1158.410 4.000 1162.630 4.280 ;
        RECT 1163.470 4.000 1168.150 4.280 ;
        RECT 1168.990 4.000 1173.210 4.280 ;
        RECT 1174.050 4.000 1178.270 4.280 ;
        RECT 1179.110 4.000 1183.330 4.280 ;
        RECT 1184.170 4.000 1188.390 4.280 ;
        RECT 1189.230 4.000 1193.450 4.280 ;
        RECT 1194.290 4.000 1198.510 4.280 ;
        RECT 1199.350 4.000 1203.570 4.280 ;
        RECT 1204.410 4.000 1208.630 4.280 ;
        RECT 1209.470 4.000 1213.690 4.280 ;
        RECT 1214.530 4.000 1218.750 4.280 ;
        RECT 1219.590 4.000 1224.270 4.280 ;
        RECT 1225.110 4.000 1229.330 4.280 ;
        RECT 1230.170 4.000 1234.390 4.280 ;
        RECT 1235.230 4.000 1239.450 4.280 ;
        RECT 1240.290 4.000 1244.510 4.280 ;
        RECT 1245.350 4.000 1249.570 4.280 ;
        RECT 1250.410 4.000 1254.630 4.280 ;
        RECT 1255.470 4.000 1259.690 4.280 ;
        RECT 1260.530 4.000 1264.750 4.280 ;
        RECT 1265.590 4.000 1269.810 4.280 ;
        RECT 1270.650 4.000 1274.870 4.280 ;
        RECT 1275.710 4.000 1280.390 4.280 ;
        RECT 1281.230 4.000 1285.450 4.280 ;
        RECT 1286.290 4.000 1290.510 4.280 ;
        RECT 1291.350 4.000 1295.570 4.280 ;
        RECT 1296.410 4.000 1300.630 4.280 ;
        RECT 1301.470 4.000 1305.690 4.280 ;
        RECT 1306.530 4.000 1310.750 4.280 ;
        RECT 1311.590 4.000 1315.810 4.280 ;
        RECT 1316.650 4.000 1320.870 4.280 ;
        RECT 1321.710 4.000 1325.930 4.280 ;
        RECT 1326.770 4.000 1330.990 4.280 ;
        RECT 1331.830 4.000 1336.510 4.280 ;
        RECT 1337.350 4.000 1341.570 4.280 ;
        RECT 1342.410 4.000 1346.630 4.280 ;
        RECT 1347.470 4.000 1351.690 4.280 ;
        RECT 1352.530 4.000 1356.750 4.280 ;
        RECT 1357.590 4.000 1361.810 4.280 ;
        RECT 1362.650 4.000 1366.870 4.280 ;
        RECT 1367.710 4.000 1371.930 4.280 ;
        RECT 1372.770 4.000 1376.990 4.280 ;
        RECT 1377.830 4.000 1382.050 4.280 ;
        RECT 1382.890 4.000 1387.110 4.280 ;
        RECT 1387.950 4.000 1392.630 4.280 ;
        RECT 1393.470 4.000 1397.690 4.280 ;
        RECT 1398.530 4.000 1402.750 4.280 ;
        RECT 1403.590 4.000 1407.810 4.280 ;
        RECT 1408.650 4.000 1412.870 4.280 ;
        RECT 1413.710 4.000 1417.930 4.280 ;
        RECT 1418.770 4.000 1422.990 4.280 ;
        RECT 1423.830 4.000 1428.050 4.280 ;
        RECT 1428.890 4.000 1433.110 4.280 ;
        RECT 1433.950 4.000 1438.170 4.280 ;
        RECT 1439.010 4.000 1443.230 4.280 ;
        RECT 1444.070 4.000 1448.750 4.280 ;
        RECT 1449.590 4.000 1453.810 4.280 ;
        RECT 1454.650 4.000 1458.870 4.280 ;
        RECT 1459.710 4.000 1463.930 4.280 ;
        RECT 1464.770 4.000 1468.990 4.280 ;
        RECT 1469.830 4.000 1474.050 4.280 ;
        RECT 1474.890 4.000 1479.110 4.280 ;
        RECT 1479.950 4.000 1484.170 4.280 ;
        RECT 1485.010 4.000 1489.230 4.280 ;
        RECT 1490.070 4.000 1494.290 4.280 ;
        RECT 1495.130 4.000 1499.810 4.280 ;
        RECT 1500.650 4.000 1504.870 4.280 ;
        RECT 1505.710 4.000 1509.930 4.280 ;
        RECT 1510.770 4.000 1514.990 4.280 ;
        RECT 1515.830 4.000 1520.050 4.280 ;
        RECT 1520.890 4.000 1525.110 4.280 ;
        RECT 1525.950 4.000 1530.170 4.280 ;
        RECT 1531.010 4.000 1535.230 4.280 ;
        RECT 1536.070 4.000 1540.290 4.280 ;
        RECT 1541.130 4.000 1545.350 4.280 ;
        RECT 1546.190 4.000 1550.410 4.280 ;
        RECT 1551.250 4.000 1555.930 4.280 ;
        RECT 1556.770 4.000 1560.990 4.280 ;
        RECT 1561.830 4.000 1566.050 4.280 ;
        RECT 1566.890 4.000 1571.110 4.280 ;
        RECT 1571.950 4.000 1576.170 4.280 ;
        RECT 1577.010 4.000 1581.230 4.280 ;
        RECT 1582.070 4.000 1586.290 4.280 ;
        RECT 1587.130 4.000 1591.350 4.280 ;
        RECT 1592.190 4.000 1596.410 4.280 ;
        RECT 1597.250 4.000 1601.470 4.280 ;
        RECT 1602.310 4.000 1606.530 4.280 ;
        RECT 1607.370 4.000 1612.050 4.280 ;
        RECT 1612.890 4.000 1617.110 4.280 ;
        RECT 1617.950 4.000 1622.170 4.280 ;
        RECT 1623.010 4.000 1627.230 4.280 ;
        RECT 1628.070 4.000 1632.290 4.280 ;
        RECT 1633.130 4.000 1637.350 4.280 ;
        RECT 1638.190 4.000 1642.410 4.280 ;
        RECT 1643.250 4.000 1647.470 4.280 ;
        RECT 1648.310 4.000 1652.530 4.280 ;
        RECT 1653.370 4.000 1657.590 4.280 ;
        RECT 1658.430 4.000 1662.650 4.280 ;
        RECT 1663.490 4.000 1668.170 4.280 ;
        RECT 1669.010 4.000 1673.230 4.280 ;
        RECT 1674.070 4.000 1678.290 4.280 ;
        RECT 1679.130 4.000 1683.350 4.280 ;
        RECT 1684.190 4.000 1688.410 4.280 ;
        RECT 1689.250 4.000 1693.470 4.280 ;
        RECT 1694.310 4.000 1698.530 4.280 ;
        RECT 1699.370 4.000 1703.590 4.280 ;
        RECT 1704.430 4.000 1708.650 4.280 ;
        RECT 1709.490 4.000 1713.710 4.280 ;
        RECT 1714.550 4.000 1718.770 4.280 ;
        RECT 1719.610 4.000 1724.290 4.280 ;
        RECT 1725.130 4.000 1729.350 4.280 ;
        RECT 1730.190 4.000 1734.410 4.280 ;
        RECT 1735.250 4.000 1739.470 4.280 ;
        RECT 1740.310 4.000 1744.530 4.280 ;
        RECT 1745.370 4.000 1749.590 4.280 ;
        RECT 1750.430 4.000 1754.650 4.280 ;
        RECT 1755.490 4.000 1759.710 4.280 ;
        RECT 1760.550 4.000 1764.770 4.280 ;
        RECT 1765.610 4.000 1769.830 4.280 ;
        RECT 1770.670 4.000 1774.890 4.280 ;
        RECT 1775.730 4.000 1780.410 4.280 ;
        RECT 1781.250 4.000 1785.470 4.280 ;
        RECT 1786.310 4.000 1790.530 4.280 ;
        RECT 1791.370 4.000 1795.590 4.280 ;
        RECT 1796.430 4.000 1800.650 4.280 ;
        RECT 1801.490 4.000 1805.710 4.280 ;
        RECT 1806.550 4.000 1810.770 4.280 ;
        RECT 1811.610 4.000 1815.830 4.280 ;
        RECT 1816.670 4.000 1820.890 4.280 ;
        RECT 1821.730 4.000 1825.950 4.280 ;
        RECT 1826.790 4.000 1831.010 4.280 ;
        RECT 1831.850 4.000 1836.530 4.280 ;
        RECT 1837.370 4.000 1841.590 4.280 ;
        RECT 1842.430 4.000 1846.650 4.280 ;
        RECT 1847.490 4.000 1851.710 4.280 ;
        RECT 1852.550 4.000 1856.770 4.280 ;
        RECT 1857.610 4.000 1861.830 4.280 ;
        RECT 1862.670 4.000 1866.890 4.280 ;
        RECT 1867.730 4.000 1871.950 4.280 ;
        RECT 1872.790 4.000 1877.010 4.280 ;
        RECT 1877.850 4.000 1882.070 4.280 ;
        RECT 1882.910 4.000 1887.130 4.280 ;
        RECT 1887.970 4.000 1892.650 4.280 ;
        RECT 1893.490 4.000 1897.710 4.280 ;
        RECT 1898.550 4.000 1902.770 4.280 ;
        RECT 1903.610 4.000 1907.830 4.280 ;
        RECT 1908.670 4.000 1912.890 4.280 ;
        RECT 1913.730 4.000 1917.950 4.280 ;
        RECT 1918.790 4.000 1923.010 4.280 ;
        RECT 1923.850 4.000 1928.070 4.280 ;
        RECT 1928.910 4.000 1933.130 4.280 ;
        RECT 1933.970 4.000 1938.190 4.280 ;
        RECT 1939.030 4.000 1943.250 4.280 ;
        RECT 1944.090 4.000 1948.770 4.280 ;
        RECT 1949.610 4.000 1953.830 4.280 ;
        RECT 1954.670 4.000 1958.890 4.280 ;
        RECT 1959.730 4.000 1963.950 4.280 ;
        RECT 1964.790 4.000 1969.010 4.280 ;
        RECT 1969.850 4.000 1974.070 4.280 ;
        RECT 1974.910 4.000 1979.130 4.280 ;
        RECT 1979.970 4.000 1984.190 4.280 ;
        RECT 1985.030 4.000 1989.250 4.280 ;
        RECT 1990.090 4.000 1994.310 4.280 ;
        RECT 1995.150 4.000 1999.830 4.280 ;
        RECT 2000.670 4.000 2004.890 4.280 ;
        RECT 2005.730 4.000 2009.950 4.280 ;
        RECT 2010.790 4.000 2015.010 4.280 ;
        RECT 2015.850 4.000 2020.070 4.280 ;
        RECT 2020.910 4.000 2025.130 4.280 ;
        RECT 2025.970 4.000 2030.190 4.280 ;
        RECT 2031.030 4.000 2035.250 4.280 ;
        RECT 2036.090 4.000 2040.310 4.280 ;
        RECT 2041.150 4.000 2045.370 4.280 ;
        RECT 2046.210 4.000 2050.430 4.280 ;
        RECT 2051.270 4.000 2055.950 4.280 ;
        RECT 2056.790 4.000 2061.010 4.280 ;
        RECT 2061.850 4.000 2066.070 4.280 ;
        RECT 2066.910 4.000 2071.130 4.280 ;
        RECT 2071.970 4.000 2076.190 4.280 ;
        RECT 2077.030 4.000 2081.250 4.280 ;
        RECT 2082.090 4.000 2086.310 4.280 ;
        RECT 2087.150 4.000 2091.370 4.280 ;
        RECT 2092.210 4.000 2096.430 4.280 ;
        RECT 2097.270 4.000 2101.490 4.280 ;
        RECT 2102.330 4.000 2106.550 4.280 ;
        RECT 2107.390 4.000 2112.070 4.280 ;
        RECT 2112.910 4.000 2117.130 4.280 ;
        RECT 2117.970 4.000 2122.190 4.280 ;
        RECT 2123.030 4.000 2127.250 4.280 ;
        RECT 2128.090 4.000 2132.310 4.280 ;
        RECT 2133.150 4.000 2137.370 4.280 ;
        RECT 2138.210 4.000 2142.430 4.280 ;
        RECT 2143.270 4.000 2147.490 4.280 ;
        RECT 2148.330 4.000 2152.550 4.280 ;
        RECT 2153.390 4.000 2157.610 4.280 ;
        RECT 2158.450 4.000 2162.670 4.280 ;
        RECT 2163.510 4.000 2168.190 4.280 ;
        RECT 2169.030 4.000 2173.250 4.280 ;
        RECT 2174.090 4.000 2178.310 4.280 ;
        RECT 2179.150 4.000 2183.370 4.280 ;
        RECT 2184.210 4.000 2188.430 4.280 ;
        RECT 2189.270 4.000 2193.490 4.280 ;
        RECT 2194.330 4.000 2198.550 4.280 ;
        RECT 2199.390 4.000 2203.610 4.280 ;
        RECT 2204.450 4.000 2208.670 4.280 ;
        RECT 2209.510 4.000 2213.730 4.280 ;
        RECT 2214.570 4.000 2218.790 4.280 ;
        RECT 2219.630 4.000 2224.310 4.280 ;
        RECT 2225.150 4.000 2229.370 4.280 ;
        RECT 2230.210 4.000 2234.430 4.280 ;
        RECT 2235.270 4.000 2239.490 4.280 ;
        RECT 2240.330 4.000 2244.550 4.280 ;
        RECT 2245.390 4.000 2249.610 4.280 ;
        RECT 2250.450 4.000 2254.670 4.280 ;
        RECT 2255.510 4.000 2259.730 4.280 ;
        RECT 2260.570 4.000 2264.790 4.280 ;
        RECT 2265.630 4.000 2269.850 4.280 ;
        RECT 2270.690 4.000 2274.910 4.280 ;
        RECT 2275.750 4.000 2280.430 4.280 ;
        RECT 2281.270 4.000 2285.490 4.280 ;
        RECT 2286.330 4.000 2290.550 4.280 ;
        RECT 2291.390 4.000 2295.610 4.280 ;
        RECT 2296.450 4.000 2300.670 4.280 ;
        RECT 2301.510 4.000 2305.730 4.280 ;
        RECT 2306.570 4.000 2310.790 4.280 ;
        RECT 2311.630 4.000 2315.850 4.280 ;
        RECT 2316.690 4.000 2320.910 4.280 ;
        RECT 2321.750 4.000 2325.970 4.280 ;
        RECT 2326.810 4.000 2331.030 4.280 ;
        RECT 2331.870 4.000 2336.550 4.280 ;
        RECT 2337.390 4.000 2341.610 4.280 ;
        RECT 2342.450 4.000 2346.670 4.280 ;
        RECT 2347.510 4.000 2351.730 4.280 ;
        RECT 2352.570 4.000 2356.790 4.280 ;
        RECT 2357.630 4.000 2361.850 4.280 ;
        RECT 2362.690 4.000 2366.910 4.280 ;
        RECT 2367.750 4.000 2371.970 4.280 ;
        RECT 2372.810 4.000 2377.030 4.280 ;
        RECT 2377.870 4.000 2382.090 4.280 ;
        RECT 2382.930 4.000 2387.150 4.280 ;
        RECT 2387.990 4.000 2392.670 4.280 ;
        RECT 2393.510 4.000 2397.730 4.280 ;
        RECT 2398.570 4.000 2402.790 4.280 ;
        RECT 2403.630 4.000 2407.850 4.280 ;
        RECT 2408.690 4.000 2412.910 4.280 ;
        RECT 2413.750 4.000 2417.970 4.280 ;
        RECT 2418.810 4.000 2423.030 4.280 ;
        RECT 2423.870 4.000 2428.090 4.280 ;
        RECT 2428.930 4.000 2433.150 4.280 ;
        RECT 2433.990 4.000 2438.210 4.280 ;
        RECT 2439.050 4.000 2443.270 4.280 ;
        RECT 2444.110 4.000 2448.790 4.280 ;
        RECT 2449.630 4.000 2453.850 4.280 ;
        RECT 2454.690 4.000 2458.910 4.280 ;
        RECT 2459.750 4.000 2463.970 4.280 ;
        RECT 2464.810 4.000 2469.030 4.280 ;
        RECT 2469.870 4.000 2474.090 4.280 ;
        RECT 2474.930 4.000 2479.150 4.280 ;
        RECT 2479.990 4.000 2484.210 4.280 ;
        RECT 2485.050 4.000 2489.270 4.280 ;
      LAYER met3 ;
        RECT 0.005 4.255 2482.495 3087.365 ;
      LAYER met4 ;
        RECT 25.535 10.640 95.080 3087.440 ;
        RECT 97.480 10.640 2477.880 3087.440 ;
  END
END user_proj_example
END LIBRARY

