VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 229.150 3216.440 229.470 3216.700 ;
        RECT 229.240 3215.960 229.380 3216.440 ;
        RECT 2611.490 3215.960 2611.810 3216.020 ;
        RECT 229.240 3215.820 2611.810 3215.960 ;
        RECT 2611.490 3215.760 2611.810 3215.820 ;
        RECT 2611.490 89.660 2611.810 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2611.490 89.520 2899.310 89.660 ;
        RECT 2611.490 89.460 2611.810 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 229.180 3216.440 229.440 3216.700 ;
        RECT 2611.520 3215.760 2611.780 3216.020 ;
        RECT 2611.520 89.460 2611.780 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 227.840 3216.810 228.120 3220.000 ;
        RECT 227.840 3216.730 229.380 3216.810 ;
        RECT 227.840 3216.670 229.440 3216.730 ;
        RECT 227.840 3216.000 228.120 3216.670 ;
        RECT 229.180 3216.410 229.440 3216.670 ;
        RECT 2611.520 3215.730 2611.780 3216.050 ;
        RECT 2611.580 89.750 2611.720 3215.730 ;
        RECT 2611.520 89.430 2611.780 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 860.730 3218.680 861.050 3218.740 ;
        RECT 2839.190 3218.680 2839.510 3218.740 ;
        RECT 860.730 3218.540 2839.510 3218.680 ;
        RECT 860.730 3218.480 861.050 3218.540 ;
        RECT 2839.190 3218.480 2839.510 3218.540 ;
        RECT 2839.190 2435.660 2839.510 2435.720 ;
        RECT 2898.070 2435.660 2898.390 2435.720 ;
        RECT 2839.190 2435.520 2898.390 2435.660 ;
        RECT 2839.190 2435.460 2839.510 2435.520 ;
        RECT 2898.070 2435.460 2898.390 2435.520 ;
      LAYER via ;
        RECT 860.760 3218.480 861.020 3218.740 ;
        RECT 2839.220 3218.480 2839.480 3218.740 ;
        RECT 2839.220 2435.460 2839.480 2435.720 ;
        RECT 2898.100 2435.460 2898.360 2435.720 ;
      LAYER met2 ;
        RECT 858.960 3218.850 859.240 3220.000 ;
        RECT 858.960 3218.770 860.960 3218.850 ;
        RECT 858.960 3218.710 861.020 3218.770 ;
        RECT 858.960 3216.000 859.240 3218.710 ;
        RECT 860.760 3218.450 861.020 3218.710 ;
        RECT 2839.220 3218.450 2839.480 3218.770 ;
        RECT 2839.280 2435.750 2839.420 3218.450 ;
        RECT 2839.220 2435.430 2839.480 2435.750 ;
        RECT 2898.100 2435.430 2898.360 2435.750 ;
        RECT 2898.160 2434.245 2898.300 2435.430 ;
        RECT 2898.090 2433.875 2898.370 2434.245 ;
      LAYER via2 ;
        RECT 2898.090 2433.920 2898.370 2434.200 ;
      LAYER met3 ;
        RECT 2898.065 2434.210 2898.395 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2898.065 2433.910 2924.800 2434.210 ;
        RECT 2898.065 2433.895 2898.395 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 922.370 3221.400 922.690 3221.460 ;
        RECT 2617.930 3221.400 2618.250 3221.460 ;
        RECT 922.370 3221.260 2618.250 3221.400 ;
        RECT 922.370 3221.200 922.690 3221.260 ;
        RECT 2617.930 3221.200 2618.250 3221.260 ;
        RECT 2617.930 2670.260 2618.250 2670.320 ;
        RECT 2898.990 2670.260 2899.310 2670.320 ;
        RECT 2617.930 2670.120 2899.310 2670.260 ;
        RECT 2617.930 2670.060 2618.250 2670.120 ;
        RECT 2898.990 2670.060 2899.310 2670.120 ;
      LAYER via ;
        RECT 922.400 3221.200 922.660 3221.460 ;
        RECT 2617.960 3221.200 2618.220 3221.460 ;
        RECT 2617.960 2670.060 2618.220 2670.320 ;
        RECT 2899.020 2670.060 2899.280 2670.320 ;
      LAYER met2 ;
        RECT 922.400 3221.170 922.660 3221.490 ;
        RECT 2617.960 3221.170 2618.220 3221.490 ;
        RECT 922.460 3220.000 922.600 3221.170 ;
        RECT 922.440 3216.000 922.720 3220.000 ;
        RECT 2618.020 2670.350 2618.160 3221.170 ;
        RECT 2617.960 2670.030 2618.220 2670.350 ;
        RECT 2899.020 2670.030 2899.280 2670.350 ;
        RECT 2899.080 2669.525 2899.220 2670.030 ;
        RECT 2899.010 2669.155 2899.290 2669.525 ;
      LAYER via2 ;
        RECT 2899.010 2669.200 2899.290 2669.480 ;
      LAYER met3 ;
        RECT 2898.985 2669.490 2899.315 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2898.985 2669.190 2924.800 2669.490 ;
        RECT 2898.985 2669.175 2899.315 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 985.390 3221.740 985.710 3221.800 ;
        RECT 2617.470 3221.740 2617.790 3221.800 ;
        RECT 985.390 3221.600 2617.790 3221.740 ;
        RECT 985.390 3221.540 985.710 3221.600 ;
        RECT 2617.470 3221.540 2617.790 3221.600 ;
        RECT 2617.470 2904.860 2617.790 2904.920 ;
        RECT 2898.990 2904.860 2899.310 2904.920 ;
        RECT 2617.470 2904.720 2899.310 2904.860 ;
        RECT 2617.470 2904.660 2617.790 2904.720 ;
        RECT 2898.990 2904.660 2899.310 2904.720 ;
      LAYER via ;
        RECT 985.420 3221.540 985.680 3221.800 ;
        RECT 2617.500 3221.540 2617.760 3221.800 ;
        RECT 2617.500 2904.660 2617.760 2904.920 ;
        RECT 2899.020 2904.660 2899.280 2904.920 ;
      LAYER met2 ;
        RECT 985.420 3221.510 985.680 3221.830 ;
        RECT 2617.500 3221.510 2617.760 3221.830 ;
        RECT 985.480 3220.000 985.620 3221.510 ;
        RECT 985.460 3216.000 985.740 3220.000 ;
        RECT 2617.560 2904.950 2617.700 3221.510 ;
        RECT 2617.500 2904.630 2617.760 2904.950 ;
        RECT 2899.020 2904.630 2899.280 2904.950 ;
        RECT 2899.080 2904.125 2899.220 2904.630 ;
        RECT 2899.010 2903.755 2899.290 2904.125 ;
      LAYER via2 ;
        RECT 2899.010 2903.800 2899.290 2904.080 ;
      LAYER met3 ;
        RECT 2898.985 2904.090 2899.315 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2898.985 2903.790 2924.800 2904.090 ;
        RECT 2898.985 2903.775 2899.315 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1048.410 3222.080 1048.730 3222.140 ;
        RECT 2617.010 3222.080 2617.330 3222.140 ;
        RECT 1048.410 3221.940 2617.330 3222.080 ;
        RECT 1048.410 3221.880 1048.730 3221.940 ;
        RECT 2617.010 3221.880 2617.330 3221.940 ;
        RECT 2617.010 3139.460 2617.330 3139.520 ;
        RECT 2898.990 3139.460 2899.310 3139.520 ;
        RECT 2617.010 3139.320 2899.310 3139.460 ;
        RECT 2617.010 3139.260 2617.330 3139.320 ;
        RECT 2898.990 3139.260 2899.310 3139.320 ;
      LAYER via ;
        RECT 1048.440 3221.880 1048.700 3222.140 ;
        RECT 2617.040 3221.880 2617.300 3222.140 ;
        RECT 2617.040 3139.260 2617.300 3139.520 ;
        RECT 2899.020 3139.260 2899.280 3139.520 ;
      LAYER met2 ;
        RECT 1048.440 3221.850 1048.700 3222.170 ;
        RECT 2617.040 3221.850 2617.300 3222.170 ;
        RECT 1048.500 3220.000 1048.640 3221.850 ;
        RECT 1048.480 3216.000 1048.760 3220.000 ;
        RECT 2617.100 3139.550 2617.240 3221.850 ;
        RECT 2617.040 3139.230 2617.300 3139.550 ;
        RECT 2899.020 3139.230 2899.280 3139.550 ;
        RECT 2617.100 3139.015 2617.240 3139.230 ;
        RECT 2899.080 3138.725 2899.220 3139.230 ;
        RECT 2899.010 3138.355 2899.290 3138.725 ;
      LAYER via2 ;
        RECT 2899.010 3138.400 2899.290 3138.680 ;
      LAYER met3 ;
        RECT 2898.985 3138.690 2899.315 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2898.985 3138.390 2924.800 3138.690 ;
        RECT 2898.985 3138.375 2899.315 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1117.410 3367.600 1117.730 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 1117.410 3367.460 2901.150 3367.600 ;
        RECT 1117.410 3367.400 1117.730 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
      LAYER via ;
        RECT 1117.440 3367.400 1117.700 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 1117.440 3367.370 1117.700 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 1111.960 3218.850 1112.240 3220.000 ;
        RECT 1117.500 3218.850 1117.640 3367.370 ;
        RECT 1111.960 3218.710 1117.640 3218.850 ;
        RECT 1111.960 3216.000 1112.240 3218.710 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2796.025 3332.765 2796.195 3422.355 ;
        RECT 2795.105 3239.265 2795.275 3284.315 ;
      LAYER mcon ;
        RECT 2796.025 3422.185 2796.195 3422.355 ;
        RECT 2795.105 3284.145 2795.275 3284.315 ;
      LAYER met1 ;
        RECT 2795.490 3443.080 2795.810 3443.140 ;
        RECT 2798.250 3443.080 2798.570 3443.140 ;
        RECT 2795.490 3442.940 2798.570 3443.080 ;
        RECT 2795.490 3442.880 2795.810 3442.940 ;
        RECT 2798.250 3442.880 2798.570 3442.940 ;
        RECT 2795.030 3422.340 2795.350 3422.400 ;
        RECT 2795.965 3422.340 2796.255 3422.385 ;
        RECT 2795.030 3422.200 2796.255 3422.340 ;
        RECT 2795.030 3422.140 2795.350 3422.200 ;
        RECT 2795.965 3422.155 2796.255 3422.200 ;
        RECT 2795.950 3332.920 2796.270 3332.980 ;
        RECT 2795.755 3332.780 2796.270 3332.920 ;
        RECT 2795.950 3332.720 2796.270 3332.780 ;
        RECT 2795.030 3284.300 2795.350 3284.360 ;
        RECT 2794.835 3284.160 2795.350 3284.300 ;
        RECT 2795.030 3284.100 2795.350 3284.160 ;
        RECT 1174.910 3239.420 1175.230 3239.480 ;
        RECT 2795.045 3239.420 2795.335 3239.465 ;
        RECT 1174.910 3239.280 2795.335 3239.420 ;
        RECT 1174.910 3239.220 1175.230 3239.280 ;
        RECT 2795.045 3239.235 2795.335 3239.280 ;
      LAYER via ;
        RECT 2795.520 3442.880 2795.780 3443.140 ;
        RECT 2798.280 3442.880 2798.540 3443.140 ;
        RECT 2795.060 3422.140 2795.320 3422.400 ;
        RECT 2795.980 3332.720 2796.240 3332.980 ;
        RECT 2795.060 3284.100 2795.320 3284.360 ;
        RECT 1174.940 3239.220 1175.200 3239.480 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3443.170 2798.480 3517.600 ;
        RECT 2795.520 3442.850 2795.780 3443.170 ;
        RECT 2798.280 3442.850 2798.540 3443.170 ;
        RECT 2795.580 3429.650 2795.720 3442.850 ;
        RECT 2795.120 3429.510 2795.720 3429.650 ;
        RECT 2795.120 3422.430 2795.260 3429.510 ;
        RECT 2795.060 3422.110 2795.320 3422.430 ;
        RECT 2795.980 3332.690 2796.240 3333.010 ;
        RECT 2796.040 3298.410 2796.180 3332.690 ;
        RECT 2795.120 3298.270 2796.180 3298.410 ;
        RECT 2795.120 3284.390 2795.260 3298.270 ;
        RECT 2795.060 3284.070 2795.320 3284.390 ;
        RECT 1174.940 3239.190 1175.200 3239.510 ;
        RECT 1175.000 3220.000 1175.140 3239.190 ;
        RECT 1174.980 3216.000 1175.260 3220.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2470.345 3332.765 2470.515 3380.875 ;
      LAYER mcon ;
        RECT 2470.345 3380.705 2470.515 3380.875 ;
      LAYER met1 ;
        RECT 2470.270 3380.860 2470.590 3380.920 ;
        RECT 2470.075 3380.720 2470.590 3380.860 ;
        RECT 2470.270 3380.660 2470.590 3380.720 ;
        RECT 2470.285 3332.920 2470.575 3332.965 ;
        RECT 2470.730 3332.920 2471.050 3332.980 ;
        RECT 2470.285 3332.780 2471.050 3332.920 ;
        RECT 2470.285 3332.735 2470.575 3332.780 ;
        RECT 2470.730 3332.720 2471.050 3332.780 ;
        RECT 2470.270 3270.700 2470.590 3270.760 ;
        RECT 2471.190 3270.700 2471.510 3270.760 ;
        RECT 2470.270 3270.560 2471.510 3270.700 ;
        RECT 2470.270 3270.500 2470.590 3270.560 ;
        RECT 2471.190 3270.500 2471.510 3270.560 ;
        RECT 1237.930 3239.760 1238.250 3239.820 ;
        RECT 2470.270 3239.760 2470.590 3239.820 ;
        RECT 1237.930 3239.620 2470.590 3239.760 ;
        RECT 1237.930 3239.560 1238.250 3239.620 ;
        RECT 2470.270 3239.560 2470.590 3239.620 ;
      LAYER via ;
        RECT 2470.300 3380.660 2470.560 3380.920 ;
        RECT 2470.760 3332.720 2471.020 3332.980 ;
        RECT 2470.300 3270.500 2470.560 3270.760 ;
        RECT 2471.220 3270.500 2471.480 3270.760 ;
        RECT 1237.960 3239.560 1238.220 3239.820 ;
        RECT 2470.300 3239.560 2470.560 3239.820 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3430.445 2474.640 3517.230 ;
        RECT 2474.430 3430.075 2474.710 3430.445 ;
        RECT 2471.210 3429.395 2471.490 3429.765 ;
        RECT 2471.280 3394.970 2471.420 3429.395 ;
        RECT 2470.360 3394.830 2471.420 3394.970 ;
        RECT 2470.360 3380.950 2470.500 3394.830 ;
        RECT 2470.300 3380.630 2470.560 3380.950 ;
        RECT 2470.760 3332.690 2471.020 3333.010 ;
        RECT 2470.820 3298.410 2470.960 3332.690 ;
        RECT 2470.820 3298.270 2471.420 3298.410 ;
        RECT 2471.280 3270.790 2471.420 3298.270 ;
        RECT 2470.300 3270.470 2470.560 3270.790 ;
        RECT 2471.220 3270.470 2471.480 3270.790 ;
        RECT 2470.360 3239.850 2470.500 3270.470 ;
        RECT 1237.960 3239.530 1238.220 3239.850 ;
        RECT 2470.300 3239.530 2470.560 3239.850 ;
        RECT 1238.020 3220.000 1238.160 3239.530 ;
        RECT 1238.000 3216.000 1238.280 3220.000 ;
      LAYER via2 ;
        RECT 2474.430 3430.120 2474.710 3430.400 ;
        RECT 2471.210 3429.440 2471.490 3429.720 ;
      LAYER met3 ;
        RECT 2474.405 3430.410 2474.735 3430.425 ;
        RECT 2470.510 3430.110 2474.735 3430.410 ;
        RECT 2470.510 3429.730 2470.810 3430.110 ;
        RECT 2474.405 3430.095 2474.735 3430.110 ;
        RECT 2471.185 3429.730 2471.515 3429.745 ;
        RECT 2470.510 3429.430 2471.515 3429.730 ;
        RECT 2471.185 3429.415 2471.515 3429.430 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2147.425 3332.765 2147.595 3422.355 ;
        RECT 2146.505 3239.945 2146.675 3284.315 ;
      LAYER mcon ;
        RECT 2147.425 3422.185 2147.595 3422.355 ;
        RECT 2146.505 3284.145 2146.675 3284.315 ;
      LAYER met1 ;
        RECT 2146.890 3443.080 2147.210 3443.140 ;
        RECT 2149.190 3443.080 2149.510 3443.140 ;
        RECT 2146.890 3442.940 2149.510 3443.080 ;
        RECT 2146.890 3442.880 2147.210 3442.940 ;
        RECT 2149.190 3442.880 2149.510 3442.940 ;
        RECT 2146.430 3422.340 2146.750 3422.400 ;
        RECT 2147.365 3422.340 2147.655 3422.385 ;
        RECT 2146.430 3422.200 2147.655 3422.340 ;
        RECT 2146.430 3422.140 2146.750 3422.200 ;
        RECT 2147.365 3422.155 2147.655 3422.200 ;
        RECT 2147.350 3332.920 2147.670 3332.980 ;
        RECT 2147.155 3332.780 2147.670 3332.920 ;
        RECT 2147.350 3332.720 2147.670 3332.780 ;
        RECT 2146.430 3284.300 2146.750 3284.360 ;
        RECT 2146.235 3284.160 2146.750 3284.300 ;
        RECT 2146.430 3284.100 2146.750 3284.160 ;
        RECT 1300.950 3240.100 1301.270 3240.160 ;
        RECT 2146.445 3240.100 2146.735 3240.145 ;
        RECT 1300.950 3239.960 2146.735 3240.100 ;
        RECT 1300.950 3239.900 1301.270 3239.960 ;
        RECT 2146.445 3239.915 2146.735 3239.960 ;
      LAYER via ;
        RECT 2146.920 3442.880 2147.180 3443.140 ;
        RECT 2149.220 3442.880 2149.480 3443.140 ;
        RECT 2146.460 3422.140 2146.720 3422.400 ;
        RECT 2147.380 3332.720 2147.640 3332.980 ;
        RECT 2146.460 3284.100 2146.720 3284.360 ;
        RECT 1300.980 3239.900 1301.240 3240.160 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3443.170 2149.420 3517.600 ;
        RECT 2146.920 3442.850 2147.180 3443.170 ;
        RECT 2149.220 3442.850 2149.480 3443.170 ;
        RECT 2146.980 3429.650 2147.120 3442.850 ;
        RECT 2146.520 3429.510 2147.120 3429.650 ;
        RECT 2146.520 3422.430 2146.660 3429.510 ;
        RECT 2146.460 3422.110 2146.720 3422.430 ;
        RECT 2147.380 3332.690 2147.640 3333.010 ;
        RECT 2147.440 3298.410 2147.580 3332.690 ;
        RECT 2146.520 3298.270 2147.580 3298.410 ;
        RECT 2146.520 3284.390 2146.660 3298.270 ;
        RECT 2146.460 3284.070 2146.720 3284.390 ;
        RECT 1300.980 3239.870 1301.240 3240.190 ;
        RECT 1301.040 3220.000 1301.180 3239.870 ;
        RECT 1301.020 3216.000 1301.300 3220.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1821.745 3332.765 1821.915 3380.875 ;
      LAYER mcon ;
        RECT 1821.745 3380.705 1821.915 3380.875 ;
      LAYER met1 ;
        RECT 1821.670 3380.860 1821.990 3380.920 ;
        RECT 1821.475 3380.720 1821.990 3380.860 ;
        RECT 1821.670 3380.660 1821.990 3380.720 ;
        RECT 1821.685 3332.920 1821.975 3332.965 ;
        RECT 1822.130 3332.920 1822.450 3332.980 ;
        RECT 1821.685 3332.780 1822.450 3332.920 ;
        RECT 1821.685 3332.735 1821.975 3332.780 ;
        RECT 1822.130 3332.720 1822.450 3332.780 ;
        RECT 1821.670 3270.700 1821.990 3270.760 ;
        RECT 1822.590 3270.700 1822.910 3270.760 ;
        RECT 1821.670 3270.560 1822.910 3270.700 ;
        RECT 1821.670 3270.500 1821.990 3270.560 ;
        RECT 1822.590 3270.500 1822.910 3270.560 ;
        RECT 1364.430 3240.440 1364.750 3240.500 ;
        RECT 1821.670 3240.440 1821.990 3240.500 ;
        RECT 1364.430 3240.300 1821.990 3240.440 ;
        RECT 1364.430 3240.240 1364.750 3240.300 ;
        RECT 1821.670 3240.240 1821.990 3240.300 ;
      LAYER via ;
        RECT 1821.700 3380.660 1821.960 3380.920 ;
        RECT 1822.160 3332.720 1822.420 3332.980 ;
        RECT 1821.700 3270.500 1821.960 3270.760 ;
        RECT 1822.620 3270.500 1822.880 3270.760 ;
        RECT 1364.460 3240.240 1364.720 3240.500 ;
        RECT 1821.700 3240.240 1821.960 3240.500 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3517.370 1825.120 3517.600 ;
        RECT 1824.980 3517.230 1825.580 3517.370 ;
        RECT 1825.440 3430.445 1825.580 3517.230 ;
        RECT 1825.370 3430.075 1825.650 3430.445 ;
        RECT 1822.610 3429.395 1822.890 3429.765 ;
        RECT 1822.680 3394.970 1822.820 3429.395 ;
        RECT 1821.760 3394.830 1822.820 3394.970 ;
        RECT 1821.760 3380.950 1821.900 3394.830 ;
        RECT 1821.700 3380.630 1821.960 3380.950 ;
        RECT 1822.160 3332.690 1822.420 3333.010 ;
        RECT 1822.220 3298.410 1822.360 3332.690 ;
        RECT 1822.220 3298.270 1822.820 3298.410 ;
        RECT 1822.680 3270.790 1822.820 3298.270 ;
        RECT 1821.700 3270.470 1821.960 3270.790 ;
        RECT 1822.620 3270.470 1822.880 3270.790 ;
        RECT 1821.760 3240.530 1821.900 3270.470 ;
        RECT 1364.460 3240.210 1364.720 3240.530 ;
        RECT 1821.700 3240.210 1821.960 3240.530 ;
        RECT 1364.520 3220.000 1364.660 3240.210 ;
        RECT 1364.500 3216.000 1364.780 3220.000 ;
      LAYER via2 ;
        RECT 1825.370 3430.120 1825.650 3430.400 ;
        RECT 1822.610 3429.440 1822.890 3429.720 ;
      LAYER met3 ;
        RECT 1825.345 3430.410 1825.675 3430.425 ;
        RECT 1821.910 3430.110 1825.675 3430.410 ;
        RECT 1821.910 3429.730 1822.210 3430.110 ;
        RECT 1825.345 3430.095 1825.675 3430.110 ;
        RECT 1822.585 3429.730 1822.915 3429.745 ;
        RECT 1821.910 3429.430 1822.915 3429.730 ;
        RECT 1822.585 3429.415 1822.915 3429.430 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1498.825 3332.765 1498.995 3422.355 ;
        RECT 1498.825 3284.825 1498.995 3298.595 ;
        RECT 1497.905 3240.965 1498.075 3284.315 ;
      LAYER mcon ;
        RECT 1498.825 3422.185 1498.995 3422.355 ;
        RECT 1498.825 3298.425 1498.995 3298.595 ;
        RECT 1497.905 3284.145 1498.075 3284.315 ;
      LAYER met1 ;
        RECT 1498.290 3443.080 1498.610 3443.140 ;
        RECT 1500.590 3443.080 1500.910 3443.140 ;
        RECT 1498.290 3442.940 1500.910 3443.080 ;
        RECT 1498.290 3442.880 1498.610 3442.940 ;
        RECT 1500.590 3442.880 1500.910 3442.940 ;
        RECT 1497.830 3422.340 1498.150 3422.400 ;
        RECT 1498.765 3422.340 1499.055 3422.385 ;
        RECT 1497.830 3422.200 1499.055 3422.340 ;
        RECT 1497.830 3422.140 1498.150 3422.200 ;
        RECT 1498.765 3422.155 1499.055 3422.200 ;
        RECT 1498.750 3332.920 1499.070 3332.980 ;
        RECT 1498.555 3332.780 1499.070 3332.920 ;
        RECT 1498.750 3332.720 1499.070 3332.780 ;
        RECT 1498.750 3298.580 1499.070 3298.640 ;
        RECT 1498.555 3298.440 1499.070 3298.580 ;
        RECT 1498.750 3298.380 1499.070 3298.440 ;
        RECT 1498.290 3284.980 1498.610 3285.040 ;
        RECT 1498.765 3284.980 1499.055 3285.025 ;
        RECT 1498.290 3284.840 1499.055 3284.980 ;
        RECT 1498.290 3284.780 1498.610 3284.840 ;
        RECT 1498.765 3284.795 1499.055 3284.840 ;
        RECT 1497.830 3284.300 1498.150 3284.360 ;
        RECT 1497.635 3284.160 1498.150 3284.300 ;
        RECT 1497.830 3284.100 1498.150 3284.160 ;
        RECT 1427.450 3241.120 1427.770 3241.180 ;
        RECT 1497.845 3241.120 1498.135 3241.165 ;
        RECT 1427.450 3240.980 1498.135 3241.120 ;
        RECT 1427.450 3240.920 1427.770 3240.980 ;
        RECT 1497.845 3240.935 1498.135 3240.980 ;
      LAYER via ;
        RECT 1498.320 3442.880 1498.580 3443.140 ;
        RECT 1500.620 3442.880 1500.880 3443.140 ;
        RECT 1497.860 3422.140 1498.120 3422.400 ;
        RECT 1498.780 3332.720 1499.040 3332.980 ;
        RECT 1498.780 3298.380 1499.040 3298.640 ;
        RECT 1498.320 3284.780 1498.580 3285.040 ;
        RECT 1497.860 3284.100 1498.120 3284.360 ;
        RECT 1427.480 3240.920 1427.740 3241.180 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3443.170 1500.820 3517.600 ;
        RECT 1498.320 3442.850 1498.580 3443.170 ;
        RECT 1500.620 3442.850 1500.880 3443.170 ;
        RECT 1498.380 3429.650 1498.520 3442.850 ;
        RECT 1497.920 3429.510 1498.520 3429.650 ;
        RECT 1497.920 3422.430 1498.060 3429.510 ;
        RECT 1497.860 3422.110 1498.120 3422.430 ;
        RECT 1498.780 3332.690 1499.040 3333.010 ;
        RECT 1498.840 3298.670 1498.980 3332.690 ;
        RECT 1498.780 3298.350 1499.040 3298.670 ;
        RECT 1498.320 3284.810 1498.580 3285.070 ;
        RECT 1497.920 3284.750 1498.580 3284.810 ;
        RECT 1497.920 3284.670 1498.520 3284.750 ;
        RECT 1497.920 3284.390 1498.060 3284.670 ;
        RECT 1497.860 3284.070 1498.120 3284.390 ;
        RECT 1427.480 3240.890 1427.740 3241.210 ;
        RECT 1427.540 3220.000 1427.680 3240.890 ;
        RECT 1427.520 3216.000 1427.800 3220.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 292.170 3216.640 292.490 3216.700 ;
        RECT 2611.950 3216.640 2612.270 3216.700 ;
        RECT 292.170 3216.500 2612.270 3216.640 ;
        RECT 292.170 3216.440 292.490 3216.500 ;
        RECT 2611.950 3216.440 2612.270 3216.500 ;
        RECT 2612.410 324.260 2612.730 324.320 ;
        RECT 2900.830 324.260 2901.150 324.320 ;
        RECT 2612.410 324.120 2901.150 324.260 ;
        RECT 2612.410 324.060 2612.730 324.120 ;
        RECT 2900.830 324.060 2901.150 324.120 ;
      LAYER via ;
        RECT 292.200 3216.440 292.460 3216.700 ;
        RECT 2611.980 3216.440 2612.240 3216.700 ;
        RECT 2612.440 324.060 2612.700 324.320 ;
        RECT 2900.860 324.060 2901.120 324.320 ;
      LAYER met2 ;
        RECT 290.860 3216.810 291.140 3220.000 ;
        RECT 290.860 3216.730 292.400 3216.810 ;
        RECT 290.860 3216.670 292.460 3216.730 ;
        RECT 290.860 3216.000 291.140 3216.670 ;
        RECT 292.200 3216.410 292.460 3216.670 ;
        RECT 2611.980 3216.410 2612.240 3216.730 ;
        RECT 2612.040 330.890 2612.180 3216.410 ;
        RECT 2612.040 330.750 2612.640 330.890 ;
        RECT 2612.500 324.350 2612.640 330.750 ;
        RECT 2612.440 324.030 2612.700 324.350 ;
        RECT 2900.860 324.030 2901.120 324.350 ;
        RECT 2900.920 322.845 2901.060 324.030 ;
        RECT 2900.850 322.475 2901.130 322.845 ;
      LAYER via2 ;
        RECT 2900.850 322.520 2901.130 322.800 ;
      LAYER met3 ;
        RECT 2900.825 322.810 2901.155 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2900.825 322.510 2924.800 322.810 ;
        RECT 2900.825 322.495 2901.155 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1179.510 3240.780 1179.830 3240.840 ;
        RECT 1490.470 3240.780 1490.790 3240.840 ;
        RECT 1179.510 3240.640 1490.790 3240.780 ;
        RECT 1179.510 3240.580 1179.830 3240.640 ;
        RECT 1490.470 3240.580 1490.790 3240.640 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1179.540 3240.580 1179.800 3240.840 ;
        RECT 1490.500 3240.580 1490.760 3240.840 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 3240.870 1179.740 3498.270 ;
        RECT 1179.540 3240.550 1179.800 3240.870 ;
        RECT 1490.500 3240.550 1490.760 3240.870 ;
        RECT 1490.560 3220.000 1490.700 3240.550 ;
        RECT 1490.540 3216.000 1490.820 3220.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3500.880 851.850 3500.940 ;
        RECT 1552.570 3500.880 1552.890 3500.940 ;
        RECT 851.530 3500.740 1552.890 3500.880 ;
        RECT 851.530 3500.680 851.850 3500.740 ;
        RECT 1552.570 3500.680 1552.890 3500.740 ;
      LAYER via ;
        RECT 851.560 3500.680 851.820 3500.940 ;
        RECT 1552.600 3500.680 1552.860 3500.940 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3500.970 851.760 3517.600 ;
        RECT 851.560 3500.650 851.820 3500.970 ;
        RECT 1552.600 3500.650 1552.860 3500.970 ;
        RECT 1552.660 3219.530 1552.800 3500.650 ;
        RECT 1554.020 3219.530 1554.300 3220.000 ;
        RECT 1552.660 3219.390 1554.300 3219.530 ;
        RECT 1554.020 3216.000 1554.300 3219.390 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3503.940 527.550 3504.000 ;
        RECT 1614.670 3503.940 1614.990 3504.000 ;
        RECT 527.230 3503.800 1614.990 3503.940 ;
        RECT 527.230 3503.740 527.550 3503.800 ;
        RECT 1614.670 3503.740 1614.990 3503.800 ;
      LAYER via ;
        RECT 527.260 3503.740 527.520 3504.000 ;
        RECT 1614.700 3503.740 1614.960 3504.000 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3504.030 527.460 3517.600 ;
        RECT 527.260 3503.710 527.520 3504.030 ;
        RECT 1614.700 3503.710 1614.960 3504.030 ;
        RECT 1614.760 3218.850 1614.900 3503.710 ;
        RECT 1617.040 3218.850 1617.320 3220.000 ;
        RECT 1614.760 3218.710 1617.320 3218.850 ;
        RECT 1617.040 3216.000 1617.320 3218.710 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3502.240 202.790 3502.300 ;
        RECT 1676.770 3502.240 1677.090 3502.300 ;
        RECT 202.470 3502.100 1677.090 3502.240 ;
        RECT 202.470 3502.040 202.790 3502.100 ;
        RECT 1676.770 3502.040 1677.090 3502.100 ;
      LAYER via ;
        RECT 202.500 3502.040 202.760 3502.300 ;
        RECT 1676.800 3502.040 1677.060 3502.300 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3502.330 202.700 3517.600 ;
        RECT 202.500 3502.010 202.760 3502.330 ;
        RECT 1676.800 3502.010 1677.060 3502.330 ;
        RECT 1676.860 3218.850 1677.000 3502.010 ;
        RECT 1680.060 3218.850 1680.340 3220.000 ;
        RECT 1676.860 3218.710 1680.340 3218.850 ;
        RECT 1680.060 3216.000 1680.340 3218.710 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 1738.870 3408.740 1739.190 3408.800 ;
        RECT 17.550 3408.600 1739.190 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 1738.870 3408.540 1739.190 3408.600 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 1738.900 3408.540 1739.160 3408.800 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 1738.900 3408.510 1739.160 3408.830 ;
        RECT 1738.960 3218.850 1739.100 3408.510 ;
        RECT 1743.080 3218.850 1743.360 3220.000 ;
        RECT 1738.960 3218.710 1743.360 3218.850 ;
        RECT 1743.080 3216.000 1743.360 3218.710 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 40.550 3220.380 40.870 3220.440 ;
        RECT 1806.490 3220.380 1806.810 3220.440 ;
        RECT 40.550 3220.240 1806.810 3220.380 ;
        RECT 40.550 3220.180 40.870 3220.240 ;
        RECT 1806.490 3220.180 1806.810 3220.240 ;
        RECT 16.630 3124.500 16.950 3124.560 ;
        RECT 40.550 3124.500 40.870 3124.560 ;
        RECT 16.630 3124.360 40.870 3124.500 ;
        RECT 16.630 3124.300 16.950 3124.360 ;
        RECT 40.550 3124.300 40.870 3124.360 ;
      LAYER via ;
        RECT 40.580 3220.180 40.840 3220.440 ;
        RECT 1806.520 3220.180 1806.780 3220.440 ;
        RECT 16.660 3124.300 16.920 3124.560 ;
        RECT 40.580 3124.300 40.840 3124.560 ;
      LAYER met2 ;
        RECT 40.580 3220.150 40.840 3220.470 ;
        RECT 1806.520 3220.150 1806.780 3220.470 ;
        RECT 40.640 3124.590 40.780 3220.150 ;
        RECT 1806.580 3220.000 1806.720 3220.150 ;
        RECT 1806.560 3216.000 1806.840 3220.000 ;
        RECT 16.660 3124.445 16.920 3124.590 ;
        RECT 16.650 3124.075 16.930 3124.445 ;
        RECT 40.580 3124.270 40.840 3124.590 ;
      LAYER via2 ;
        RECT 16.650 3124.120 16.930 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 16.625 3124.410 16.955 3124.425 ;
        RECT -4.800 3124.110 16.955 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 16.625 3124.095 16.955 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 40.090 3220.040 40.410 3220.100 ;
        RECT 1867.670 3220.040 1867.990 3220.100 ;
        RECT 40.090 3219.900 1867.990 3220.040 ;
        RECT 40.090 3219.840 40.410 3219.900 ;
        RECT 1867.670 3219.840 1867.990 3219.900 ;
        RECT 16.170 2840.600 16.490 2840.660 ;
        RECT 40.090 2840.600 40.410 2840.660 ;
        RECT 16.170 2840.460 40.410 2840.600 ;
        RECT 16.170 2840.400 16.490 2840.460 ;
        RECT 40.090 2840.400 40.410 2840.460 ;
      LAYER via ;
        RECT 40.120 3219.840 40.380 3220.100 ;
        RECT 1867.700 3219.840 1867.960 3220.100 ;
        RECT 16.200 2840.400 16.460 2840.660 ;
        RECT 40.120 2840.400 40.380 2840.660 ;
      LAYER met2 ;
        RECT 40.120 3219.810 40.380 3220.130 ;
        RECT 1867.700 3219.810 1867.960 3220.130 ;
        RECT 40.180 2840.690 40.320 3219.810 ;
        RECT 1867.760 3219.530 1867.900 3219.810 ;
        RECT 1869.580 3219.530 1869.860 3220.000 ;
        RECT 1867.760 3219.390 1869.860 3219.530 ;
        RECT 1869.580 3216.000 1869.860 3219.390 ;
        RECT 16.200 2840.370 16.460 2840.690 ;
        RECT 40.120 2840.370 40.380 2840.690 ;
        RECT 16.260 2836.805 16.400 2840.370 ;
        RECT 16.190 2836.435 16.470 2836.805 ;
      LAYER via2 ;
        RECT 16.190 2836.480 16.470 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 16.165 2836.770 16.495 2836.785 ;
        RECT -4.800 2836.470 16.495 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 16.165 2836.455 16.495 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 39.630 3227.520 39.950 3227.580 ;
        RECT 1932.530 3227.520 1932.850 3227.580 ;
        RECT 39.630 3227.380 1932.850 3227.520 ;
        RECT 39.630 3227.320 39.950 3227.380 ;
        RECT 1932.530 3227.320 1932.850 3227.380 ;
        RECT 16.630 2549.900 16.950 2549.960 ;
        RECT 39.630 2549.900 39.950 2549.960 ;
        RECT 16.630 2549.760 39.950 2549.900 ;
        RECT 16.630 2549.700 16.950 2549.760 ;
        RECT 39.630 2549.700 39.950 2549.760 ;
      LAYER via ;
        RECT 39.660 3227.320 39.920 3227.580 ;
        RECT 1932.560 3227.320 1932.820 3227.580 ;
        RECT 16.660 2549.700 16.920 2549.960 ;
        RECT 39.660 2549.700 39.920 2549.960 ;
      LAYER met2 ;
        RECT 39.660 3227.290 39.920 3227.610 ;
        RECT 1932.560 3227.290 1932.820 3227.610 ;
        RECT 39.720 2549.990 39.860 3227.290 ;
        RECT 1932.620 3220.000 1932.760 3227.290 ;
        RECT 1932.600 3216.000 1932.880 3220.000 ;
        RECT 16.660 2549.845 16.920 2549.990 ;
        RECT 16.650 2549.475 16.930 2549.845 ;
        RECT 39.660 2549.670 39.920 2549.990 ;
      LAYER via2 ;
        RECT 16.650 2549.520 16.930 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 16.625 2549.810 16.955 2549.825 ;
        RECT -4.800 2549.510 16.955 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 16.625 2549.495 16.955 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 39.170 3226.840 39.490 3226.900 ;
        RECT 1996.010 3226.840 1996.330 3226.900 ;
        RECT 39.170 3226.700 1996.330 3226.840 ;
        RECT 39.170 3226.640 39.490 3226.700 ;
        RECT 1996.010 3226.640 1996.330 3226.700 ;
        RECT 16.630 2262.600 16.950 2262.660 ;
        RECT 39.170 2262.600 39.490 2262.660 ;
        RECT 16.630 2262.460 39.490 2262.600 ;
        RECT 16.630 2262.400 16.950 2262.460 ;
        RECT 39.170 2262.400 39.490 2262.460 ;
      LAYER via ;
        RECT 39.200 3226.640 39.460 3226.900 ;
        RECT 1996.040 3226.640 1996.300 3226.900 ;
        RECT 16.660 2262.400 16.920 2262.660 ;
        RECT 39.200 2262.400 39.460 2262.660 ;
      LAYER met2 ;
        RECT 39.200 3226.610 39.460 3226.930 ;
        RECT 1996.040 3226.610 1996.300 3226.930 ;
        RECT 39.260 2262.690 39.400 3226.610 ;
        RECT 1996.100 3220.000 1996.240 3226.610 ;
        RECT 1996.080 3216.000 1996.360 3220.000 ;
        RECT 16.660 2262.370 16.920 2262.690 ;
        RECT 39.200 2262.370 39.460 2262.690 ;
        RECT 16.720 2262.205 16.860 2262.370 ;
        RECT 16.650 2261.835 16.930 2262.205 ;
      LAYER via2 ;
        RECT 16.650 2261.880 16.930 2262.160 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 16.625 2262.170 16.955 2262.185 ;
        RECT -4.800 2261.870 16.955 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 16.625 2261.855 16.955 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.710 3226.500 39.030 3226.560 ;
        RECT 2059.030 3226.500 2059.350 3226.560 ;
        RECT 38.710 3226.360 2059.350 3226.500 ;
        RECT 38.710 3226.300 39.030 3226.360 ;
        RECT 2059.030 3226.300 2059.350 3226.360 ;
        RECT 15.250 1976.320 15.570 1976.380 ;
        RECT 38.710 1976.320 39.030 1976.380 ;
        RECT 15.250 1976.180 39.030 1976.320 ;
        RECT 15.250 1976.120 15.570 1976.180 ;
        RECT 38.710 1976.120 39.030 1976.180 ;
      LAYER via ;
        RECT 38.740 3226.300 39.000 3226.560 ;
        RECT 2059.060 3226.300 2059.320 3226.560 ;
        RECT 15.280 1976.120 15.540 1976.380 ;
        RECT 38.740 1976.120 39.000 1976.380 ;
      LAYER met2 ;
        RECT 38.740 3226.270 39.000 3226.590 ;
        RECT 2059.060 3226.270 2059.320 3226.590 ;
        RECT 38.800 1976.410 38.940 3226.270 ;
        RECT 2059.120 3220.000 2059.260 3226.270 ;
        RECT 2059.100 3216.000 2059.380 3220.000 ;
        RECT 15.280 1976.090 15.540 1976.410 ;
        RECT 38.740 1976.090 39.000 1976.410 ;
        RECT 15.340 1975.245 15.480 1976.090 ;
        RECT 15.270 1974.875 15.550 1975.245 ;
      LAYER via2 ;
        RECT 15.270 1974.920 15.550 1975.200 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 15.245 1975.210 15.575 1975.225 ;
        RECT -4.800 1974.910 15.575 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 15.245 1974.895 15.575 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 353.810 3224.120 354.130 3224.180 ;
        RECT 2612.410 3224.120 2612.730 3224.180 ;
        RECT 353.810 3223.980 2612.730 3224.120 ;
        RECT 353.810 3223.920 354.130 3223.980 ;
        RECT 2612.410 3223.920 2612.730 3223.980 ;
        RECT 2612.410 558.860 2612.730 558.920 ;
        RECT 2898.070 558.860 2898.390 558.920 ;
        RECT 2612.410 558.720 2898.390 558.860 ;
        RECT 2612.410 558.660 2612.730 558.720 ;
        RECT 2898.070 558.660 2898.390 558.720 ;
      LAYER via ;
        RECT 353.840 3223.920 354.100 3224.180 ;
        RECT 2612.440 3223.920 2612.700 3224.180 ;
        RECT 2612.440 558.660 2612.700 558.920 ;
        RECT 2898.100 558.660 2898.360 558.920 ;
      LAYER met2 ;
        RECT 353.840 3223.890 354.100 3224.210 ;
        RECT 2612.440 3223.890 2612.700 3224.210 ;
        RECT 353.900 3220.000 354.040 3223.890 ;
        RECT 353.880 3216.000 354.160 3220.000 ;
        RECT 2612.500 558.950 2612.640 3223.890 ;
        RECT 2612.440 558.630 2612.700 558.950 ;
        RECT 2898.100 558.630 2898.360 558.950 ;
        RECT 2898.160 557.445 2898.300 558.630 ;
        RECT 2898.090 557.075 2898.370 557.445 ;
      LAYER via2 ;
        RECT 2898.090 557.120 2898.370 557.400 ;
      LAYER met3 ;
        RECT 2898.065 557.410 2898.395 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.065 557.110 2924.800 557.410 ;
        RECT 2898.065 557.095 2898.395 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 3225.820 38.570 3225.880 ;
        RECT 2122.050 3225.820 2122.370 3225.880 ;
        RECT 38.250 3225.680 2122.370 3225.820 ;
        RECT 38.250 3225.620 38.570 3225.680 ;
        RECT 2122.050 3225.620 2122.370 3225.680 ;
        RECT 15.710 1689.020 16.030 1689.080 ;
        RECT 38.250 1689.020 38.570 1689.080 ;
        RECT 15.710 1688.880 38.570 1689.020 ;
        RECT 15.710 1688.820 16.030 1688.880 ;
        RECT 38.250 1688.820 38.570 1688.880 ;
      LAYER via ;
        RECT 38.280 3225.620 38.540 3225.880 ;
        RECT 2122.080 3225.620 2122.340 3225.880 ;
        RECT 15.740 1688.820 16.000 1689.080 ;
        RECT 38.280 1688.820 38.540 1689.080 ;
      LAYER met2 ;
        RECT 38.280 3225.590 38.540 3225.910 ;
        RECT 2122.080 3225.590 2122.340 3225.910 ;
        RECT 38.340 1689.110 38.480 3225.590 ;
        RECT 2122.140 3220.000 2122.280 3225.590 ;
        RECT 2122.120 3216.000 2122.400 3220.000 ;
        RECT 15.740 1688.790 16.000 1689.110 ;
        RECT 38.280 1688.790 38.540 1689.110 ;
        RECT 15.800 1687.605 15.940 1688.790 ;
        RECT 15.730 1687.235 16.010 1687.605 ;
      LAYER via2 ;
        RECT 15.730 1687.280 16.010 1687.560 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 15.705 1687.570 16.035 1687.585 ;
        RECT -4.800 1687.270 16.035 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 15.705 1687.255 16.035 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 46.070 3225.140 46.390 3225.200 ;
        RECT 2185.070 3225.140 2185.390 3225.200 ;
        RECT 46.070 3225.000 2185.390 3225.140 ;
        RECT 46.070 3224.940 46.390 3225.000 ;
        RECT 2185.070 3224.940 2185.390 3225.000 ;
        RECT 18.010 1474.820 18.330 1474.880 ;
        RECT 46.070 1474.820 46.390 1474.880 ;
        RECT 18.010 1474.680 46.390 1474.820 ;
        RECT 18.010 1474.620 18.330 1474.680 ;
        RECT 46.070 1474.620 46.390 1474.680 ;
      LAYER via ;
        RECT 46.100 3224.940 46.360 3225.200 ;
        RECT 2185.100 3224.940 2185.360 3225.200 ;
        RECT 18.040 1474.620 18.300 1474.880 ;
        RECT 46.100 1474.620 46.360 1474.880 ;
      LAYER met2 ;
        RECT 46.100 3224.910 46.360 3225.230 ;
        RECT 2185.100 3224.910 2185.360 3225.230 ;
        RECT 46.160 1474.910 46.300 3224.910 ;
        RECT 2185.160 3220.000 2185.300 3224.910 ;
        RECT 2185.140 3216.000 2185.420 3220.000 ;
        RECT 18.040 1474.590 18.300 1474.910 ;
        RECT 46.100 1474.590 46.360 1474.910 ;
        RECT 18.100 1472.045 18.240 1474.590 ;
        RECT 18.030 1471.675 18.310 1472.045 ;
      LAYER via2 ;
        RECT 18.030 1471.720 18.310 1472.000 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 18.005 1472.010 18.335 1472.025 ;
        RECT -4.800 1471.710 18.335 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 18.005 1471.695 18.335 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 31.810 3224.460 32.130 3224.520 ;
        RECT 2248.550 3224.460 2248.870 3224.520 ;
        RECT 31.810 3224.320 2248.870 3224.460 ;
        RECT 31.810 3224.260 32.130 3224.320 ;
        RECT 2248.550 3224.260 2248.870 3224.320 ;
        RECT 15.710 1256.540 16.030 1256.600 ;
        RECT 31.810 1256.540 32.130 1256.600 ;
        RECT 15.710 1256.400 32.130 1256.540 ;
        RECT 15.710 1256.340 16.030 1256.400 ;
        RECT 31.810 1256.340 32.130 1256.400 ;
      LAYER via ;
        RECT 31.840 3224.260 32.100 3224.520 ;
        RECT 2248.580 3224.260 2248.840 3224.520 ;
        RECT 15.740 1256.340 16.000 1256.600 ;
        RECT 31.840 1256.340 32.100 1256.600 ;
      LAYER met2 ;
        RECT 31.840 3224.230 32.100 3224.550 ;
        RECT 2248.580 3224.230 2248.840 3224.550 ;
        RECT 31.900 1256.630 32.040 3224.230 ;
        RECT 2248.640 3220.000 2248.780 3224.230 ;
        RECT 2248.620 3216.000 2248.900 3220.000 ;
        RECT 15.740 1256.485 16.000 1256.630 ;
        RECT 15.730 1256.115 16.010 1256.485 ;
        RECT 31.840 1256.310 32.100 1256.630 ;
      LAYER via2 ;
        RECT 15.730 1256.160 16.010 1256.440 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 15.705 1256.450 16.035 1256.465 ;
        RECT -4.800 1256.150 16.035 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 15.705 1256.135 16.035 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 37.790 3223.780 38.110 3223.840 ;
        RECT 2311.570 3223.780 2311.890 3223.840 ;
        RECT 37.790 3223.640 2311.890 3223.780 ;
        RECT 37.790 3223.580 38.110 3223.640 ;
        RECT 2311.570 3223.580 2311.890 3223.640 ;
        RECT 16.630 1040.980 16.950 1041.040 ;
        RECT 37.790 1040.980 38.110 1041.040 ;
        RECT 16.630 1040.840 38.110 1040.980 ;
        RECT 16.630 1040.780 16.950 1040.840 ;
        RECT 37.790 1040.780 38.110 1040.840 ;
      LAYER via ;
        RECT 37.820 3223.580 38.080 3223.840 ;
        RECT 2311.600 3223.580 2311.860 3223.840 ;
        RECT 16.660 1040.780 16.920 1041.040 ;
        RECT 37.820 1040.780 38.080 1041.040 ;
      LAYER met2 ;
        RECT 37.820 3223.550 38.080 3223.870 ;
        RECT 2311.600 3223.550 2311.860 3223.870 ;
        RECT 37.880 1041.070 38.020 3223.550 ;
        RECT 2311.660 3220.000 2311.800 3223.550 ;
        RECT 2311.640 3216.000 2311.920 3220.000 ;
        RECT 16.660 1040.925 16.920 1041.070 ;
        RECT 16.650 1040.555 16.930 1040.925 ;
        RECT 37.820 1040.750 38.080 1041.070 ;
      LAYER via2 ;
        RECT 16.650 1040.600 16.930 1040.880 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 16.625 1040.890 16.955 1040.905 ;
        RECT -4.800 1040.590 16.955 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 16.625 1040.575 16.955 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 45.610 3223.440 45.930 3223.500 ;
        RECT 2374.590 3223.440 2374.910 3223.500 ;
        RECT 45.610 3223.300 2374.910 3223.440 ;
        RECT 45.610 3223.240 45.930 3223.300 ;
        RECT 2374.590 3223.240 2374.910 3223.300 ;
        RECT 15.710 826.100 16.030 826.160 ;
        RECT 45.610 826.100 45.930 826.160 ;
        RECT 15.710 825.960 45.930 826.100 ;
        RECT 15.710 825.900 16.030 825.960 ;
        RECT 45.610 825.900 45.930 825.960 ;
      LAYER via ;
        RECT 45.640 3223.240 45.900 3223.500 ;
        RECT 2374.620 3223.240 2374.880 3223.500 ;
        RECT 15.740 825.900 16.000 826.160 ;
        RECT 45.640 825.900 45.900 826.160 ;
      LAYER met2 ;
        RECT 45.640 3223.210 45.900 3223.530 ;
        RECT 2374.620 3223.210 2374.880 3223.530 ;
        RECT 45.700 826.190 45.840 3223.210 ;
        RECT 2374.680 3220.000 2374.820 3223.210 ;
        RECT 2374.660 3216.000 2374.940 3220.000 ;
        RECT 15.740 825.870 16.000 826.190 ;
        RECT 45.640 825.870 45.900 826.190 ;
        RECT 15.800 825.365 15.940 825.870 ;
        RECT 15.730 824.995 16.010 825.365 ;
      LAYER via2 ;
        RECT 15.730 825.040 16.010 825.320 ;
      LAYER met3 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 15.705 825.330 16.035 825.345 ;
        RECT -4.800 825.030 16.035 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 15.705 825.015 16.035 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 45.150 3223.100 45.470 3223.160 ;
        RECT 2438.070 3223.100 2438.390 3223.160 ;
        RECT 45.150 3222.960 2438.390 3223.100 ;
        RECT 45.150 3222.900 45.470 3222.960 ;
        RECT 2438.070 3222.900 2438.390 3222.960 ;
        RECT 14.790 613.940 15.110 614.000 ;
        RECT 45.150 613.940 45.470 614.000 ;
        RECT 14.790 613.800 45.470 613.940 ;
        RECT 14.790 613.740 15.110 613.800 ;
        RECT 45.150 613.740 45.470 613.800 ;
      LAYER via ;
        RECT 45.180 3222.900 45.440 3223.160 ;
        RECT 2438.100 3222.900 2438.360 3223.160 ;
        RECT 14.820 613.740 15.080 614.000 ;
        RECT 45.180 613.740 45.440 614.000 ;
      LAYER met2 ;
        RECT 45.180 3222.870 45.440 3223.190 ;
        RECT 2438.100 3222.870 2438.360 3223.190 ;
        RECT 45.240 614.030 45.380 3222.870 ;
        RECT 2438.160 3220.000 2438.300 3222.870 ;
        RECT 2438.140 3216.000 2438.420 3220.000 ;
        RECT 14.820 613.710 15.080 614.030 ;
        RECT 45.180 613.710 45.440 614.030 ;
        RECT 14.880 610.485 15.020 613.710 ;
        RECT 14.810 610.115 15.090 610.485 ;
      LAYER via2 ;
        RECT 14.810 610.160 15.090 610.440 ;
      LAYER met3 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 14.785 610.450 15.115 610.465 ;
        RECT -4.800 610.150 15.115 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 14.785 610.135 15.115 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.690 3222.420 45.010 3222.480 ;
        RECT 2501.090 3222.420 2501.410 3222.480 ;
        RECT 44.690 3222.280 2501.410 3222.420 ;
        RECT 44.690 3222.220 45.010 3222.280 ;
        RECT 2501.090 3222.220 2501.410 3222.280 ;
        RECT 15.250 399.400 15.570 399.460 ;
        RECT 44.690 399.400 45.010 399.460 ;
        RECT 15.250 399.260 45.010 399.400 ;
        RECT 15.250 399.200 15.570 399.260 ;
        RECT 44.690 399.200 45.010 399.260 ;
      LAYER via ;
        RECT 44.720 3222.220 44.980 3222.480 ;
        RECT 2501.120 3222.220 2501.380 3222.480 ;
        RECT 15.280 399.200 15.540 399.460 ;
        RECT 44.720 399.200 44.980 399.460 ;
      LAYER met2 ;
        RECT 44.720 3222.190 44.980 3222.510 ;
        RECT 2501.120 3222.190 2501.380 3222.510 ;
        RECT 44.780 399.490 44.920 3222.190 ;
        RECT 2501.180 3220.000 2501.320 3222.190 ;
        RECT 2501.160 3216.000 2501.440 3220.000 ;
        RECT 15.280 399.170 15.540 399.490 ;
        RECT 44.720 399.170 44.980 399.490 ;
        RECT 15.340 394.925 15.480 399.170 ;
        RECT 15.270 394.555 15.550 394.925 ;
      LAYER via2 ;
        RECT 15.270 394.600 15.550 394.880 ;
      LAYER met3 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 15.245 394.890 15.575 394.905 ;
        RECT -4.800 394.590 15.575 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 15.245 394.575 15.575 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 127.490 3222.760 127.810 3222.820 ;
        RECT 2564.110 3222.760 2564.430 3222.820 ;
        RECT 127.490 3222.620 2564.430 3222.760 ;
        RECT 127.490 3222.560 127.810 3222.620 ;
        RECT 2564.110 3222.560 2564.430 3222.620 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 127.490 179.420 127.810 179.480 ;
        RECT 17.090 179.280 127.810 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 127.490 179.220 127.810 179.280 ;
      LAYER via ;
        RECT 127.520 3222.560 127.780 3222.820 ;
        RECT 2564.140 3222.560 2564.400 3222.820 ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 127.520 179.220 127.780 179.480 ;
      LAYER met2 ;
        RECT 127.520 3222.530 127.780 3222.850 ;
        RECT 2564.140 3222.530 2564.400 3222.850 ;
        RECT 127.580 179.510 127.720 3222.530 ;
        RECT 2564.200 3220.000 2564.340 3222.530 ;
        RECT 2564.180 3216.000 2564.460 3220.000 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 127.520 179.190 127.780 179.510 ;
      LAYER via2 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 416.830 3224.800 417.150 3224.860 ;
        RECT 2612.870 3224.800 2613.190 3224.860 ;
        RECT 416.830 3224.660 2613.190 3224.800 ;
        RECT 416.830 3224.600 417.150 3224.660 ;
        RECT 2612.870 3224.600 2613.190 3224.660 ;
        RECT 2612.870 793.460 2613.190 793.520 ;
        RECT 2900.830 793.460 2901.150 793.520 ;
        RECT 2612.870 793.320 2901.150 793.460 ;
        RECT 2612.870 793.260 2613.190 793.320 ;
        RECT 2900.830 793.260 2901.150 793.320 ;
      LAYER via ;
        RECT 416.860 3224.600 417.120 3224.860 ;
        RECT 2612.900 3224.600 2613.160 3224.860 ;
        RECT 2612.900 793.260 2613.160 793.520 ;
        RECT 2900.860 793.260 2901.120 793.520 ;
      LAYER met2 ;
        RECT 416.860 3224.570 417.120 3224.890 ;
        RECT 2612.900 3224.570 2613.160 3224.890 ;
        RECT 416.920 3220.000 417.060 3224.570 ;
        RECT 416.900 3216.000 417.180 3220.000 ;
        RECT 2612.960 793.550 2613.100 3224.570 ;
        RECT 2612.900 793.230 2613.160 793.550 ;
        RECT 2900.860 793.230 2901.120 793.550 ;
        RECT 2900.920 792.045 2901.060 793.230 ;
        RECT 2900.850 791.675 2901.130 792.045 ;
      LAYER via2 ;
        RECT 2900.850 791.720 2901.130 792.000 ;
      LAYER met3 ;
        RECT 2900.825 792.010 2901.155 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2900.825 791.710 2924.800 792.010 ;
        RECT 2900.825 791.695 2901.155 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 481.690 3217.660 482.010 3217.720 ;
        RECT 2619.310 3217.660 2619.630 3217.720 ;
        RECT 481.690 3217.520 2619.630 3217.660 ;
        RECT 481.690 3217.460 482.010 3217.520 ;
        RECT 2619.310 3217.460 2619.630 3217.520 ;
        RECT 2619.310 1028.060 2619.630 1028.120 ;
        RECT 2900.830 1028.060 2901.150 1028.120 ;
        RECT 2619.310 1027.920 2901.150 1028.060 ;
        RECT 2619.310 1027.860 2619.630 1027.920 ;
        RECT 2900.830 1027.860 2901.150 1027.920 ;
      LAYER via ;
        RECT 481.720 3217.460 481.980 3217.720 ;
        RECT 2619.340 3217.460 2619.600 3217.720 ;
        RECT 2619.340 1027.860 2619.600 1028.120 ;
        RECT 2900.860 1027.860 2901.120 1028.120 ;
      LAYER met2 ;
        RECT 480.380 3217.490 480.660 3220.000 ;
        RECT 481.720 3217.490 481.980 3217.750 ;
        RECT 480.380 3217.430 481.980 3217.490 ;
        RECT 2619.340 3217.430 2619.600 3217.750 ;
        RECT 480.380 3217.350 481.920 3217.430 ;
        RECT 480.380 3216.000 480.660 3217.350 ;
        RECT 2619.400 1028.150 2619.540 3217.430 ;
        RECT 2619.340 1027.830 2619.600 1028.150 ;
        RECT 2900.860 1027.830 2901.120 1028.150 ;
        RECT 2900.920 1026.645 2901.060 1027.830 ;
        RECT 2900.850 1026.275 2901.130 1026.645 ;
      LAYER via2 ;
        RECT 2900.850 1026.320 2901.130 1026.600 ;
      LAYER met3 ;
        RECT 2900.825 1026.610 2901.155 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2900.825 1026.310 2924.800 1026.610 ;
        RECT 2900.825 1026.295 2901.155 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 543.330 3225.480 543.650 3225.540 ;
        RECT 2619.770 3225.480 2620.090 3225.540 ;
        RECT 543.330 3225.340 2620.090 3225.480 ;
        RECT 543.330 3225.280 543.650 3225.340 ;
        RECT 2619.770 3225.280 2620.090 3225.340 ;
        RECT 2619.770 1262.660 2620.090 1262.720 ;
        RECT 2898.530 1262.660 2898.850 1262.720 ;
        RECT 2619.770 1262.520 2898.850 1262.660 ;
        RECT 2619.770 1262.460 2620.090 1262.520 ;
        RECT 2898.530 1262.460 2898.850 1262.520 ;
      LAYER via ;
        RECT 543.360 3225.280 543.620 3225.540 ;
        RECT 2619.800 3225.280 2620.060 3225.540 ;
        RECT 2619.800 1262.460 2620.060 1262.720 ;
        RECT 2898.560 1262.460 2898.820 1262.720 ;
      LAYER met2 ;
        RECT 543.360 3225.250 543.620 3225.570 ;
        RECT 2619.800 3225.250 2620.060 3225.570 ;
        RECT 543.420 3220.000 543.560 3225.250 ;
        RECT 543.400 3216.000 543.680 3220.000 ;
        RECT 2619.860 1262.750 2620.000 3225.250 ;
        RECT 2619.800 1262.430 2620.060 1262.750 ;
        RECT 2898.560 1262.430 2898.820 1262.750 ;
        RECT 2898.620 1261.245 2898.760 1262.430 ;
        RECT 2898.550 1260.875 2898.830 1261.245 ;
      LAYER via2 ;
        RECT 2898.550 1260.920 2898.830 1261.200 ;
      LAYER met3 ;
        RECT 2898.525 1261.210 2898.855 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.525 1260.910 2924.800 1261.210 ;
        RECT 2898.525 1260.895 2898.855 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 3218.340 607.130 3218.400 ;
        RECT 2620.230 3218.340 2620.550 3218.400 ;
        RECT 606.810 3218.200 2620.550 3218.340 ;
        RECT 606.810 3218.140 607.130 3218.200 ;
        RECT 2620.230 3218.140 2620.550 3218.200 ;
        RECT 2620.230 1497.260 2620.550 1497.320 ;
        RECT 2900.830 1497.260 2901.150 1497.320 ;
        RECT 2620.230 1497.120 2901.150 1497.260 ;
        RECT 2620.230 1497.060 2620.550 1497.120 ;
        RECT 2900.830 1497.060 2901.150 1497.120 ;
      LAYER via ;
        RECT 606.840 3218.140 607.100 3218.400 ;
        RECT 2620.260 3218.140 2620.520 3218.400 ;
        RECT 2620.260 1497.060 2620.520 1497.320 ;
        RECT 2900.860 1497.060 2901.120 1497.320 ;
      LAYER met2 ;
        RECT 606.420 3218.170 606.700 3220.000 ;
        RECT 606.840 3218.170 607.100 3218.430 ;
        RECT 606.420 3218.110 607.100 3218.170 ;
        RECT 2620.260 3218.110 2620.520 3218.430 ;
        RECT 606.420 3218.030 607.040 3218.110 ;
        RECT 606.420 3216.000 606.700 3218.030 ;
        RECT 2620.320 1497.350 2620.460 3218.110 ;
        RECT 2620.260 1497.030 2620.520 1497.350 ;
        RECT 2900.860 1497.030 2901.120 1497.350 ;
        RECT 2900.920 1495.845 2901.060 1497.030 ;
        RECT 2900.850 1495.475 2901.130 1495.845 ;
      LAYER via2 ;
        RECT 2900.850 1495.520 2901.130 1495.800 ;
      LAYER met3 ;
        RECT 2900.825 1495.810 2901.155 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2900.825 1495.510 2924.800 1495.810 ;
        RECT 2900.825 1495.495 2901.155 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 669.830 3227.180 670.150 3227.240 ;
        RECT 2620.690 3227.180 2621.010 3227.240 ;
        RECT 669.830 3227.040 2621.010 3227.180 ;
        RECT 669.830 3226.980 670.150 3227.040 ;
        RECT 2620.690 3226.980 2621.010 3227.040 ;
        RECT 2620.690 1731.860 2621.010 1731.920 ;
        RECT 2898.070 1731.860 2898.390 1731.920 ;
        RECT 2620.690 1731.720 2898.390 1731.860 ;
        RECT 2620.690 1731.660 2621.010 1731.720 ;
        RECT 2898.070 1731.660 2898.390 1731.720 ;
      LAYER via ;
        RECT 669.860 3226.980 670.120 3227.240 ;
        RECT 2620.720 3226.980 2620.980 3227.240 ;
        RECT 2620.720 1731.660 2620.980 1731.920 ;
        RECT 2898.100 1731.660 2898.360 1731.920 ;
      LAYER met2 ;
        RECT 669.860 3226.950 670.120 3227.270 ;
        RECT 2620.720 3226.950 2620.980 3227.270 ;
        RECT 669.920 3220.000 670.060 3226.950 ;
        RECT 669.900 3216.000 670.180 3220.000 ;
        RECT 2620.780 1731.950 2620.920 3226.950 ;
        RECT 2620.720 1731.630 2620.980 1731.950 ;
        RECT 2898.100 1731.630 2898.360 1731.950 ;
        RECT 2898.160 1730.445 2898.300 1731.630 ;
        RECT 2898.090 1730.075 2898.370 1730.445 ;
      LAYER via2 ;
        RECT 2898.090 1730.120 2898.370 1730.400 ;
      LAYER met3 ;
        RECT 2898.065 1730.410 2898.395 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2898.065 1730.110 2924.800 1730.410 ;
        RECT 2898.065 1730.095 2898.395 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 734.690 3219.360 735.010 3219.420 ;
        RECT 2621.150 3219.360 2621.470 3219.420 ;
        RECT 734.690 3219.220 2621.470 3219.360 ;
        RECT 734.690 3219.160 735.010 3219.220 ;
        RECT 2621.150 3219.160 2621.470 3219.220 ;
        RECT 2621.150 1966.460 2621.470 1966.520 ;
        RECT 2898.070 1966.460 2898.390 1966.520 ;
        RECT 2621.150 1966.320 2898.390 1966.460 ;
        RECT 2621.150 1966.260 2621.470 1966.320 ;
        RECT 2898.070 1966.260 2898.390 1966.320 ;
      LAYER via ;
        RECT 734.720 3219.160 734.980 3219.420 ;
        RECT 2621.180 3219.160 2621.440 3219.420 ;
        RECT 2621.180 1966.260 2621.440 1966.520 ;
        RECT 2898.100 1966.260 2898.360 1966.520 ;
      LAYER met2 ;
        RECT 732.920 3219.530 733.200 3220.000 ;
        RECT 732.920 3219.450 734.920 3219.530 ;
        RECT 732.920 3219.390 734.980 3219.450 ;
        RECT 732.920 3216.000 733.200 3219.390 ;
        RECT 734.720 3219.130 734.980 3219.390 ;
        RECT 2621.180 3219.130 2621.440 3219.450 ;
        RECT 2621.240 1966.550 2621.380 3219.130 ;
        RECT 2621.180 1966.230 2621.440 1966.550 ;
        RECT 2898.100 1966.230 2898.360 1966.550 ;
        RECT 2898.160 1965.045 2898.300 1966.230 ;
        RECT 2898.090 1964.675 2898.370 1965.045 ;
      LAYER via2 ;
        RECT 2898.090 1964.720 2898.370 1965.000 ;
      LAYER met3 ;
        RECT 2898.065 1965.010 2898.395 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2898.065 1964.710 2924.800 1965.010 ;
        RECT 2898.065 1964.695 2898.395 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 795.870 3228.200 796.190 3228.260 ;
        RECT 2628.050 3228.200 2628.370 3228.260 ;
        RECT 795.870 3228.060 2628.370 3228.200 ;
        RECT 795.870 3228.000 796.190 3228.060 ;
        RECT 2628.050 3228.000 2628.370 3228.060 ;
        RECT 2628.050 2201.060 2628.370 2201.120 ;
        RECT 2898.070 2201.060 2898.390 2201.120 ;
        RECT 2628.050 2200.920 2898.390 2201.060 ;
        RECT 2628.050 2200.860 2628.370 2200.920 ;
        RECT 2898.070 2200.860 2898.390 2200.920 ;
      LAYER via ;
        RECT 795.900 3228.000 796.160 3228.260 ;
        RECT 2628.080 3228.000 2628.340 3228.260 ;
        RECT 2628.080 2200.860 2628.340 2201.120 ;
        RECT 2898.100 2200.860 2898.360 2201.120 ;
      LAYER met2 ;
        RECT 795.900 3227.970 796.160 3228.290 ;
        RECT 2628.080 3227.970 2628.340 3228.290 ;
        RECT 795.960 3220.000 796.100 3227.970 ;
        RECT 795.940 3216.000 796.220 3220.000 ;
        RECT 2628.140 2201.150 2628.280 3227.970 ;
        RECT 2628.080 2200.830 2628.340 2201.150 ;
        RECT 2898.100 2200.830 2898.360 2201.150 ;
        RECT 2898.160 2199.645 2898.300 2200.830 ;
        RECT 2898.090 2199.275 2898.370 2199.645 ;
      LAYER via2 ;
        RECT 2898.090 2199.320 2898.370 2199.600 ;
      LAYER met3 ;
        RECT 2898.065 2199.610 2898.395 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2898.065 2199.310 2924.800 2199.610 ;
        RECT 2898.065 2199.295 2898.395 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 248.540 3216.810 248.820 3220.000 ;
        RECT 249.870 3216.810 250.150 3216.925 ;
        RECT 248.540 3216.670 250.150 3216.810 ;
        RECT 248.540 3216.000 248.820 3216.670 ;
        RECT 249.870 3216.555 250.150 3216.670 ;
        RECT 2623.470 223.195 2623.750 223.565 ;
        RECT 2623.540 202.485 2623.680 223.195 ;
        RECT 2704.430 203.475 2704.710 203.845 ;
        RECT 2623.470 202.115 2623.750 202.485 ;
        RECT 2704.500 201.805 2704.640 203.475 ;
        RECT 2825.410 202.115 2825.690 202.485 ;
        RECT 2704.430 201.435 2704.710 201.805 ;
        RECT 2801.030 200.755 2801.310 201.125 ;
        RECT 2801.100 199.085 2801.240 200.755 ;
        RECT 2825.480 200.445 2825.620 202.115 ;
        RECT 2863.130 200.755 2863.410 201.125 ;
        RECT 2825.410 200.075 2825.690 200.445 ;
        RECT 2863.200 200.330 2863.340 200.755 ;
        RECT 2863.590 200.330 2863.870 200.445 ;
        RECT 2863.200 200.190 2863.870 200.330 ;
        RECT 2863.590 200.075 2863.870 200.190 ;
        RECT 2801.030 198.715 2801.310 199.085 ;
      LAYER via2 ;
        RECT 249.870 3216.600 250.150 3216.880 ;
        RECT 2623.470 223.240 2623.750 223.520 ;
        RECT 2704.430 203.520 2704.710 203.800 ;
        RECT 2623.470 202.160 2623.750 202.440 ;
        RECT 2825.410 202.160 2825.690 202.440 ;
        RECT 2704.430 201.480 2704.710 201.760 ;
        RECT 2801.030 200.800 2801.310 201.080 ;
        RECT 2863.130 200.800 2863.410 201.080 ;
        RECT 2825.410 200.120 2825.690 200.400 ;
        RECT 2863.590 200.120 2863.870 200.400 ;
        RECT 2801.030 198.760 2801.310 199.040 ;
      LAYER met3 ;
        RECT 249.845 3216.890 250.175 3216.905 ;
        RECT 254.190 3216.890 254.570 3216.900 ;
        RECT 249.845 3216.590 254.570 3216.890 ;
        RECT 249.845 3216.575 250.175 3216.590 ;
        RECT 254.190 3216.580 254.570 3216.590 ;
        RECT 1204.550 3215.530 1204.930 3215.540 ;
        RECT 1268.950 3215.530 1269.330 3215.540 ;
        RECT 1204.550 3215.230 1269.330 3215.530 ;
        RECT 1204.550 3215.220 1204.930 3215.230 ;
        RECT 1268.950 3215.220 1269.330 3215.230 ;
        RECT 1322.310 3215.530 1322.690 3215.540 ;
        RECT 1365.550 3215.530 1365.930 3215.540 ;
        RECT 1322.310 3215.230 1365.930 3215.530 ;
        RECT 1322.310 3215.220 1322.690 3215.230 ;
        RECT 1365.550 3215.220 1365.930 3215.230 ;
        RECT 1414.310 3215.530 1414.690 3215.540 ;
        RECT 1558.750 3215.530 1559.130 3215.540 ;
        RECT 1414.310 3215.230 1559.130 3215.530 ;
        RECT 1414.310 3215.220 1414.690 3215.230 ;
        RECT 1558.750 3215.220 1559.130 3215.230 ;
        RECT 1676.510 3215.530 1676.890 3215.540 ;
        RECT 1748.270 3215.530 1748.650 3215.540 ;
        RECT 1676.510 3215.230 1748.650 3215.530 ;
        RECT 1676.510 3215.220 1676.890 3215.230 ;
        RECT 1748.270 3215.220 1748.650 3215.230 ;
        RECT 1753.790 3215.530 1754.170 3215.540 ;
        RECT 1848.550 3215.530 1848.930 3215.540 ;
        RECT 1753.790 3215.230 1848.930 3215.530 ;
        RECT 1753.790 3215.220 1754.170 3215.230 ;
        RECT 1848.550 3215.220 1848.930 3215.230 ;
        RECT 1898.230 3210.770 1898.610 3210.780 ;
        RECT 1956.190 3210.770 1956.570 3210.780 ;
        RECT 1898.230 3210.470 1956.570 3210.770 ;
        RECT 1898.230 3210.460 1898.610 3210.470 ;
        RECT 1956.190 3210.460 1956.570 3210.470 ;
        RECT 379.310 3209.410 379.690 3209.420 ;
        RECT 427.150 3209.410 427.530 3209.420 ;
        RECT 379.310 3209.110 427.530 3209.410 ;
        RECT 379.310 3209.100 379.690 3209.110 ;
        RECT 427.150 3209.100 427.530 3209.110 ;
        RECT 475.910 3209.410 476.290 3209.420 ;
        RECT 523.750 3209.410 524.130 3209.420 ;
        RECT 475.910 3209.110 524.130 3209.410 ;
        RECT 475.910 3209.100 476.290 3209.110 ;
        RECT 523.750 3209.100 524.130 3209.110 ;
        RECT 765.710 3209.410 766.090 3209.420 ;
        RECT 812.630 3209.410 813.010 3209.420 ;
        RECT 765.710 3209.110 813.010 3209.410 ;
        RECT 765.710 3209.100 766.090 3209.110 ;
        RECT 812.630 3209.100 813.010 3209.110 ;
        RECT 820.910 3209.410 821.290 3209.420 ;
        RECT 893.590 3209.410 893.970 3209.420 ;
        RECT 820.910 3209.110 893.970 3209.410 ;
        RECT 820.910 3209.100 821.290 3209.110 ;
        RECT 893.590 3209.100 893.970 3209.110 ;
        RECT 931.310 3209.410 931.690 3209.420 ;
        RECT 979.150 3209.410 979.530 3209.420 ;
        RECT 931.310 3209.110 979.530 3209.410 ;
        RECT 931.310 3209.100 931.690 3209.110 ;
        RECT 979.150 3209.100 979.530 3209.110 ;
        RECT 1993.910 3208.730 1994.290 3208.740 ;
        RECT 2052.790 3208.730 2053.170 3208.740 ;
        RECT 1993.910 3208.430 2053.170 3208.730 ;
        RECT 1993.910 3208.420 1994.290 3208.430 ;
        RECT 2052.790 3208.420 2053.170 3208.430 ;
        RECT 2090.510 3208.730 2090.890 3208.740 ;
        RECT 2138.350 3208.730 2138.730 3208.740 ;
        RECT 2090.510 3208.430 2138.730 3208.730 ;
        RECT 2090.510 3208.420 2090.890 3208.430 ;
        RECT 2138.350 3208.420 2138.730 3208.430 ;
        RECT 2214.710 3208.730 2215.090 3208.740 ;
        RECT 2262.550 3208.730 2262.930 3208.740 ;
        RECT 2214.710 3208.430 2262.930 3208.730 ;
        RECT 2214.710 3208.420 2215.090 3208.430 ;
        RECT 2262.550 3208.420 2262.930 3208.430 ;
        RECT 2312.230 3208.730 2312.610 3208.740 ;
        RECT 2359.150 3208.730 2359.530 3208.740 ;
        RECT 2312.230 3208.430 2359.530 3208.730 ;
        RECT 2312.230 3208.420 2312.610 3208.430 ;
        RECT 2359.150 3208.420 2359.530 3208.430 ;
        RECT 2407.910 3208.730 2408.290 3208.740 ;
        RECT 2455.750 3208.730 2456.130 3208.740 ;
        RECT 2407.910 3208.430 2456.130 3208.730 ;
        RECT 2407.910 3208.420 2408.290 3208.430 ;
        RECT 2455.750 3208.420 2456.130 3208.430 ;
        RECT 2504.510 3208.730 2504.890 3208.740 ;
        RECT 2597.430 3208.730 2597.810 3208.740 ;
        RECT 2504.510 3208.430 2597.810 3208.730 ;
        RECT 2504.510 3208.420 2504.890 3208.430 ;
        RECT 2597.430 3208.420 2597.810 3208.430 ;
        RECT 2611.230 223.530 2611.610 223.540 ;
        RECT 2623.445 223.530 2623.775 223.545 ;
        RECT 2611.230 223.230 2623.775 223.530 ;
        RECT 2611.230 223.220 2611.610 223.230 ;
        RECT 2623.445 223.215 2623.775 223.230 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2916.710 204.870 2924.800 205.170 ;
        RECT 2656.310 203.810 2656.690 203.820 ;
        RECT 2704.405 203.810 2704.735 203.825 ;
        RECT 2656.310 203.510 2704.735 203.810 ;
        RECT 2656.310 203.500 2656.690 203.510 ;
        RECT 2704.405 203.495 2704.735 203.510 ;
        RECT 2623.445 202.450 2623.775 202.465 ;
        RECT 2656.310 202.450 2656.690 202.460 ;
        RECT 2825.385 202.450 2825.715 202.465 ;
        RECT 2623.445 202.150 2656.690 202.450 ;
        RECT 2623.445 202.135 2623.775 202.150 ;
        RECT 2656.310 202.140 2656.690 202.150 ;
        RECT 2801.710 202.150 2825.715 202.450 ;
        RECT 2704.405 201.770 2704.735 201.785 ;
        RECT 2704.405 201.470 2719.210 201.770 ;
        RECT 2704.405 201.455 2704.735 201.470 ;
        RECT 2718.910 200.410 2719.210 201.470 ;
        RECT 2801.005 201.090 2801.335 201.105 ;
        RECT 2801.710 201.090 2802.010 202.150 ;
        RECT 2825.385 202.135 2825.715 202.150 ;
        RECT 2863.105 201.090 2863.435 201.105 ;
        RECT 2916.710 201.090 2917.010 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
        RECT 2801.005 200.790 2802.010 201.090 ;
        RECT 2849.550 200.790 2863.435 201.090 ;
        RECT 2801.005 200.775 2801.335 200.790 ;
        RECT 2752.910 200.410 2753.290 200.420 ;
        RECT 2718.910 200.110 2753.290 200.410 ;
        RECT 2752.910 200.100 2753.290 200.110 ;
        RECT 2825.385 200.410 2825.715 200.425 ;
        RECT 2849.550 200.410 2849.850 200.790 ;
        RECT 2863.105 200.775 2863.435 200.790 ;
        RECT 2884.510 200.790 2917.010 201.090 ;
        RECT 2825.385 200.110 2849.850 200.410 ;
        RECT 2863.565 200.410 2863.895 200.425 ;
        RECT 2884.510 200.410 2884.810 200.790 ;
        RECT 2863.565 200.110 2884.810 200.410 ;
        RECT 2825.385 200.095 2825.715 200.110 ;
        RECT 2863.565 200.095 2863.895 200.110 ;
        RECT 2752.910 199.050 2753.290 199.060 ;
        RECT 2801.005 199.050 2801.335 199.065 ;
        RECT 2752.910 198.750 2801.335 199.050 ;
        RECT 2752.910 198.740 2753.290 198.750 ;
        RECT 2801.005 198.735 2801.335 198.750 ;
      LAYER via3 ;
        RECT 254.220 3216.580 254.540 3216.900 ;
        RECT 1204.580 3215.220 1204.900 3215.540 ;
        RECT 1268.980 3215.220 1269.300 3215.540 ;
        RECT 1322.340 3215.220 1322.660 3215.540 ;
        RECT 1365.580 3215.220 1365.900 3215.540 ;
        RECT 1414.340 3215.220 1414.660 3215.540 ;
        RECT 1558.780 3215.220 1559.100 3215.540 ;
        RECT 1676.540 3215.220 1676.860 3215.540 ;
        RECT 1748.300 3215.220 1748.620 3215.540 ;
        RECT 1753.820 3215.220 1754.140 3215.540 ;
        RECT 1848.580 3215.220 1848.900 3215.540 ;
        RECT 1898.260 3210.460 1898.580 3210.780 ;
        RECT 1956.220 3210.460 1956.540 3210.780 ;
        RECT 379.340 3209.100 379.660 3209.420 ;
        RECT 427.180 3209.100 427.500 3209.420 ;
        RECT 475.940 3209.100 476.260 3209.420 ;
        RECT 523.780 3209.100 524.100 3209.420 ;
        RECT 765.740 3209.100 766.060 3209.420 ;
        RECT 812.660 3209.100 812.980 3209.420 ;
        RECT 820.940 3209.100 821.260 3209.420 ;
        RECT 893.620 3209.100 893.940 3209.420 ;
        RECT 931.340 3209.100 931.660 3209.420 ;
        RECT 979.180 3209.100 979.500 3209.420 ;
        RECT 1993.940 3208.420 1994.260 3208.740 ;
        RECT 2052.820 3208.420 2053.140 3208.740 ;
        RECT 2090.540 3208.420 2090.860 3208.740 ;
        RECT 2138.380 3208.420 2138.700 3208.740 ;
        RECT 2214.740 3208.420 2215.060 3208.740 ;
        RECT 2262.580 3208.420 2262.900 3208.740 ;
        RECT 2312.260 3208.420 2312.580 3208.740 ;
        RECT 2359.180 3208.420 2359.500 3208.740 ;
        RECT 2407.940 3208.420 2408.260 3208.740 ;
        RECT 2455.780 3208.420 2456.100 3208.740 ;
        RECT 2504.540 3208.420 2504.860 3208.740 ;
        RECT 2597.460 3208.420 2597.780 3208.740 ;
        RECT 2611.260 223.220 2611.580 223.540 ;
        RECT 2656.340 203.500 2656.660 203.820 ;
        RECT 2656.340 202.140 2656.660 202.460 ;
        RECT 2752.940 200.100 2753.260 200.420 ;
        RECT 2752.940 198.740 2753.260 199.060 ;
      LAYER met4 ;
        RECT 254.215 3216.575 254.545 3216.905 ;
        RECT 254.230 3208.490 254.530 3216.575 ;
        RECT 1204.575 3215.215 1204.905 3215.545 ;
        RECT 1268.975 3215.215 1269.305 3215.545 ;
        RECT 1322.335 3215.215 1322.665 3215.545 ;
        RECT 1365.575 3215.215 1365.905 3215.545 ;
        RECT 1414.335 3215.215 1414.665 3215.545 ;
        RECT 1558.775 3215.215 1559.105 3215.545 ;
        RECT 1676.535 3215.215 1676.865 3215.545 ;
        RECT 1748.295 3215.215 1748.625 3215.545 ;
        RECT 1753.815 3215.215 1754.145 3215.545 ;
        RECT 1848.575 3215.215 1848.905 3215.545 ;
        RECT 379.335 3209.095 379.665 3209.425 ;
        RECT 427.175 3209.095 427.505 3209.425 ;
        RECT 475.935 3209.095 476.265 3209.425 ;
        RECT 523.775 3209.095 524.105 3209.425 ;
        RECT 765.735 3209.095 766.065 3209.425 ;
        RECT 812.655 3209.095 812.985 3209.425 ;
        RECT 820.935 3209.095 821.265 3209.425 ;
        RECT 893.615 3209.095 893.945 3209.425 ;
        RECT 931.335 3209.095 931.665 3209.425 ;
        RECT 979.175 3209.095 979.505 3209.425 ;
        RECT 379.350 3208.490 379.650 3209.095 ;
        RECT 427.190 3208.490 427.490 3209.095 ;
        RECT 475.950 3208.490 476.250 3209.095 ;
        RECT 523.790 3208.490 524.090 3209.095 ;
        RECT 765.750 3208.490 766.050 3209.095 ;
        RECT 812.670 3208.490 812.970 3209.095 ;
        RECT 820.950 3208.490 821.250 3209.095 ;
        RECT 893.630 3208.490 893.930 3209.095 ;
        RECT 931.350 3208.490 931.650 3209.095 ;
        RECT 979.190 3208.490 979.490 3209.095 ;
        RECT 1204.590 3208.490 1204.890 3215.215 ;
        RECT 1268.990 3208.490 1269.290 3215.215 ;
        RECT 1322.350 3208.490 1322.650 3215.215 ;
        RECT 1365.590 3208.490 1365.890 3215.215 ;
        RECT 1414.350 3208.490 1414.650 3215.215 ;
        RECT 1558.790 3208.490 1559.090 3215.215 ;
        RECT 1676.550 3208.490 1676.850 3215.215 ;
        RECT 1748.310 3208.490 1748.610 3215.215 ;
        RECT 1753.830 3208.490 1754.130 3215.215 ;
        RECT 1848.590 3208.490 1848.890 3215.215 ;
        RECT 1898.255 3210.455 1898.585 3210.785 ;
        RECT 1956.215 3210.455 1956.545 3210.785 ;
        RECT 1898.270 3208.490 1898.570 3210.455 ;
        RECT 1956.230 3208.490 1956.530 3210.455 ;
        RECT 1993.935 3208.490 1994.265 3208.745 ;
        RECT 2052.815 3208.490 2053.145 3208.745 ;
        RECT 2090.535 3208.490 2090.865 3208.745 ;
        RECT 2138.375 3208.490 2138.705 3208.745 ;
        RECT 2214.735 3208.490 2215.065 3208.745 ;
        RECT 2262.575 3208.490 2262.905 3208.745 ;
        RECT 2312.255 3208.490 2312.585 3208.745 ;
        RECT 2359.175 3208.490 2359.505 3208.745 ;
        RECT 2407.935 3208.490 2408.265 3208.745 ;
        RECT 2455.775 3208.490 2456.105 3208.745 ;
        RECT 2504.535 3208.490 2504.865 3208.745 ;
        RECT 2597.455 3208.490 2597.785 3208.745 ;
        RECT 253.790 3207.310 254.970 3208.490 ;
        RECT 378.910 3207.310 380.090 3208.490 ;
        RECT 426.750 3207.310 427.930 3208.490 ;
        RECT 475.510 3207.310 476.690 3208.490 ;
        RECT 523.350 3207.310 524.530 3208.490 ;
        RECT 678.830 3208.050 680.010 3208.490 ;
        RECT 682.510 3208.050 683.690 3208.490 ;
        RECT 678.830 3207.750 683.690 3208.050 ;
        RECT 678.830 3207.310 680.010 3207.750 ;
        RECT 682.510 3207.310 683.690 3207.750 ;
        RECT 765.310 3207.310 766.490 3208.490 ;
        RECT 812.230 3207.310 813.410 3208.490 ;
        RECT 820.510 3207.310 821.690 3208.490 ;
        RECT 893.190 3207.310 894.370 3208.490 ;
        RECT 930.910 3207.310 932.090 3208.490 ;
        RECT 978.750 3207.310 979.930 3208.490 ;
        RECT 1204.150 3207.310 1205.330 3208.490 ;
        RECT 1268.550 3207.310 1269.730 3208.490 ;
        RECT 1321.910 3207.310 1323.090 3208.490 ;
        RECT 1365.150 3207.310 1366.330 3208.490 ;
        RECT 1413.910 3207.310 1415.090 3208.490 ;
        RECT 1558.350 3207.310 1559.530 3208.490 ;
        RECT 1676.110 3207.310 1677.290 3208.490 ;
        RECT 1747.870 3207.310 1749.050 3208.490 ;
        RECT 1753.390 3207.310 1754.570 3208.490 ;
        RECT 1848.150 3207.310 1849.330 3208.490 ;
        RECT 1897.830 3207.310 1899.010 3208.490 ;
        RECT 1955.790 3207.310 1956.970 3208.490 ;
        RECT 1993.510 3207.310 1994.690 3208.490 ;
        RECT 2052.390 3207.310 2053.570 3208.490 ;
        RECT 2090.110 3207.310 2091.290 3208.490 ;
        RECT 2137.950 3207.310 2139.130 3208.490 ;
        RECT 2214.310 3207.310 2215.490 3208.490 ;
        RECT 2262.150 3207.310 2263.330 3208.490 ;
        RECT 2311.830 3207.310 2313.010 3208.490 ;
        RECT 2358.750 3207.310 2359.930 3208.490 ;
        RECT 2407.510 3207.310 2408.690 3208.490 ;
        RECT 2455.350 3207.310 2456.530 3208.490 ;
        RECT 2504.110 3207.310 2505.290 3208.490 ;
        RECT 2597.030 3207.310 2598.210 3208.490 ;
        RECT 2610.830 3207.310 2612.010 3208.490 ;
        RECT 2611.270 223.545 2611.570 3207.310 ;
        RECT 2611.255 223.215 2611.585 223.545 ;
        RECT 2656.335 203.495 2656.665 203.825 ;
        RECT 2656.350 202.465 2656.650 203.495 ;
        RECT 2656.335 202.135 2656.665 202.465 ;
        RECT 2752.935 200.095 2753.265 200.425 ;
        RECT 2752.950 199.065 2753.250 200.095 ;
        RECT 2752.935 198.735 2753.265 199.065 ;
      LAYER met5 ;
        RECT 253.580 3207.100 325.100 3208.700 ;
        RECT 323.500 3201.900 325.100 3207.100 ;
        RECT 337.300 3207.100 380.300 3208.700 ;
        RECT 337.300 3201.900 338.900 3207.100 ;
        RECT 323.500 3200.300 338.900 3201.900 ;
        RECT 426.540 3201.900 428.140 3208.700 ;
        RECT 433.900 3207.100 476.900 3208.700 ;
        RECT 433.900 3201.900 435.500 3207.100 ;
        RECT 426.540 3200.300 435.500 3201.900 ;
        RECT 523.140 3201.900 524.740 3208.700 ;
        RECT 530.500 3207.100 586.380 3208.700 ;
        RECT 530.500 3201.900 532.100 3207.100 ;
        RECT 584.780 3205.300 586.380 3207.100 ;
        RECT 627.100 3207.100 680.220 3208.700 ;
        RECT 682.300 3207.100 717.940 3208.700 ;
        RECT 584.780 3203.700 621.340 3205.300 ;
        RECT 523.140 3200.300 532.100 3201.900 ;
        RECT 619.740 3201.900 621.340 3203.700 ;
        RECT 627.100 3201.900 628.700 3207.100 ;
        RECT 619.740 3200.300 628.700 3201.900 ;
        RECT 716.340 3201.900 717.940 3207.100 ;
        RECT 723.700 3207.100 766.700 3208.700 ;
        RECT 812.020 3208.460 821.900 3210.060 ;
        RECT 812.020 3207.100 813.620 3208.460 ;
        RECT 820.300 3207.100 821.900 3208.460 ;
        RECT 892.980 3207.100 932.300 3208.700 ;
        RECT 723.700 3201.900 725.300 3207.100 ;
        RECT 978.540 3205.300 980.140 3208.700 ;
        RECT 1007.060 3207.100 1050.060 3208.700 ;
        RECT 978.540 3203.700 1001.300 3205.300 ;
        RECT 716.340 3200.300 725.300 3201.900 ;
        RECT 999.700 3201.900 1001.300 3203.700 ;
        RECT 1007.060 3201.900 1008.660 3207.100 ;
        RECT 999.700 3200.300 1008.660 3201.900 ;
        RECT 1048.460 3201.900 1050.060 3207.100 ;
        RECT 1063.180 3207.100 1104.340 3208.700 ;
        RECT 1063.180 3201.900 1064.780 3207.100 ;
        RECT 1048.460 3200.300 1064.780 3201.900 ;
        RECT 1102.740 3201.900 1104.340 3207.100 ;
        RECT 1134.020 3207.100 1205.540 3208.700 ;
        RECT 1268.340 3207.100 1323.300 3208.700 ;
        RECT 1364.940 3207.100 1415.300 3208.700 ;
        RECT 1134.020 3201.900 1135.620 3207.100 ;
        RECT 1268.340 3203.700 1270.860 3207.100 ;
        RECT 1364.940 3203.700 1367.460 3207.100 ;
        RECT 1558.140 3205.300 1559.740 3208.700 ;
        RECT 1593.100 3207.100 1629.660 3208.700 ;
        RECT 1558.140 3203.700 1580.900 3205.300 ;
        RECT 1102.740 3200.300 1135.620 3201.900 ;
        RECT 1579.300 3201.900 1580.900 3203.700 ;
        RECT 1593.100 3201.900 1594.700 3207.100 ;
        RECT 1628.060 3205.300 1629.660 3207.100 ;
        RECT 1675.900 3205.300 1677.500 3208.700 ;
        RECT 1628.060 3203.700 1677.500 3205.300 ;
        RECT 1747.660 3205.300 1749.260 3208.700 ;
        RECT 1752.260 3207.100 1754.780 3208.700 ;
        RECT 1847.940 3207.100 1899.220 3208.700 ;
        RECT 1955.580 3207.100 1994.900 3208.700 ;
        RECT 2052.180 3207.100 2091.500 3208.700 ;
        RECT 1752.260 3205.300 1753.860 3207.100 ;
        RECT 1747.660 3203.700 1753.860 3205.300 ;
        RECT 1847.940 3203.700 1850.460 3207.100 ;
        RECT 2137.740 3205.300 2139.340 3208.700 ;
        RECT 2172.700 3207.100 2215.700 3208.700 ;
        RECT 2137.740 3203.700 2160.500 3205.300 ;
        RECT 1579.300 3200.300 1594.700 3201.900 ;
        RECT 2158.900 3201.900 2160.500 3203.700 ;
        RECT 2172.700 3201.900 2174.300 3207.100 ;
        RECT 2158.900 3200.300 2174.300 3201.900 ;
        RECT 2261.940 3201.900 2263.540 3208.700 ;
        RECT 2269.300 3207.100 2313.220 3208.700 ;
        RECT 2269.300 3201.900 2270.900 3207.100 ;
        RECT 2261.940 3200.300 2270.900 3201.900 ;
        RECT 2358.540 3201.900 2360.140 3208.700 ;
        RECT 2365.900 3207.100 2408.900 3208.700 ;
        RECT 2365.900 3201.900 2367.500 3207.100 ;
        RECT 2358.540 3200.300 2367.500 3201.900 ;
        RECT 2455.140 3201.900 2456.740 3208.700 ;
        RECT 2462.500 3207.100 2505.500 3208.700 ;
        RECT 2596.820 3207.100 2612.220 3208.700 ;
        RECT 2462.500 3201.900 2464.100 3207.100 ;
        RECT 2455.140 3200.300 2464.100 3201.900 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 880.050 3220.720 880.370 3220.780 ;
        RECT 2621.610 3220.720 2621.930 3220.780 ;
        RECT 880.050 3220.580 2621.930 3220.720 ;
        RECT 880.050 3220.520 880.370 3220.580 ;
        RECT 2621.610 3220.520 2621.930 3220.580 ;
        RECT 2621.610 2552.960 2621.930 2553.020 ;
        RECT 2900.830 2552.960 2901.150 2553.020 ;
        RECT 2621.610 2552.820 2901.150 2552.960 ;
        RECT 2621.610 2552.760 2621.930 2552.820 ;
        RECT 2900.830 2552.760 2901.150 2552.820 ;
      LAYER via ;
        RECT 880.080 3220.520 880.340 3220.780 ;
        RECT 2621.640 3220.520 2621.900 3220.780 ;
        RECT 2621.640 2552.760 2621.900 2553.020 ;
        RECT 2900.860 2552.760 2901.120 2553.020 ;
      LAYER met2 ;
        RECT 880.080 3220.490 880.340 3220.810 ;
        RECT 2621.640 3220.490 2621.900 3220.810 ;
        RECT 880.140 3220.000 880.280 3220.490 ;
        RECT 880.120 3216.000 880.400 3220.000 ;
        RECT 2621.700 2553.050 2621.840 3220.490 ;
        RECT 2621.640 2552.730 2621.900 2553.050 ;
        RECT 2900.860 2552.730 2901.120 2553.050 ;
        RECT 2900.920 2551.885 2901.060 2552.730 ;
        RECT 2900.850 2551.515 2901.130 2551.885 ;
      LAYER via2 ;
        RECT 2900.850 2551.560 2901.130 2551.840 ;
      LAYER met3 ;
        RECT 2900.825 2551.850 2901.155 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.825 2551.550 2924.800 2551.850 ;
        RECT 2900.825 2551.535 2901.155 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 943.090 3232.875 943.370 3233.245 ;
        RECT 943.160 3220.000 943.300 3232.875 ;
        RECT 943.140 3216.000 943.420 3220.000 ;
      LAYER via2 ;
        RECT 943.090 3232.920 943.370 3233.200 ;
      LAYER met3 ;
        RECT 943.065 3233.210 943.395 3233.225 ;
        RECT 2602.950 3233.210 2603.330 3233.220 ;
        RECT 943.065 3232.910 2603.330 3233.210 ;
        RECT 943.065 3232.895 943.395 3232.910 ;
        RECT 2602.950 3232.900 2603.330 3232.910 ;
        RECT 2602.950 3208.730 2603.330 3208.740 ;
        RECT 2606.630 3208.730 2607.010 3208.740 ;
        RECT 2602.950 3208.430 2607.010 3208.730 ;
        RECT 2602.950 3208.420 2603.330 3208.430 ;
        RECT 2606.630 3208.420 2607.010 3208.430 ;
        RECT 2609.390 2816.060 2609.770 2816.380 ;
        RECT 2607.550 2813.650 2607.930 2813.660 ;
        RECT 2609.430 2813.650 2609.730 2816.060 ;
        RECT 2607.550 2813.350 2609.730 2813.650 ;
        RECT 2607.550 2813.340 2607.930 2813.350 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2916.710 2786.150 2924.800 2786.450 ;
        RECT 2607.550 2782.740 2607.930 2783.060 ;
        RECT 2607.590 2782.370 2607.890 2782.740 ;
        RECT 2607.590 2782.070 2642.850 2782.370 ;
        RECT 2642.550 2781.690 2642.850 2782.070 ;
        RECT 2691.310 2782.070 2739.450 2782.370 ;
        RECT 2642.550 2781.390 2690.690 2781.690 ;
        RECT 2690.390 2781.010 2690.690 2781.390 ;
        RECT 2691.310 2781.010 2691.610 2782.070 ;
        RECT 2739.150 2781.690 2739.450 2782.070 ;
        RECT 2787.910 2782.070 2836.050 2782.370 ;
        RECT 2739.150 2781.390 2787.290 2781.690 ;
        RECT 2690.390 2780.710 2691.610 2781.010 ;
        RECT 2786.990 2781.010 2787.290 2781.390 ;
        RECT 2787.910 2781.010 2788.210 2782.070 ;
        RECT 2835.750 2781.690 2836.050 2782.070 ;
        RECT 2835.750 2781.390 2883.890 2781.690 ;
        RECT 2786.990 2780.710 2788.210 2781.010 ;
        RECT 2883.590 2781.010 2883.890 2781.390 ;
        RECT 2916.710 2781.010 2917.010 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 2883.590 2780.710 2917.010 2781.010 ;
      LAYER via3 ;
        RECT 2602.980 3232.900 2603.300 3233.220 ;
        RECT 2602.980 3208.420 2603.300 3208.740 ;
        RECT 2606.660 3208.420 2606.980 3208.740 ;
        RECT 2609.420 2816.060 2609.740 2816.380 ;
        RECT 2607.580 2813.340 2607.900 2813.660 ;
        RECT 2607.580 2782.740 2607.900 2783.060 ;
      LAYER met4 ;
        RECT 2602.975 3232.895 2603.305 3233.225 ;
        RECT 2602.990 3208.745 2603.290 3232.895 ;
        RECT 2602.975 3208.415 2603.305 3208.745 ;
        RECT 2606.655 3208.415 2606.985 3208.745 ;
        RECT 2606.670 3034.650 2606.970 3208.415 ;
        RECT 2606.670 3034.350 2608.810 3034.650 ;
        RECT 2608.510 2956.450 2608.810 3034.350 ;
        RECT 2607.590 2956.150 2608.810 2956.450 ;
        RECT 2607.590 2915.650 2607.890 2956.150 ;
        RECT 2607.590 2915.350 2608.810 2915.650 ;
        RECT 2608.510 2874.850 2608.810 2915.350 ;
        RECT 2608.510 2874.550 2610.650 2874.850 ;
        RECT 2610.350 2851.050 2610.650 2874.550 ;
        RECT 2609.430 2850.750 2610.650 2851.050 ;
        RECT 2609.430 2816.385 2609.730 2850.750 ;
        RECT 2609.415 2816.055 2609.745 2816.385 ;
        RECT 2607.575 2813.650 2607.905 2813.665 ;
        RECT 2606.670 2813.350 2607.905 2813.650 ;
        RECT 2606.670 2783.050 2606.970 2813.350 ;
        RECT 2607.575 2813.335 2607.905 2813.350 ;
        RECT 2607.575 2783.050 2607.905 2783.065 ;
        RECT 2606.670 2782.750 2607.905 2783.050 ;
        RECT 2607.575 2782.735 2607.905 2782.750 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1006.570 3233.555 1006.850 3233.925 ;
        RECT 1006.640 3220.000 1006.780 3233.555 ;
        RECT 1006.620 3216.000 1006.900 3220.000 ;
        RECT 2610.590 3083.955 2610.870 3084.325 ;
        RECT 2610.660 3051.005 2610.800 3083.955 ;
        RECT 2610.590 3050.635 2610.870 3051.005 ;
        RECT 2622.550 3034.995 2622.830 3035.365 ;
        RECT 2622.620 3016.325 2622.760 3034.995 ;
        RECT 2622.550 3015.955 2622.830 3016.325 ;
      LAYER via2 ;
        RECT 1006.570 3233.600 1006.850 3233.880 ;
        RECT 2610.590 3084.000 2610.870 3084.280 ;
        RECT 2610.590 3050.680 2610.870 3050.960 ;
        RECT 2622.550 3035.040 2622.830 3035.320 ;
        RECT 2622.550 3016.000 2622.830 3016.280 ;
      LAYER met3 ;
        RECT 1006.545 3233.890 1006.875 3233.905 ;
        RECT 2607.550 3233.890 2607.930 3233.900 ;
        RECT 1006.545 3233.590 2607.930 3233.890 ;
        RECT 1006.545 3233.575 1006.875 3233.590 ;
        RECT 2607.550 3233.580 2607.930 3233.590 ;
        RECT 2607.550 3183.940 2607.930 3184.260 ;
        RECT 2607.590 3182.900 2607.890 3183.940 ;
        RECT 2607.550 3182.580 2607.930 3182.900 ;
        RECT 2607.550 3143.820 2607.930 3144.140 ;
        RECT 2607.590 3140.060 2607.890 3143.820 ;
        RECT 2607.550 3139.740 2607.930 3140.060 ;
        RECT 2607.550 3084.290 2607.930 3084.300 ;
        RECT 2610.565 3084.290 2610.895 3084.305 ;
        RECT 2607.550 3083.990 2610.895 3084.290 ;
        RECT 2607.550 3083.980 2607.930 3083.990 ;
        RECT 2610.565 3083.975 2610.895 3083.990 ;
        RECT 2607.550 3050.970 2607.930 3050.980 ;
        RECT 2610.565 3050.970 2610.895 3050.985 ;
        RECT 2607.550 3050.670 2610.895 3050.970 ;
        RECT 2607.550 3050.660 2607.930 3050.670 ;
        RECT 2610.565 3050.655 2610.895 3050.670 ;
        RECT 2607.550 3035.330 2607.930 3035.340 ;
        RECT 2622.525 3035.330 2622.855 3035.345 ;
        RECT 2607.550 3035.030 2622.855 3035.330 ;
        RECT 2607.550 3035.020 2607.930 3035.030 ;
        RECT 2622.525 3035.015 2622.855 3035.030 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2916.710 3020.750 2924.800 3021.050 ;
        RECT 2691.310 3016.670 2739.450 3016.970 ;
        RECT 2622.525 3016.290 2622.855 3016.305 ;
        RECT 2622.525 3015.990 2690.690 3016.290 ;
        RECT 2622.525 3015.975 2622.855 3015.990 ;
        RECT 2690.390 3015.610 2690.690 3015.990 ;
        RECT 2691.310 3015.610 2691.610 3016.670 ;
        RECT 2739.150 3016.290 2739.450 3016.670 ;
        RECT 2787.910 3016.670 2836.050 3016.970 ;
        RECT 2739.150 3015.990 2787.290 3016.290 ;
        RECT 2690.390 3015.310 2691.610 3015.610 ;
        RECT 2786.990 3015.610 2787.290 3015.990 ;
        RECT 2787.910 3015.610 2788.210 3016.670 ;
        RECT 2835.750 3016.290 2836.050 3016.670 ;
        RECT 2835.750 3015.990 2883.890 3016.290 ;
        RECT 2786.990 3015.310 2788.210 3015.610 ;
        RECT 2883.590 3015.610 2883.890 3015.990 ;
        RECT 2916.710 3015.610 2917.010 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 2883.590 3015.310 2917.010 3015.610 ;
      LAYER via3 ;
        RECT 2607.580 3233.580 2607.900 3233.900 ;
        RECT 2607.580 3183.940 2607.900 3184.260 ;
        RECT 2607.580 3182.580 2607.900 3182.900 ;
        RECT 2607.580 3143.820 2607.900 3144.140 ;
        RECT 2607.580 3139.740 2607.900 3140.060 ;
        RECT 2607.580 3083.980 2607.900 3084.300 ;
        RECT 2607.580 3050.660 2607.900 3050.980 ;
        RECT 2607.580 3035.020 2607.900 3035.340 ;
      LAYER met4 ;
        RECT 2607.575 3233.575 2607.905 3233.905 ;
        RECT 2607.590 3184.265 2607.890 3233.575 ;
        RECT 2607.575 3183.935 2607.905 3184.265 ;
        RECT 2607.575 3182.575 2607.905 3182.905 ;
        RECT 2607.590 3144.145 2607.890 3182.575 ;
        RECT 2607.575 3143.815 2607.905 3144.145 ;
        RECT 2607.575 3139.735 2607.905 3140.065 ;
        RECT 2607.590 3084.305 2607.890 3139.735 ;
        RECT 2607.575 3083.975 2607.905 3084.305 ;
        RECT 2607.575 3050.655 2607.905 3050.985 ;
        RECT 2607.590 3035.345 2607.890 3050.655 ;
        RECT 2607.575 3035.015 2607.905 3035.345 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1076.010 3250.300 1076.330 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 1076.010 3250.160 2901.150 3250.300 ;
        RECT 1076.010 3250.100 1076.330 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
      LAYER via ;
        RECT 1076.040 3250.100 1076.300 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 1076.040 3250.070 1076.300 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 1069.640 3218.850 1069.920 3220.000 ;
        RECT 1076.100 3218.850 1076.240 3250.070 ;
        RECT 1069.640 3218.710 1076.240 3218.850 ;
        RECT 1069.640 3216.000 1069.920 3218.710 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1138.110 3484.900 1138.430 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 1138.110 3484.760 2901.150 3484.900 ;
        RECT 1138.110 3484.700 1138.430 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 1138.140 3484.700 1138.400 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 1138.140 3484.670 1138.400 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 1138.200 3220.210 1138.340 3484.670 ;
        RECT 1134.980 3220.070 1138.340 3220.210 ;
        RECT 1132.660 3218.850 1132.940 3220.000 ;
        RECT 1134.980 3218.850 1135.120 3220.070 ;
        RECT 1132.660 3218.710 1135.120 3218.850 ;
        RECT 1132.660 3216.000 1132.940 3218.710 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1200.210 3502.580 1200.530 3502.640 ;
        RECT 2635.870 3502.580 2636.190 3502.640 ;
        RECT 1200.210 3502.440 2636.190 3502.580 ;
        RECT 1200.210 3502.380 1200.530 3502.440 ;
        RECT 2635.870 3502.380 2636.190 3502.440 ;
      LAYER via ;
        RECT 1200.240 3502.380 1200.500 3502.640 ;
        RECT 2635.900 3502.380 2636.160 3502.640 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3502.670 2636.100 3517.600 ;
        RECT 1200.240 3502.350 1200.500 3502.670 ;
        RECT 2635.900 3502.350 2636.160 3502.670 ;
        RECT 1196.140 3218.850 1196.420 3220.000 ;
        RECT 1200.300 3218.850 1200.440 3502.350 ;
        RECT 1196.140 3218.710 1200.440 3218.850 ;
        RECT 1196.140 3216.000 1196.420 3218.710 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1262.310 3504.280 1262.630 3504.340 ;
        RECT 2311.570 3504.280 2311.890 3504.340 ;
        RECT 1262.310 3504.140 2311.890 3504.280 ;
        RECT 1262.310 3504.080 1262.630 3504.140 ;
        RECT 2311.570 3504.080 2311.890 3504.140 ;
      LAYER via ;
        RECT 1262.340 3504.080 1262.600 3504.340 ;
        RECT 2311.600 3504.080 2311.860 3504.340 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3504.370 2311.800 3517.600 ;
        RECT 1262.340 3504.050 1262.600 3504.370 ;
        RECT 2311.600 3504.050 2311.860 3504.370 ;
        RECT 1259.160 3218.850 1259.440 3220.000 ;
        RECT 1262.400 3218.850 1262.540 3504.050 ;
        RECT 1259.160 3218.710 1262.540 3218.850 ;
        RECT 1259.160 3216.000 1259.440 3218.710 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1324.410 3500.540 1324.730 3500.600 ;
        RECT 1987.270 3500.540 1987.590 3500.600 ;
        RECT 1324.410 3500.400 1987.590 3500.540 ;
        RECT 1324.410 3500.340 1324.730 3500.400 ;
        RECT 1987.270 3500.340 1987.590 3500.400 ;
      LAYER via ;
        RECT 1324.440 3500.340 1324.700 3500.600 ;
        RECT 1987.300 3500.340 1987.560 3500.600 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3500.630 1987.500 3517.600 ;
        RECT 1324.440 3500.310 1324.700 3500.630 ;
        RECT 1987.300 3500.310 1987.560 3500.630 ;
        RECT 1322.180 3218.850 1322.460 3220.000 ;
        RECT 1324.500 3218.850 1324.640 3500.310 ;
        RECT 1322.180 3218.710 1324.640 3218.850 ;
        RECT 1322.180 3216.000 1322.460 3218.710 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1386.510 3499.180 1386.830 3499.240 ;
        RECT 1662.510 3499.180 1662.830 3499.240 ;
        RECT 1386.510 3499.040 1662.830 3499.180 ;
        RECT 1386.510 3498.980 1386.830 3499.040 ;
        RECT 1662.510 3498.980 1662.830 3499.040 ;
      LAYER via ;
        RECT 1386.540 3498.980 1386.800 3499.240 ;
        RECT 1662.540 3498.980 1662.800 3499.240 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3499.270 1662.740 3517.600 ;
        RECT 1386.540 3498.950 1386.800 3499.270 ;
        RECT 1662.540 3498.950 1662.800 3499.270 ;
        RECT 1385.200 3219.530 1385.480 3220.000 ;
        RECT 1386.600 3219.530 1386.740 3498.950 ;
        RECT 1385.200 3219.390 1386.740 3219.530 ;
        RECT 1385.200 3216.000 1385.480 3219.390 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3498.840 1338.530 3498.900 ;
        RECT 1442.170 3498.840 1442.490 3498.900 ;
        RECT 1338.210 3498.700 1442.490 3498.840 ;
        RECT 1338.210 3498.640 1338.530 3498.700 ;
        RECT 1442.170 3498.640 1442.490 3498.700 ;
      LAYER via ;
        RECT 1338.240 3498.640 1338.500 3498.900 ;
        RECT 1442.200 3498.640 1442.460 3498.900 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3498.930 1338.440 3517.600 ;
        RECT 1338.240 3498.610 1338.500 3498.930 ;
        RECT 1442.200 3498.610 1442.460 3498.930 ;
        RECT 1442.260 3220.210 1442.400 3498.610 ;
        RECT 1442.260 3220.070 1446.540 3220.210 ;
        RECT 1446.400 3218.850 1446.540 3220.070 ;
        RECT 1448.680 3218.850 1448.960 3220.000 ;
        RECT 1446.400 3218.710 1448.960 3218.850 ;
        RECT 1448.680 3216.000 1448.960 3218.710 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2766.510 435.780 2766.830 435.840 ;
        RECT 2801.010 435.780 2801.330 435.840 ;
        RECT 2766.510 435.640 2801.330 435.780 ;
        RECT 2766.510 435.580 2766.830 435.640 ;
        RECT 2801.010 435.580 2801.330 435.640 ;
      LAYER via ;
        RECT 2766.540 435.580 2766.800 435.840 ;
        RECT 2801.040 435.580 2801.300 435.840 ;
      LAYER met2 ;
        RECT 311.970 3230.835 312.250 3231.205 ;
        RECT 312.040 3220.000 312.180 3230.835 ;
        RECT 312.020 3216.000 312.300 3220.000 ;
        RECT 2745.830 436.715 2746.110 437.085 ;
        RECT 2669.930 436.035 2670.210 436.405 ;
        RECT 2670.000 435.610 2670.140 436.035 ;
        RECT 2670.850 435.610 2671.130 435.725 ;
        RECT 2670.000 435.470 2671.130 435.610 ;
        RECT 2670.850 435.355 2671.130 435.470 ;
        RECT 2745.900 435.045 2746.040 436.715 ;
        RECT 2801.030 436.035 2801.310 436.405 ;
        RECT 2801.100 435.870 2801.240 436.035 ;
        RECT 2766.540 435.725 2766.800 435.870 ;
        RECT 2766.530 435.355 2766.810 435.725 ;
        RECT 2801.040 435.550 2801.300 435.870 ;
        RECT 2745.830 434.675 2746.110 435.045 ;
      LAYER via2 ;
        RECT 311.970 3230.880 312.250 3231.160 ;
        RECT 2745.830 436.760 2746.110 437.040 ;
        RECT 2669.930 436.080 2670.210 436.360 ;
        RECT 2670.850 435.400 2671.130 435.680 ;
        RECT 2801.030 436.080 2801.310 436.360 ;
        RECT 2766.530 435.400 2766.810 435.680 ;
        RECT 2745.830 434.720 2746.110 435.000 ;
      LAYER met3 ;
        RECT 311.945 3231.170 312.275 3231.185 ;
        RECT 2603.870 3231.170 2604.250 3231.180 ;
        RECT 311.945 3230.870 2604.250 3231.170 ;
        RECT 311.945 3230.855 312.275 3230.870 ;
        RECT 2603.870 3230.860 2604.250 3230.870 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2916.710 439.470 2924.800 439.770 ;
        RECT 2697.710 437.050 2698.090 437.060 ;
        RECT 2745.805 437.050 2746.135 437.065 ;
        RECT 2697.710 436.750 2746.135 437.050 ;
        RECT 2697.710 436.740 2698.090 436.750 ;
        RECT 2745.805 436.735 2746.135 436.750 ;
        RECT 2669.905 436.370 2670.235 436.385 ;
        RECT 2622.310 436.070 2670.235 436.370 ;
        RECT 2607.550 435.010 2607.930 435.020 ;
        RECT 2622.310 435.010 2622.610 436.070 ;
        RECT 2669.905 436.055 2670.235 436.070 ;
        RECT 2801.005 436.370 2801.335 436.385 ;
        RECT 2801.005 436.070 2836.050 436.370 ;
        RECT 2801.005 436.055 2801.335 436.070 ;
        RECT 2670.825 435.690 2671.155 435.705 ;
        RECT 2697.710 435.690 2698.090 435.700 ;
        RECT 2766.505 435.690 2766.835 435.705 ;
        RECT 2670.825 435.390 2698.090 435.690 ;
        RECT 2670.825 435.375 2671.155 435.390 ;
        RECT 2697.710 435.380 2698.090 435.390 ;
        RECT 2752.950 435.390 2766.835 435.690 ;
        RECT 2835.750 435.690 2836.050 436.070 ;
        RECT 2916.710 435.690 2917.010 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
        RECT 2835.750 435.390 2883.890 435.690 ;
        RECT 2607.550 434.710 2622.610 435.010 ;
        RECT 2745.805 435.010 2746.135 435.025 ;
        RECT 2752.950 435.010 2753.250 435.390 ;
        RECT 2766.505 435.375 2766.835 435.390 ;
        RECT 2745.805 434.710 2753.250 435.010 ;
        RECT 2883.590 435.010 2883.890 435.390 ;
        RECT 2884.510 435.390 2917.010 435.690 ;
        RECT 2884.510 435.010 2884.810 435.390 ;
        RECT 2883.590 434.710 2884.810 435.010 ;
        RECT 2607.550 434.700 2607.930 434.710 ;
        RECT 2745.805 434.695 2746.135 434.710 ;
      LAYER via3 ;
        RECT 2603.900 3230.860 2604.220 3231.180 ;
        RECT 2697.740 436.740 2698.060 437.060 ;
        RECT 2607.580 434.700 2607.900 435.020 ;
        RECT 2697.740 435.380 2698.060 435.700 ;
      LAYER met4 ;
        RECT 2603.895 3230.855 2604.225 3231.185 ;
        RECT 2603.910 3058.450 2604.210 3230.855 ;
        RECT 2601.150 3058.150 2604.210 3058.450 ;
        RECT 2601.150 3051.650 2601.450 3058.150 ;
        RECT 2601.150 3051.350 2604.210 3051.650 ;
        RECT 2603.910 443.850 2604.210 3051.350 ;
        RECT 2603.910 443.550 2606.970 443.850 ;
        RECT 2606.670 433.650 2606.970 443.550 ;
        RECT 2697.735 436.735 2698.065 437.065 ;
        RECT 2697.750 435.705 2698.050 436.735 ;
        RECT 2697.735 435.375 2698.065 435.705 ;
        RECT 2607.575 434.695 2607.905 435.025 ;
        RECT 2607.590 433.650 2607.890 434.695 ;
        RECT 2606.670 433.350 2607.890 433.650 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3500.200 1014.230 3500.260 ;
        RECT 1511.170 3500.200 1511.490 3500.260 ;
        RECT 1013.910 3500.060 1511.490 3500.200 ;
        RECT 1013.910 3500.000 1014.230 3500.060 ;
        RECT 1511.170 3500.000 1511.490 3500.060 ;
      LAYER via ;
        RECT 1013.940 3500.000 1014.200 3500.260 ;
        RECT 1511.200 3500.000 1511.460 3500.260 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3500.290 1014.140 3517.600 ;
        RECT 1013.940 3499.970 1014.200 3500.290 ;
        RECT 1511.200 3499.970 1511.460 3500.290 ;
        RECT 1511.260 3219.530 1511.400 3499.970 ;
        RECT 1511.700 3219.530 1511.980 3220.000 ;
        RECT 1511.260 3219.390 1511.980 3219.530 ;
        RECT 1511.700 3216.000 1511.980 3219.390 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3504.620 689.470 3504.680 ;
        RECT 1573.270 3504.620 1573.590 3504.680 ;
        RECT 689.150 3504.480 1573.590 3504.620 ;
        RECT 689.150 3504.420 689.470 3504.480 ;
        RECT 1573.270 3504.420 1573.590 3504.480 ;
      LAYER via ;
        RECT 689.180 3504.420 689.440 3504.680 ;
        RECT 1573.300 3504.420 1573.560 3504.680 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3504.710 689.380 3517.600 ;
        RECT 689.180 3504.390 689.440 3504.710 ;
        RECT 1573.300 3504.390 1573.560 3504.710 ;
        RECT 1573.360 3219.530 1573.500 3504.390 ;
        RECT 1574.720 3219.530 1575.000 3220.000 ;
        RECT 1573.360 3219.390 1575.000 3219.530 ;
        RECT 1574.720 3216.000 1575.000 3219.390 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 3502.920 365.170 3502.980 ;
        RECT 1635.370 3502.920 1635.690 3502.980 ;
        RECT 364.850 3502.780 1635.690 3502.920 ;
        RECT 364.850 3502.720 365.170 3502.780 ;
        RECT 1635.370 3502.720 1635.690 3502.780 ;
      LAYER via ;
        RECT 364.880 3502.720 365.140 3502.980 ;
        RECT 1635.400 3502.720 1635.660 3502.980 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3503.010 365.080 3517.600 ;
        RECT 364.880 3502.690 365.140 3503.010 ;
        RECT 1635.400 3502.690 1635.660 3503.010 ;
        RECT 1635.460 3218.850 1635.600 3502.690 ;
        RECT 1638.200 3218.850 1638.480 3220.000 ;
        RECT 1635.460 3218.710 1638.480 3218.850 ;
        RECT 1638.200 3216.000 1638.480 3218.710 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.845 40.780 3517.600 ;
        RECT 40.570 3501.475 40.850 3501.845 ;
        RECT 1697.490 3501.475 1697.770 3501.845 ;
        RECT 1697.560 3218.850 1697.700 3501.475 ;
        RECT 1701.220 3218.850 1701.500 3220.000 ;
        RECT 1697.560 3218.710 1701.500 3218.850 ;
        RECT 1701.220 3216.000 1701.500 3218.710 ;
      LAYER via2 ;
        RECT 40.570 3501.520 40.850 3501.800 ;
        RECT 1697.490 3501.520 1697.770 3501.800 ;
      LAYER met3 ;
        RECT 40.545 3501.810 40.875 3501.825 ;
        RECT 1697.465 3501.810 1697.795 3501.825 ;
        RECT 40.545 3501.510 1697.795 3501.810 ;
        RECT 40.545 3501.495 40.875 3501.510 ;
        RECT 1697.465 3501.495 1697.795 3501.510 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 1759.570 3263.900 1759.890 3263.960 ;
        RECT 15.250 3263.760 1759.890 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 1759.570 3263.700 1759.890 3263.760 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 1759.600 3263.700 1759.860 3263.960 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 1759.600 3263.670 1759.860 3263.990 ;
        RECT 1759.660 3218.850 1759.800 3263.670 ;
        RECT 1764.240 3218.850 1764.520 3220.000 ;
        RECT 1759.660 3218.710 1764.520 3218.850 ;
        RECT 1764.240 3216.000 1764.520 3218.710 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.850 3235.000 20.170 3235.060 ;
        RECT 1827.650 3235.000 1827.970 3235.060 ;
        RECT 19.850 3234.860 1827.970 3235.000 ;
        RECT 19.850 3234.800 20.170 3234.860 ;
        RECT 1827.650 3234.800 1827.970 3234.860 ;
      LAYER via ;
        RECT 19.880 3234.800 20.140 3235.060 ;
        RECT 1827.680 3234.800 1827.940 3235.060 ;
      LAYER met2 ;
        RECT 19.880 3234.770 20.140 3235.090 ;
        RECT 1827.680 3234.770 1827.940 3235.090 ;
        RECT 19.940 2980.285 20.080 3234.770 ;
        RECT 1827.740 3220.000 1827.880 3234.770 ;
        RECT 1827.720 3216.000 1828.000 3220.000 ;
        RECT 19.870 2979.915 20.150 2980.285 ;
      LAYER via2 ;
        RECT 19.870 2979.960 20.150 2980.240 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 19.845 2980.250 20.175 2980.265 ;
        RECT -4.800 2979.950 20.175 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 19.845 2979.935 20.175 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 127.950 3228.540 128.270 3228.600 ;
        RECT 1890.670 3228.540 1890.990 3228.600 ;
        RECT 127.950 3228.400 1890.990 3228.540 ;
        RECT 127.950 3228.340 128.270 3228.400 ;
        RECT 1890.670 3228.340 1890.990 3228.400 ;
        RECT 15.250 2697.800 15.570 2697.860 ;
        RECT 127.950 2697.800 128.270 2697.860 ;
        RECT 15.250 2697.660 128.270 2697.800 ;
        RECT 15.250 2697.600 15.570 2697.660 ;
        RECT 127.950 2697.600 128.270 2697.660 ;
      LAYER via ;
        RECT 127.980 3228.340 128.240 3228.600 ;
        RECT 1890.700 3228.340 1890.960 3228.600 ;
        RECT 15.280 2697.600 15.540 2697.860 ;
        RECT 127.980 2697.600 128.240 2697.860 ;
      LAYER met2 ;
        RECT 127.980 3228.310 128.240 3228.630 ;
        RECT 1890.700 3228.310 1890.960 3228.630 ;
        RECT 128.040 2697.890 128.180 3228.310 ;
        RECT 1890.760 3220.000 1890.900 3228.310 ;
        RECT 1890.740 3216.000 1891.020 3220.000 ;
        RECT 15.280 2697.570 15.540 2697.890 ;
        RECT 127.980 2697.570 128.240 2697.890 ;
        RECT 15.340 2693.325 15.480 2697.570 ;
        RECT 15.270 2692.955 15.550 2693.325 ;
      LAYER via2 ;
        RECT 15.270 2693.000 15.550 2693.280 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 15.245 2693.290 15.575 2693.305 ;
        RECT -4.800 2692.990 15.575 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 15.245 2692.975 15.575 2692.990 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2405.740 16.950 2405.800 ;
        RECT 47.450 2405.740 47.770 2405.800 ;
        RECT 16.630 2405.600 47.770 2405.740 ;
        RECT 16.630 2405.540 16.950 2405.600 ;
        RECT 47.450 2405.540 47.770 2405.600 ;
      LAYER via ;
        RECT 16.660 2405.540 16.920 2405.800 ;
        RECT 47.480 2405.540 47.740 2405.800 ;
      LAYER met2 ;
        RECT 1952.790 3216.810 1953.070 3216.925 ;
        RECT 1953.760 3216.810 1954.040 3220.000 ;
        RECT 1952.790 3216.670 1954.040 3216.810 ;
        RECT 1952.790 3216.555 1953.070 3216.670 ;
        RECT 1953.760 3216.000 1954.040 3216.670 ;
        RECT 47.470 3211.115 47.750 3211.485 ;
        RECT 47.540 2405.830 47.680 3211.115 ;
        RECT 16.660 2405.685 16.920 2405.830 ;
        RECT 16.650 2405.315 16.930 2405.685 ;
        RECT 47.480 2405.510 47.740 2405.830 ;
      LAYER via2 ;
        RECT 1952.790 3216.600 1953.070 3216.880 ;
        RECT 47.470 3211.160 47.750 3211.440 ;
        RECT 16.650 2405.360 16.930 2405.640 ;
      LAYER met3 ;
        RECT 1952.765 3216.900 1953.095 3216.905 ;
        RECT 1952.510 3216.890 1953.095 3216.900 ;
        RECT 1952.310 3216.590 1953.095 3216.890 ;
        RECT 1952.510 3216.580 1953.095 3216.590 ;
        RECT 1952.765 3216.575 1953.095 3216.580 ;
        RECT 47.445 3211.450 47.775 3211.465 ;
        RECT 1952.510 3211.450 1952.890 3211.460 ;
        RECT 47.445 3211.150 1952.890 3211.450 ;
        RECT 47.445 3211.135 47.775 3211.150 ;
        RECT 1952.510 3211.140 1952.890 3211.150 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 16.625 2405.650 16.955 2405.665 ;
        RECT -4.800 2405.350 16.955 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 16.625 2405.335 16.955 2405.350 ;
      LAYER via3 ;
        RECT 1952.540 3216.580 1952.860 3216.900 ;
        RECT 1952.540 3211.140 1952.860 3211.460 ;
      LAYER met4 ;
        RECT 1952.535 3216.575 1952.865 3216.905 ;
        RECT 1952.550 3211.465 1952.850 3216.575 ;
        RECT 1952.535 3211.135 1952.865 3211.465 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 46.990 3219.020 47.310 3219.080 ;
        RECT 2014.870 3219.020 2015.190 3219.080 ;
        RECT 46.990 3218.880 2015.190 3219.020 ;
        RECT 46.990 3218.820 47.310 3218.880 ;
        RECT 2014.870 3218.820 2015.190 3218.880 ;
        RECT 16.630 2120.480 16.950 2120.540 ;
        RECT 46.990 2120.480 47.310 2120.540 ;
        RECT 16.630 2120.340 47.310 2120.480 ;
        RECT 16.630 2120.280 16.950 2120.340 ;
        RECT 46.990 2120.280 47.310 2120.340 ;
      LAYER via ;
        RECT 47.020 3218.820 47.280 3219.080 ;
        RECT 2014.900 3218.820 2015.160 3219.080 ;
        RECT 16.660 2120.280 16.920 2120.540 ;
        RECT 47.020 2120.280 47.280 2120.540 ;
      LAYER met2 ;
        RECT 47.020 3218.790 47.280 3219.110 ;
        RECT 2014.900 3218.850 2015.160 3219.110 ;
        RECT 2016.780 3218.850 2017.060 3220.000 ;
        RECT 2014.900 3218.790 2017.060 3218.850 ;
        RECT 47.080 2120.570 47.220 3218.790 ;
        RECT 2014.960 3218.710 2017.060 3218.790 ;
        RECT 2016.780 3216.000 2017.060 3218.710 ;
        RECT 16.660 2120.250 16.920 2120.570 ;
        RECT 47.020 2120.250 47.280 2120.570 ;
        RECT 16.720 2118.725 16.860 2120.250 ;
        RECT 16.650 2118.355 16.930 2118.725 ;
      LAYER via2 ;
        RECT 16.650 2118.400 16.930 2118.680 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.625 2118.690 16.955 2118.705 ;
        RECT -4.800 2118.390 16.955 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.625 2118.375 16.955 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 203.390 3227.860 203.710 3227.920 ;
        RECT 2080.190 3227.860 2080.510 3227.920 ;
        RECT 203.390 3227.720 2080.510 3227.860 ;
        RECT 203.390 3227.660 203.710 3227.720 ;
        RECT 2080.190 3227.660 2080.510 3227.720 ;
        RECT 15.710 1835.220 16.030 1835.280 ;
        RECT 203.390 1835.220 203.710 1835.280 ;
        RECT 15.710 1835.080 203.710 1835.220 ;
        RECT 15.710 1835.020 16.030 1835.080 ;
        RECT 203.390 1835.020 203.710 1835.080 ;
      LAYER via ;
        RECT 203.420 3227.660 203.680 3227.920 ;
        RECT 2080.220 3227.660 2080.480 3227.920 ;
        RECT 15.740 1835.020 16.000 1835.280 ;
        RECT 203.420 1835.020 203.680 1835.280 ;
      LAYER met2 ;
        RECT 203.420 3227.630 203.680 3227.950 ;
        RECT 2080.220 3227.630 2080.480 3227.950 ;
        RECT 203.480 1835.310 203.620 3227.630 ;
        RECT 2080.280 3220.000 2080.420 3227.630 ;
        RECT 2080.260 3216.000 2080.540 3220.000 ;
        RECT 15.740 1834.990 16.000 1835.310 ;
        RECT 203.420 1834.990 203.680 1835.310 ;
        RECT 15.800 1831.085 15.940 1834.990 ;
        RECT 15.730 1830.715 16.010 1831.085 ;
      LAYER via2 ;
        RECT 15.730 1830.760 16.010 1831.040 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 15.705 1831.050 16.035 1831.065 ;
        RECT -4.800 1830.750 16.035 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 15.705 1830.735 16.035 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 676.160 2618.710 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 2618.390 676.020 2901.150 676.160 ;
        RECT 2618.390 675.960 2618.710 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 2618.420 675.960 2618.680 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 375.040 3216.810 375.320 3220.000 ;
        RECT 376.370 3216.810 376.650 3216.925 ;
        RECT 375.040 3216.670 376.650 3216.810 ;
        RECT 375.040 3216.000 375.320 3216.670 ;
        RECT 376.370 3216.555 376.650 3216.670 ;
        RECT 2618.410 3213.155 2618.690 3213.525 ;
        RECT 2618.480 676.250 2618.620 3213.155 ;
        RECT 2618.420 675.930 2618.680 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 376.370 3216.600 376.650 3216.880 ;
        RECT 2618.410 3213.200 2618.690 3213.480 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 376.345 3216.900 376.675 3216.905 ;
        RECT 376.345 3216.890 376.930 3216.900 ;
        RECT 376.345 3216.590 377.130 3216.890 ;
        RECT 376.345 3216.580 376.930 3216.590 ;
        RECT 376.345 3216.575 376.675 3216.580 ;
        RECT 376.550 3213.490 376.930 3213.500 ;
        RECT 2618.385 3213.490 2618.715 3213.505 ;
        RECT 376.550 3213.190 2618.715 3213.490 ;
        RECT 376.550 3213.180 376.930 3213.190 ;
        RECT 2618.385 3213.175 2618.715 3213.190 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
      LAYER via3 ;
        RECT 376.580 3216.580 376.900 3216.900 ;
        RECT 376.580 3213.180 376.900 3213.500 ;
      LAYER met4 ;
        RECT 376.575 3216.575 376.905 3216.905 ;
        RECT 376.590 3213.505 376.890 3216.575 ;
        RECT 376.575 3213.175 376.905 3213.505 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 1544.180 16.950 1544.240 ;
        RECT 46.530 1544.180 46.850 1544.240 ;
        RECT 16.630 1544.040 46.850 1544.180 ;
        RECT 16.630 1543.980 16.950 1544.040 ;
        RECT 46.530 1543.980 46.850 1544.040 ;
      LAYER via ;
        RECT 16.660 1543.980 16.920 1544.240 ;
        RECT 46.560 1543.980 46.820 1544.240 ;
      LAYER met2 ;
        RECT 2142.310 3216.810 2142.590 3216.925 ;
        RECT 2143.280 3216.810 2143.560 3220.000 ;
        RECT 2142.310 3216.670 2143.560 3216.810 ;
        RECT 2142.310 3216.555 2142.590 3216.670 ;
        RECT 2143.280 3216.000 2143.560 3216.670 ;
        RECT 46.550 3214.515 46.830 3214.885 ;
        RECT 46.620 1544.270 46.760 3214.515 ;
        RECT 16.660 1544.125 16.920 1544.270 ;
        RECT 16.650 1543.755 16.930 1544.125 ;
        RECT 46.560 1543.950 46.820 1544.270 ;
      LAYER via2 ;
        RECT 2142.310 3216.600 2142.590 3216.880 ;
        RECT 46.550 3214.560 46.830 3214.840 ;
        RECT 16.650 1543.800 16.930 1544.080 ;
      LAYER met3 ;
        RECT 2142.285 3216.890 2142.615 3216.905 ;
        RECT 2142.070 3216.575 2142.615 3216.890 ;
        RECT 46.525 3214.850 46.855 3214.865 ;
        RECT 2142.070 3214.850 2142.370 3216.575 ;
        RECT 46.525 3214.550 2142.370 3214.850 ;
        RECT 46.525 3214.535 46.855 3214.550 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 16.625 1544.090 16.955 1544.105 ;
        RECT -4.800 1543.790 16.955 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 16.625 1543.775 16.955 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 24.910 3232.280 25.230 3232.340 ;
        RECT 2206.230 3232.280 2206.550 3232.340 ;
        RECT 24.910 3232.140 2206.550 3232.280 ;
        RECT 24.910 3232.080 25.230 3232.140 ;
        RECT 2206.230 3232.080 2206.550 3232.140 ;
        RECT 13.870 1331.000 14.190 1331.060 ;
        RECT 24.910 1331.000 25.230 1331.060 ;
        RECT 13.870 1330.860 25.230 1331.000 ;
        RECT 13.870 1330.800 14.190 1330.860 ;
        RECT 24.910 1330.800 25.230 1330.860 ;
      LAYER via ;
        RECT 24.940 3232.080 25.200 3232.340 ;
        RECT 2206.260 3232.080 2206.520 3232.340 ;
        RECT 13.900 1330.800 14.160 1331.060 ;
        RECT 24.940 1330.800 25.200 1331.060 ;
      LAYER met2 ;
        RECT 24.940 3232.050 25.200 3232.370 ;
        RECT 2206.260 3232.050 2206.520 3232.370 ;
        RECT 25.000 1331.090 25.140 3232.050 ;
        RECT 2206.320 3220.000 2206.460 3232.050 ;
        RECT 2206.300 3216.000 2206.580 3220.000 ;
        RECT 13.900 1330.770 14.160 1331.090 ;
        RECT 24.940 1330.770 25.200 1331.090 ;
        RECT 13.960 1328.565 14.100 1330.770 ;
        RECT 13.890 1328.195 14.170 1328.565 ;
      LAYER via2 ;
        RECT 13.890 1328.240 14.170 1328.520 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 13.865 1328.530 14.195 1328.545 ;
        RECT -4.800 1328.230 14.195 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 13.865 1328.215 14.195 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2268.350 3216.810 2268.630 3216.925 ;
        RECT 2269.780 3216.810 2270.060 3220.000 ;
        RECT 2268.350 3216.670 2270.060 3216.810 ;
        RECT 2268.350 3216.555 2268.630 3216.670 ;
        RECT 2269.780 3216.000 2270.060 3216.670 ;
        RECT 18.490 3212.475 18.770 3212.845 ;
        RECT 18.560 1113.005 18.700 3212.475 ;
        RECT 18.490 1112.635 18.770 1113.005 ;
      LAYER via2 ;
        RECT 2268.350 3216.600 2268.630 3216.880 ;
        RECT 18.490 3212.520 18.770 3212.800 ;
        RECT 18.490 1112.680 18.770 1112.960 ;
      LAYER met3 ;
        RECT 2268.325 3216.900 2268.655 3216.905 ;
        RECT 2268.070 3216.890 2268.655 3216.900 ;
        RECT 2267.870 3216.590 2268.655 3216.890 ;
        RECT 2268.070 3216.580 2268.655 3216.590 ;
        RECT 2268.325 3216.575 2268.655 3216.580 ;
        RECT 18.465 3212.810 18.795 3212.825 ;
        RECT 2268.070 3212.810 2268.450 3212.820 ;
        RECT 18.465 3212.510 2268.450 3212.810 ;
        RECT 18.465 3212.495 18.795 3212.510 ;
        RECT 2268.070 3212.500 2268.450 3212.510 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 18.465 1112.970 18.795 1112.985 ;
        RECT -4.800 1112.670 18.795 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 18.465 1112.655 18.795 1112.670 ;
      LAYER via3 ;
        RECT 2268.100 3216.580 2268.420 3216.900 ;
        RECT 2268.100 3212.500 2268.420 3212.820 ;
      LAYER met4 ;
        RECT 2268.095 3216.575 2268.425 3216.905 ;
        RECT 2268.110 3212.825 2268.410 3216.575 ;
        RECT 2268.095 3212.495 2268.425 3212.825 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 24.450 3231.260 24.770 3231.320 ;
        RECT 2332.730 3231.260 2333.050 3231.320 ;
        RECT 24.450 3231.120 2333.050 3231.260 ;
        RECT 24.450 3231.060 24.770 3231.120 ;
        RECT 2332.730 3231.060 2333.050 3231.120 ;
        RECT 13.870 897.500 14.190 897.560 ;
        RECT 24.450 897.500 24.770 897.560 ;
        RECT 13.870 897.360 24.770 897.500 ;
        RECT 13.870 897.300 14.190 897.360 ;
        RECT 24.450 897.300 24.770 897.360 ;
      LAYER via ;
        RECT 24.480 3231.060 24.740 3231.320 ;
        RECT 2332.760 3231.060 2333.020 3231.320 ;
        RECT 13.900 897.300 14.160 897.560 ;
        RECT 24.480 897.300 24.740 897.560 ;
      LAYER met2 ;
        RECT 24.480 3231.030 24.740 3231.350 ;
        RECT 2332.760 3231.030 2333.020 3231.350 ;
        RECT 24.540 897.590 24.680 3231.030 ;
        RECT 2332.820 3220.000 2332.960 3231.030 ;
        RECT 2332.800 3216.000 2333.080 3220.000 ;
        RECT 13.900 897.445 14.160 897.590 ;
        RECT 13.890 897.075 14.170 897.445 ;
        RECT 24.480 897.270 24.740 897.590 ;
      LAYER via2 ;
        RECT 13.890 897.120 14.170 897.400 ;
      LAYER met3 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 13.865 897.410 14.195 897.425 ;
        RECT -4.800 897.110 14.195 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 13.865 897.095 14.195 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2395.770 3229.475 2396.050 3229.845 ;
        RECT 2395.840 3220.000 2395.980 3229.475 ;
        RECT 2395.820 3216.000 2396.100 3220.000 ;
        RECT 17.570 3211.795 17.850 3212.165 ;
        RECT 17.640 681.885 17.780 3211.795 ;
        RECT 17.570 681.515 17.850 681.885 ;
      LAYER via2 ;
        RECT 2395.770 3229.520 2396.050 3229.800 ;
        RECT 17.570 3211.840 17.850 3212.120 ;
        RECT 17.570 681.560 17.850 681.840 ;
      LAYER met3 ;
        RECT 2356.390 3229.810 2356.770 3229.820 ;
        RECT 2395.745 3229.810 2396.075 3229.825 ;
        RECT 2356.390 3229.510 2396.075 3229.810 ;
        RECT 2356.390 3229.500 2356.770 3229.510 ;
        RECT 2395.745 3229.495 2396.075 3229.510 ;
        RECT 17.545 3212.130 17.875 3212.145 ;
        RECT 2356.390 3212.130 2356.770 3212.140 ;
        RECT 17.545 3211.830 2356.770 3212.130 ;
        RECT 17.545 3211.815 17.875 3211.830 ;
        RECT 2356.390 3211.820 2356.770 3211.830 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 17.545 681.850 17.875 681.865 ;
        RECT -4.800 681.550 17.875 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 17.545 681.535 17.875 681.550 ;
      LAYER via3 ;
        RECT 2356.420 3229.500 2356.740 3229.820 ;
        RECT 2356.420 3211.820 2356.740 3212.140 ;
      LAYER met4 ;
        RECT 2356.415 3229.495 2356.745 3229.825 ;
        RECT 2356.430 3212.145 2356.730 3229.495 ;
        RECT 2356.415 3211.815 2356.745 3212.145 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 23.990 3229.900 24.310 3229.960 ;
        RECT 2458.770 3229.900 2459.090 3229.960 ;
        RECT 23.990 3229.760 2459.090 3229.900 ;
        RECT 23.990 3229.700 24.310 3229.760 ;
        RECT 2458.770 3229.700 2459.090 3229.760 ;
        RECT 13.870 466.380 14.190 466.440 ;
        RECT 23.990 466.380 24.310 466.440 ;
        RECT 13.870 466.240 24.310 466.380 ;
        RECT 13.870 466.180 14.190 466.240 ;
        RECT 23.990 466.180 24.310 466.240 ;
      LAYER via ;
        RECT 24.020 3229.700 24.280 3229.960 ;
        RECT 2458.800 3229.700 2459.060 3229.960 ;
        RECT 13.900 466.180 14.160 466.440 ;
        RECT 24.020 466.180 24.280 466.440 ;
      LAYER met2 ;
        RECT 24.020 3229.670 24.280 3229.990 ;
        RECT 2458.800 3229.670 2459.060 3229.990 ;
        RECT 24.080 466.470 24.220 3229.670 ;
        RECT 2458.860 3220.000 2459.000 3229.670 ;
        RECT 2458.840 3216.000 2459.120 3220.000 ;
        RECT 13.900 466.325 14.160 466.470 ;
        RECT 13.890 465.955 14.170 466.325 ;
        RECT 24.020 466.150 24.280 466.470 ;
      LAYER via2 ;
        RECT 13.890 466.000 14.170 466.280 ;
      LAYER met3 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 13.865 466.290 14.195 466.305 ;
        RECT -4.800 465.990 14.195 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 13.865 465.975 14.195 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.110 3230.155 17.390 3230.525 ;
        RECT 2522.270 3230.155 2522.550 3230.525 ;
        RECT 17.180 250.765 17.320 3230.155 ;
        RECT 2522.340 3220.000 2522.480 3230.155 ;
        RECT 2522.320 3216.000 2522.600 3220.000 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 17.110 3230.200 17.390 3230.480 ;
        RECT 2522.270 3230.200 2522.550 3230.480 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT 17.085 3230.490 17.415 3230.505 ;
        RECT 2522.245 3230.490 2522.575 3230.505 ;
        RECT 17.085 3230.190 2522.575 3230.490 ;
        RECT 17.085 3230.175 17.415 3230.190 ;
        RECT 2522.245 3230.175 2522.575 3230.190 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.450 3216.810 2583.730 3216.925 ;
        RECT 2585.340 3216.810 2585.620 3220.000 ;
        RECT 2583.450 3216.670 2585.620 3216.810 ;
        RECT 2583.450 3216.555 2583.730 3216.670 ;
        RECT 2585.340 3216.000 2585.620 3216.670 ;
        RECT 17.110 40.955 17.390 41.325 ;
        RECT 17.180 35.885 17.320 40.955 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 2583.450 3216.600 2583.730 3216.880 ;
        RECT 17.110 41.000 17.390 41.280 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 2581.790 3216.890 2582.170 3216.900 ;
        RECT 2583.425 3216.890 2583.755 3216.905 ;
        RECT 2581.790 3216.590 2583.755 3216.890 ;
        RECT 2581.790 3216.580 2582.170 3216.590 ;
        RECT 2583.425 3216.575 2583.755 3216.590 ;
        RECT 17.085 41.290 17.415 41.305 ;
        RECT 2581.790 41.290 2582.170 41.300 ;
        RECT 17.085 40.990 2582.170 41.290 ;
        RECT 17.085 40.975 17.415 40.990 ;
        RECT 2581.790 40.980 2582.170 40.990 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
      LAYER via3 ;
        RECT 2581.820 3216.580 2582.140 3216.900 ;
        RECT 2581.820 40.980 2582.140 41.300 ;
      LAYER met4 ;
        RECT 2581.815 3216.575 2582.145 3216.905 ;
        RECT 2581.830 41.305 2582.130 3216.575 ;
        RECT 2581.815 40.975 2582.145 41.305 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 439.370 3216.980 439.690 3217.040 ;
        RECT 2618.850 3216.980 2619.170 3217.040 ;
        RECT 439.370 3216.840 2619.170 3216.980 ;
        RECT 439.370 3216.780 439.690 3216.840 ;
        RECT 2618.850 3216.780 2619.170 3216.840 ;
        RECT 2618.850 910.760 2619.170 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 2618.850 910.620 2901.150 910.760 ;
        RECT 2618.850 910.560 2619.170 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 439.400 3216.780 439.660 3217.040 ;
        RECT 2618.880 3216.780 2619.140 3217.040 ;
        RECT 2618.880 910.560 2619.140 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 438.060 3216.810 438.340 3220.000 ;
        RECT 439.400 3216.810 439.660 3217.070 ;
        RECT 438.060 3216.750 439.660 3216.810 ;
        RECT 2618.880 3216.750 2619.140 3217.070 ;
        RECT 438.060 3216.670 439.600 3216.750 ;
        RECT 438.060 3216.000 438.340 3216.670 ;
        RECT 2618.940 910.850 2619.080 3216.750 ;
        RECT 2618.880 910.530 2619.140 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2625.750 1145.360 2626.070 1145.420 ;
        RECT 2900.830 1145.360 2901.150 1145.420 ;
        RECT 2625.750 1145.220 2901.150 1145.360 ;
        RECT 2625.750 1145.160 2626.070 1145.220 ;
        RECT 2900.830 1145.160 2901.150 1145.220 ;
      LAYER via ;
        RECT 2625.780 1145.160 2626.040 1145.420 ;
        RECT 2900.860 1145.160 2901.120 1145.420 ;
      LAYER met2 ;
        RECT 501.080 3216.810 501.360 3220.000 ;
        RECT 502.410 3216.810 502.690 3216.925 ;
        RECT 501.080 3216.670 502.690 3216.810 ;
        RECT 501.080 3216.000 501.360 3216.670 ;
        RECT 502.410 3216.555 502.690 3216.670 ;
        RECT 2625.770 3213.835 2626.050 3214.205 ;
        RECT 2625.840 1145.450 2625.980 3213.835 ;
        RECT 2625.780 1145.130 2626.040 1145.450 ;
        RECT 2900.860 1145.130 2901.120 1145.450 ;
        RECT 2900.920 1144.285 2901.060 1145.130 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
      LAYER via2 ;
        RECT 502.410 3216.600 502.690 3216.880 ;
        RECT 2625.770 3213.880 2626.050 3214.160 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
      LAYER met3 ;
        RECT 502.385 3216.900 502.715 3216.905 ;
        RECT 502.385 3216.890 502.970 3216.900 ;
        RECT 502.385 3216.590 503.170 3216.890 ;
        RECT 502.385 3216.580 502.970 3216.590 ;
        RECT 502.385 3216.575 502.715 3216.580 ;
        RECT 502.590 3214.170 502.970 3214.180 ;
        RECT 2625.745 3214.170 2626.075 3214.185 ;
        RECT 502.590 3213.870 2626.075 3214.170 ;
        RECT 502.590 3213.860 502.970 3213.870 ;
        RECT 2625.745 3213.855 2626.075 3213.870 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
      LAYER via3 ;
        RECT 502.620 3216.580 502.940 3216.900 ;
        RECT 502.620 3213.860 502.940 3214.180 ;
      LAYER met4 ;
        RECT 502.615 3216.575 502.945 3216.905 ;
        RECT 502.630 3214.185 502.930 3216.575 ;
        RECT 502.615 3213.855 502.945 3214.185 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2766.510 1374.180 2766.830 1374.240 ;
        RECT 2801.010 1374.180 2801.330 1374.240 ;
        RECT 2766.510 1374.040 2801.330 1374.180 ;
        RECT 2766.510 1373.980 2766.830 1374.040 ;
        RECT 2801.010 1373.980 2801.330 1374.040 ;
      LAYER via ;
        RECT 2766.540 1373.980 2766.800 1374.240 ;
        RECT 2801.040 1373.980 2801.300 1374.240 ;
      LAYER met2 ;
        RECT 564.510 3231.515 564.790 3231.885 ;
        RECT 564.580 3220.000 564.720 3231.515 ;
        RECT 564.560 3216.000 564.840 3220.000 ;
        RECT 2745.830 1375.115 2746.110 1375.485 ;
        RECT 2632.210 1374.435 2632.490 1374.805 ;
        RECT 2669.930 1374.435 2670.210 1374.805 ;
        RECT 2632.280 1372.085 2632.420 1374.435 ;
        RECT 2670.000 1374.010 2670.140 1374.435 ;
        RECT 2670.850 1374.010 2671.130 1374.125 ;
        RECT 2670.000 1373.870 2671.130 1374.010 ;
        RECT 2670.850 1373.755 2671.130 1373.870 ;
        RECT 2745.900 1373.445 2746.040 1375.115 ;
        RECT 2801.030 1374.435 2801.310 1374.805 ;
        RECT 2801.100 1374.270 2801.240 1374.435 ;
        RECT 2766.540 1374.125 2766.800 1374.270 ;
        RECT 2766.530 1373.755 2766.810 1374.125 ;
        RECT 2801.040 1373.950 2801.300 1374.270 ;
        RECT 2745.830 1373.075 2746.110 1373.445 ;
        RECT 2632.210 1371.715 2632.490 1372.085 ;
      LAYER via2 ;
        RECT 564.510 3231.560 564.790 3231.840 ;
        RECT 2745.830 1375.160 2746.110 1375.440 ;
        RECT 2632.210 1374.480 2632.490 1374.760 ;
        RECT 2669.930 1374.480 2670.210 1374.760 ;
        RECT 2670.850 1373.800 2671.130 1374.080 ;
        RECT 2801.030 1374.480 2801.310 1374.760 ;
        RECT 2766.530 1373.800 2766.810 1374.080 ;
        RECT 2745.830 1373.120 2746.110 1373.400 ;
        RECT 2632.210 1371.760 2632.490 1372.040 ;
      LAYER met3 ;
        RECT 564.485 3231.850 564.815 3231.865 ;
        RECT 2604.790 3231.850 2605.170 3231.860 ;
        RECT 564.485 3231.550 2605.170 3231.850 ;
        RECT 564.485 3231.535 564.815 3231.550 ;
        RECT 2604.790 3231.540 2605.170 3231.550 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2916.710 1378.550 2924.800 1378.850 ;
        RECT 2697.710 1375.450 2698.090 1375.460 ;
        RECT 2745.805 1375.450 2746.135 1375.465 ;
        RECT 2697.710 1375.150 2746.135 1375.450 ;
        RECT 2697.710 1375.140 2698.090 1375.150 ;
        RECT 2745.805 1375.135 2746.135 1375.150 ;
        RECT 2632.185 1374.770 2632.515 1374.785 ;
        RECT 2669.905 1374.770 2670.235 1374.785 ;
        RECT 2632.185 1374.470 2670.235 1374.770 ;
        RECT 2632.185 1374.455 2632.515 1374.470 ;
        RECT 2669.905 1374.455 2670.235 1374.470 ;
        RECT 2801.005 1374.770 2801.335 1374.785 ;
        RECT 2801.005 1374.470 2836.050 1374.770 ;
        RECT 2801.005 1374.455 2801.335 1374.470 ;
        RECT 2670.825 1374.090 2671.155 1374.105 ;
        RECT 2697.710 1374.090 2698.090 1374.100 ;
        RECT 2766.505 1374.090 2766.835 1374.105 ;
        RECT 2670.825 1373.790 2698.090 1374.090 ;
        RECT 2670.825 1373.775 2671.155 1373.790 ;
        RECT 2697.710 1373.780 2698.090 1373.790 ;
        RECT 2752.950 1373.790 2766.835 1374.090 ;
        RECT 2835.750 1374.090 2836.050 1374.470 ;
        RECT 2916.710 1374.090 2917.010 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
        RECT 2835.750 1373.790 2883.890 1374.090 ;
        RECT 2607.550 1373.410 2607.930 1373.420 ;
        RECT 2745.805 1373.410 2746.135 1373.425 ;
        RECT 2752.950 1373.410 2753.250 1373.790 ;
        RECT 2766.505 1373.775 2766.835 1373.790 ;
        RECT 2607.550 1373.110 2608.810 1373.410 ;
        RECT 2607.550 1373.100 2607.930 1373.110 ;
        RECT 2608.510 1372.050 2608.810 1373.110 ;
        RECT 2745.805 1373.110 2753.250 1373.410 ;
        RECT 2883.590 1373.410 2883.890 1373.790 ;
        RECT 2884.510 1373.790 2917.010 1374.090 ;
        RECT 2884.510 1373.410 2884.810 1373.790 ;
        RECT 2883.590 1373.110 2884.810 1373.410 ;
        RECT 2745.805 1373.095 2746.135 1373.110 ;
        RECT 2632.185 1372.050 2632.515 1372.065 ;
        RECT 2608.510 1371.750 2632.515 1372.050 ;
        RECT 2632.185 1371.735 2632.515 1371.750 ;
      LAYER via3 ;
        RECT 2604.820 3231.540 2605.140 3231.860 ;
        RECT 2697.740 1375.140 2698.060 1375.460 ;
        RECT 2697.740 1373.780 2698.060 1374.100 ;
        RECT 2607.580 1373.100 2607.900 1373.420 ;
      LAYER met4 ;
        RECT 2604.815 3231.535 2605.145 3231.865 ;
        RECT 2604.830 1395.850 2605.130 3231.535 ;
        RECT 2604.830 1395.550 2606.970 1395.850 ;
        RECT 2606.670 1372.050 2606.970 1395.550 ;
        RECT 2697.735 1375.135 2698.065 1375.465 ;
        RECT 2697.750 1374.105 2698.050 1375.135 ;
        RECT 2697.735 1373.775 2698.065 1374.105 ;
        RECT 2607.575 1373.095 2607.905 1373.425 ;
        RECT 2607.590 1372.050 2607.890 1373.095 ;
        RECT 2606.670 1371.750 2607.890 1372.050 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.510 3235.680 627.830 3235.740 ;
        RECT 840.950 3235.680 841.270 3235.740 ;
        RECT 627.510 3235.540 841.270 3235.680 ;
        RECT 627.510 3235.480 627.830 3235.540 ;
        RECT 840.950 3235.480 841.270 3235.540 ;
        RECT 840.950 3226.160 841.270 3226.220 ;
        RECT 2903.590 3226.160 2903.910 3226.220 ;
        RECT 840.950 3226.020 2903.910 3226.160 ;
        RECT 840.950 3225.960 841.270 3226.020 ;
        RECT 2903.590 3225.960 2903.910 3226.020 ;
      LAYER via ;
        RECT 627.540 3235.480 627.800 3235.740 ;
        RECT 840.980 3235.480 841.240 3235.740 ;
        RECT 840.980 3225.960 841.240 3226.220 ;
        RECT 2903.620 3225.960 2903.880 3226.220 ;
      LAYER met2 ;
        RECT 627.540 3235.450 627.800 3235.770 ;
        RECT 840.980 3235.450 841.240 3235.770 ;
        RECT 627.600 3220.000 627.740 3235.450 ;
        RECT 841.040 3226.250 841.180 3235.450 ;
        RECT 840.980 3225.930 841.240 3226.250 ;
        RECT 2903.620 3225.930 2903.880 3226.250 ;
        RECT 627.580 3216.000 627.860 3220.000 ;
        RECT 2903.680 1613.485 2903.820 3225.930 ;
        RECT 2903.610 1613.115 2903.890 1613.485 ;
      LAYER via2 ;
        RECT 2903.610 1613.160 2903.890 1613.440 ;
      LAYER met3 ;
        RECT 2903.585 1613.450 2903.915 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2903.585 1613.150 2924.800 1613.450 ;
        RECT 2903.585 1613.135 2903.915 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 690.530 3233.300 690.850 3233.360 ;
        RECT 2627.130 3233.300 2627.450 3233.360 ;
        RECT 690.530 3233.160 2627.450 3233.300 ;
        RECT 690.530 3233.100 690.850 3233.160 ;
        RECT 2627.130 3233.100 2627.450 3233.160 ;
        RECT 2627.130 1849.160 2627.450 1849.220 ;
        RECT 2900.830 1849.160 2901.150 1849.220 ;
        RECT 2627.130 1849.020 2901.150 1849.160 ;
        RECT 2627.130 1848.960 2627.450 1849.020 ;
        RECT 2900.830 1848.960 2901.150 1849.020 ;
      LAYER via ;
        RECT 690.560 3233.100 690.820 3233.360 ;
        RECT 2627.160 3233.100 2627.420 3233.360 ;
        RECT 2627.160 1848.960 2627.420 1849.220 ;
        RECT 2900.860 1848.960 2901.120 1849.220 ;
      LAYER met2 ;
        RECT 690.560 3233.070 690.820 3233.390 ;
        RECT 2627.160 3233.070 2627.420 3233.390 ;
        RECT 690.620 3220.000 690.760 3233.070 ;
        RECT 690.600 3216.000 690.880 3220.000 ;
        RECT 2627.220 1849.250 2627.360 3233.070 ;
        RECT 2627.160 1848.930 2627.420 1849.250 ;
        RECT 2900.860 1848.930 2901.120 1849.250 ;
        RECT 2900.920 1848.085 2901.060 1848.930 ;
        RECT 2900.850 1847.715 2901.130 1848.085 ;
      LAYER via2 ;
        RECT 2900.850 1847.760 2901.130 1848.040 ;
      LAYER met3 ;
        RECT 2900.825 1848.050 2901.155 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2900.825 1847.750 2924.800 1848.050 ;
        RECT 2900.825 1847.735 2901.155 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 754.010 3234.660 754.330 3234.720 ;
        RECT 2627.590 3234.660 2627.910 3234.720 ;
        RECT 754.010 3234.520 2627.910 3234.660 ;
        RECT 754.010 3234.460 754.330 3234.520 ;
        RECT 2627.590 3234.460 2627.910 3234.520 ;
        RECT 2627.590 2083.760 2627.910 2083.820 ;
        RECT 2900.830 2083.760 2901.150 2083.820 ;
        RECT 2627.590 2083.620 2901.150 2083.760 ;
        RECT 2627.590 2083.560 2627.910 2083.620 ;
        RECT 2900.830 2083.560 2901.150 2083.620 ;
      LAYER via ;
        RECT 754.040 3234.460 754.300 3234.720 ;
        RECT 2627.620 3234.460 2627.880 3234.720 ;
        RECT 2627.620 2083.560 2627.880 2083.820 ;
        RECT 2900.860 2083.560 2901.120 2083.820 ;
      LAYER met2 ;
        RECT 754.040 3234.430 754.300 3234.750 ;
        RECT 2627.620 3234.430 2627.880 3234.750 ;
        RECT 754.100 3220.000 754.240 3234.430 ;
        RECT 754.080 3216.000 754.360 3220.000 ;
        RECT 2627.680 2083.850 2627.820 3234.430 ;
        RECT 2627.620 2083.530 2627.880 2083.850 ;
        RECT 2900.860 2083.530 2901.120 2083.850 ;
        RECT 2900.920 2082.685 2901.060 2083.530 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
      LAYER met3 ;
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2766.510 2312.580 2766.830 2312.640 ;
        RECT 2801.010 2312.580 2801.330 2312.640 ;
        RECT 2766.510 2312.440 2801.330 2312.580 ;
        RECT 2766.510 2312.380 2766.830 2312.440 ;
        RECT 2801.010 2312.380 2801.330 2312.440 ;
      LAYER via ;
        RECT 2766.540 2312.380 2766.800 2312.640 ;
        RECT 2801.040 2312.380 2801.300 2312.640 ;
      LAYER met2 ;
        RECT 817.050 3232.195 817.330 3232.565 ;
        RECT 817.120 3220.000 817.260 3232.195 ;
        RECT 817.100 3216.000 817.380 3220.000 ;
        RECT 2745.830 2313.515 2746.110 2313.885 ;
        RECT 2632.210 2312.835 2632.490 2313.205 ;
        RECT 2669.930 2312.835 2670.210 2313.205 ;
        RECT 2632.280 2310.485 2632.420 2312.835 ;
        RECT 2670.000 2312.410 2670.140 2312.835 ;
        RECT 2670.850 2312.410 2671.130 2312.525 ;
        RECT 2670.000 2312.270 2671.130 2312.410 ;
        RECT 2670.850 2312.155 2671.130 2312.270 ;
        RECT 2745.900 2311.845 2746.040 2313.515 ;
        RECT 2801.030 2312.835 2801.310 2313.205 ;
        RECT 2801.100 2312.670 2801.240 2312.835 ;
        RECT 2766.540 2312.525 2766.800 2312.670 ;
        RECT 2766.530 2312.155 2766.810 2312.525 ;
        RECT 2801.040 2312.350 2801.300 2312.670 ;
        RECT 2745.830 2311.475 2746.110 2311.845 ;
        RECT 2632.210 2310.115 2632.490 2310.485 ;
      LAYER via2 ;
        RECT 817.050 3232.240 817.330 3232.520 ;
        RECT 2745.830 2313.560 2746.110 2313.840 ;
        RECT 2632.210 2312.880 2632.490 2313.160 ;
        RECT 2669.930 2312.880 2670.210 2313.160 ;
        RECT 2670.850 2312.200 2671.130 2312.480 ;
        RECT 2801.030 2312.880 2801.310 2313.160 ;
        RECT 2766.530 2312.200 2766.810 2312.480 ;
        RECT 2745.830 2311.520 2746.110 2311.800 ;
        RECT 2632.210 2310.160 2632.490 2310.440 ;
      LAYER met3 ;
        RECT 817.025 3232.530 817.355 3232.545 ;
        RECT 2605.710 3232.530 2606.090 3232.540 ;
        RECT 817.025 3232.230 2606.090 3232.530 ;
        RECT 817.025 3232.215 817.355 3232.230 ;
        RECT 2605.710 3232.220 2606.090 3232.230 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2916.710 2316.950 2924.800 2317.250 ;
        RECT 2697.710 2313.850 2698.090 2313.860 ;
        RECT 2745.805 2313.850 2746.135 2313.865 ;
        RECT 2697.710 2313.550 2746.135 2313.850 ;
        RECT 2697.710 2313.540 2698.090 2313.550 ;
        RECT 2745.805 2313.535 2746.135 2313.550 ;
        RECT 2632.185 2313.170 2632.515 2313.185 ;
        RECT 2669.905 2313.170 2670.235 2313.185 ;
        RECT 2632.185 2312.870 2670.235 2313.170 ;
        RECT 2632.185 2312.855 2632.515 2312.870 ;
        RECT 2669.905 2312.855 2670.235 2312.870 ;
        RECT 2801.005 2313.170 2801.335 2313.185 ;
        RECT 2801.005 2312.870 2836.050 2313.170 ;
        RECT 2801.005 2312.855 2801.335 2312.870 ;
        RECT 2670.825 2312.490 2671.155 2312.505 ;
        RECT 2697.710 2312.490 2698.090 2312.500 ;
        RECT 2766.505 2312.490 2766.835 2312.505 ;
        RECT 2670.825 2312.190 2698.090 2312.490 ;
        RECT 2670.825 2312.175 2671.155 2312.190 ;
        RECT 2697.710 2312.180 2698.090 2312.190 ;
        RECT 2752.950 2312.190 2766.835 2312.490 ;
        RECT 2835.750 2312.490 2836.050 2312.870 ;
        RECT 2916.710 2312.490 2917.010 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 2835.750 2312.190 2883.890 2312.490 ;
        RECT 2607.550 2311.810 2607.930 2311.820 ;
        RECT 2745.805 2311.810 2746.135 2311.825 ;
        RECT 2752.950 2311.810 2753.250 2312.190 ;
        RECT 2766.505 2312.175 2766.835 2312.190 ;
        RECT 2607.550 2311.510 2608.810 2311.810 ;
        RECT 2607.550 2311.500 2607.930 2311.510 ;
        RECT 2608.510 2310.450 2608.810 2311.510 ;
        RECT 2745.805 2311.510 2753.250 2311.810 ;
        RECT 2883.590 2311.810 2883.890 2312.190 ;
        RECT 2884.510 2312.190 2917.010 2312.490 ;
        RECT 2884.510 2311.810 2884.810 2312.190 ;
        RECT 2883.590 2311.510 2884.810 2311.810 ;
        RECT 2745.805 2311.495 2746.135 2311.510 ;
        RECT 2632.185 2310.450 2632.515 2310.465 ;
        RECT 2608.510 2310.150 2632.515 2310.450 ;
        RECT 2632.185 2310.135 2632.515 2310.150 ;
      LAYER via3 ;
        RECT 2605.740 3232.220 2606.060 3232.540 ;
        RECT 2697.740 2313.540 2698.060 2313.860 ;
        RECT 2697.740 2312.180 2698.060 2312.500 ;
        RECT 2607.580 2311.500 2607.900 2311.820 ;
      LAYER met4 ;
        RECT 2605.735 3232.215 2606.065 3232.545 ;
        RECT 2605.750 2324.050 2606.050 3232.215 ;
        RECT 2605.750 2323.750 2606.970 2324.050 ;
        RECT 2606.670 2310.450 2606.970 2323.750 ;
        RECT 2697.735 2313.535 2698.065 2313.865 ;
        RECT 2697.750 2312.505 2698.050 2313.535 ;
        RECT 2697.735 2312.175 2698.065 2312.505 ;
        RECT 2607.575 2311.495 2607.905 2311.825 ;
        RECT 2607.590 2310.450 2607.890 2311.495 ;
        RECT 2606.670 2310.150 2607.890 2310.450 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.650 3234.235 269.930 3234.605 ;
        RECT 2901.310 3234.235 2901.590 3234.605 ;
        RECT 269.720 3220.000 269.860 3234.235 ;
        RECT 269.700 3216.000 269.980 3220.000 ;
        RECT 2901.380 146.725 2901.520 3234.235 ;
        RECT 2901.310 146.355 2901.590 146.725 ;
      LAYER via2 ;
        RECT 269.650 3234.280 269.930 3234.560 ;
        RECT 2901.310 3234.280 2901.590 3234.560 ;
        RECT 2901.310 146.400 2901.590 146.680 ;
      LAYER met3 ;
        RECT 269.625 3234.570 269.955 3234.585 ;
        RECT 2901.285 3234.570 2901.615 3234.585 ;
        RECT 269.625 3234.270 2901.615 3234.570 ;
        RECT 269.625 3234.255 269.955 3234.270 ;
        RECT 2901.285 3234.255 2901.615 3234.270 ;
        RECT 2901.285 146.690 2901.615 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2901.285 146.390 2924.800 146.690 ;
        RECT 2901.285 146.375 2901.615 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 901.210 3236.020 901.530 3236.080 ;
        RECT 1932.990 3236.020 1933.310 3236.080 ;
        RECT 901.210 3235.880 1933.310 3236.020 ;
        RECT 901.210 3235.820 901.530 3235.880 ;
        RECT 1932.990 3235.820 1933.310 3235.880 ;
        RECT 1932.990 3227.520 1933.310 3227.580 ;
        RECT 2904.050 3227.520 2904.370 3227.580 ;
        RECT 1932.990 3227.380 2904.370 3227.520 ;
        RECT 1932.990 3227.320 1933.310 3227.380 ;
        RECT 2904.050 3227.320 2904.370 3227.380 ;
      LAYER via ;
        RECT 901.240 3235.820 901.500 3236.080 ;
        RECT 1933.020 3235.820 1933.280 3236.080 ;
        RECT 1933.020 3227.320 1933.280 3227.580 ;
        RECT 2904.080 3227.320 2904.340 3227.580 ;
      LAYER met2 ;
        RECT 901.240 3235.790 901.500 3236.110 ;
        RECT 1933.020 3235.790 1933.280 3236.110 ;
        RECT 901.300 3220.000 901.440 3235.790 ;
        RECT 1933.080 3227.610 1933.220 3235.790 ;
        RECT 1933.020 3227.290 1933.280 3227.610 ;
        RECT 2904.080 3227.290 2904.340 3227.610 ;
        RECT 901.280 3216.000 901.560 3220.000 ;
        RECT 2904.140 2493.405 2904.280 3227.290 ;
        RECT 2904.070 2493.035 2904.350 2493.405 ;
      LAYER via2 ;
        RECT 2904.070 2493.080 2904.350 2493.360 ;
      LAYER met3 ;
        RECT 2904.045 2493.370 2904.375 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2904.045 2493.070 2924.800 2493.370 ;
        RECT 2904.045 2493.055 2904.375 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 964.230 3221.060 964.550 3221.120 ;
        RECT 2659.790 3221.060 2660.110 3221.120 ;
        RECT 964.230 3220.920 2660.110 3221.060 ;
        RECT 964.230 3220.860 964.550 3220.920 ;
        RECT 2659.790 3220.860 2660.110 3220.920 ;
        RECT 2659.790 2732.140 2660.110 2732.200 ;
        RECT 2899.910 2732.140 2900.230 2732.200 ;
        RECT 2659.790 2732.000 2900.230 2732.140 ;
        RECT 2659.790 2731.940 2660.110 2732.000 ;
        RECT 2899.910 2731.940 2900.230 2732.000 ;
      LAYER via ;
        RECT 964.260 3220.860 964.520 3221.120 ;
        RECT 2659.820 3220.860 2660.080 3221.120 ;
        RECT 2659.820 2731.940 2660.080 2732.200 ;
        RECT 2899.940 2731.940 2900.200 2732.200 ;
      LAYER met2 ;
        RECT 964.260 3220.830 964.520 3221.150 ;
        RECT 2659.820 3220.830 2660.080 3221.150 ;
        RECT 964.320 3220.000 964.460 3220.830 ;
        RECT 964.300 3216.000 964.580 3220.000 ;
        RECT 2659.880 2732.230 2660.020 3220.830 ;
        RECT 2659.820 2731.910 2660.080 2732.230 ;
        RECT 2899.940 2731.910 2900.200 2732.230 ;
        RECT 2900.000 2728.005 2900.140 2731.910 ;
        RECT 2899.930 2727.635 2900.210 2728.005 ;
      LAYER via2 ;
        RECT 2899.930 2727.680 2900.210 2727.960 ;
      LAYER met3 ;
        RECT 2899.905 2727.970 2900.235 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2899.905 2727.670 2924.800 2727.970 ;
        RECT 2899.905 2727.655 2900.235 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2721.890 2966.740 2722.210 2966.800 ;
        RECT 2899.910 2966.740 2900.230 2966.800 ;
        RECT 2721.890 2966.600 2900.230 2966.740 ;
        RECT 2721.890 2966.540 2722.210 2966.600 ;
        RECT 2899.910 2966.540 2900.230 2966.600 ;
      LAYER via ;
        RECT 2721.920 2966.540 2722.180 2966.800 ;
        RECT 2899.940 2966.540 2900.200 2966.800 ;
      LAYER met2 ;
        RECT 1027.270 3216.810 1027.550 3216.925 ;
        RECT 1027.780 3216.810 1028.060 3220.000 ;
        RECT 1027.270 3216.670 1028.060 3216.810 ;
        RECT 1027.270 3216.555 1027.550 3216.670 ;
        RECT 1027.780 3216.000 1028.060 3216.670 ;
        RECT 2721.910 3209.075 2722.190 3209.445 ;
        RECT 2721.980 2966.830 2722.120 3209.075 ;
        RECT 2721.920 2966.510 2722.180 2966.830 ;
        RECT 2899.940 2966.510 2900.200 2966.830 ;
        RECT 2900.000 2962.605 2900.140 2966.510 ;
        RECT 2899.930 2962.235 2900.210 2962.605 ;
      LAYER via2 ;
        RECT 1027.270 3216.600 1027.550 3216.880 ;
        RECT 2721.910 3209.120 2722.190 3209.400 ;
        RECT 2899.930 2962.280 2900.210 2962.560 ;
      LAYER met3 ;
        RECT 1027.245 3216.900 1027.575 3216.905 ;
        RECT 1026.990 3216.890 1027.575 3216.900 ;
        RECT 1026.790 3216.590 1027.575 3216.890 ;
        RECT 1026.990 3216.580 1027.575 3216.590 ;
        RECT 1027.245 3216.575 1027.575 3216.580 ;
        RECT 1026.990 3209.410 1027.370 3209.420 ;
        RECT 2721.885 3209.410 2722.215 3209.425 ;
        RECT 1026.990 3209.110 2722.215 3209.410 ;
        RECT 1026.990 3209.100 1027.370 3209.110 ;
        RECT 2721.885 3209.095 2722.215 3209.110 ;
        RECT 2899.905 2962.570 2900.235 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2899.905 2962.270 2924.800 2962.570 ;
        RECT 2899.905 2962.255 2900.235 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
      LAYER via3 ;
        RECT 1027.020 3216.580 1027.340 3216.900 ;
        RECT 1027.020 3209.100 1027.340 3209.420 ;
      LAYER met4 ;
        RECT 1027.015 3216.575 1027.345 3216.905 ;
        RECT 1027.030 3209.425 1027.330 3216.575 ;
        RECT 1027.015 3209.095 1027.345 3209.425 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2859.890 3201.340 2860.210 3201.400 ;
        RECT 2900.830 3201.340 2901.150 3201.400 ;
        RECT 2859.890 3201.200 2901.150 3201.340 ;
        RECT 2859.890 3201.140 2860.210 3201.200 ;
        RECT 2900.830 3201.140 2901.150 3201.200 ;
      LAYER via ;
        RECT 2859.920 3201.140 2860.180 3201.400 ;
        RECT 2900.860 3201.140 2901.120 3201.400 ;
      LAYER met2 ;
        RECT 1090.800 3216.810 1091.080 3220.000 ;
        RECT 1092.130 3216.810 1092.410 3216.925 ;
        RECT 1090.800 3216.670 1092.410 3216.810 ;
        RECT 1090.800 3216.000 1091.080 3216.670 ;
        RECT 1092.130 3216.555 1092.410 3216.670 ;
        RECT 2859.910 3209.755 2860.190 3210.125 ;
        RECT 2859.980 3201.430 2860.120 3209.755 ;
        RECT 2859.920 3201.110 2860.180 3201.430 ;
        RECT 2900.860 3201.110 2901.120 3201.430 ;
        RECT 2900.920 3197.205 2901.060 3201.110 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
      LAYER via2 ;
        RECT 1092.130 3216.600 1092.410 3216.880 ;
        RECT 2859.910 3209.800 2860.190 3210.080 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
      LAYER met3 ;
        RECT 1092.105 3216.900 1092.435 3216.905 ;
        RECT 1092.105 3216.890 1092.690 3216.900 ;
        RECT 1092.105 3216.590 1092.890 3216.890 ;
        RECT 1092.105 3216.580 1092.690 3216.590 ;
        RECT 1092.105 3216.575 1092.435 3216.580 ;
        RECT 1092.310 3210.090 1092.690 3210.100 ;
        RECT 2859.885 3210.090 2860.215 3210.105 ;
        RECT 1092.310 3209.790 2860.215 3210.090 ;
        RECT 1092.310 3209.780 1092.690 3209.790 ;
        RECT 2859.885 3209.775 2860.215 3209.790 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
      LAYER via3 ;
        RECT 1092.340 3216.580 1092.660 3216.900 ;
        RECT 1092.340 3209.780 1092.660 3210.100 ;
      LAYER met4 ;
        RECT 1092.335 3216.575 1092.665 3216.905 ;
        RECT 1092.350 3210.105 1092.650 3216.575 ;
        RECT 1092.335 3209.775 1092.665 3210.105 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1497.460 3429.680 1506.340 3429.820 ;
        RECT 1158.810 3429.480 1159.130 3429.540 ;
        RECT 1497.460 3429.480 1497.600 3429.680 ;
        RECT 1158.810 3429.340 1497.600 3429.480 ;
        RECT 1506.200 3429.480 1506.340 3429.680 ;
        RECT 2146.060 3429.680 2149.880 3429.820 ;
        RECT 2146.060 3429.480 2146.200 3429.680 ;
        RECT 1506.200 3429.340 2146.200 3429.480 ;
        RECT 2149.740 3429.480 2149.880 3429.680 ;
        RECT 2762.920 3429.680 2798.940 3429.820 ;
        RECT 2762.920 3429.480 2763.060 3429.680 ;
        RECT 2149.740 3429.340 2763.060 3429.480 ;
        RECT 2798.800 3429.480 2798.940 3429.680 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2798.800 3429.340 2901.150 3429.480 ;
        RECT 1158.810 3429.280 1159.130 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 1158.840 3429.280 1159.100 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 1158.840 3429.250 1159.100 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 1153.820 3218.850 1154.100 3220.000 ;
        RECT 1158.900 3218.850 1159.040 3429.250 ;
        RECT 1153.820 3218.710 1159.040 3218.850 ;
        RECT 1153.820 3216.000 1154.100 3218.710 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1220.910 3501.900 1221.230 3501.960 ;
        RECT 2717.290 3501.900 2717.610 3501.960 ;
        RECT 1220.910 3501.760 2717.610 3501.900 ;
        RECT 1220.910 3501.700 1221.230 3501.760 ;
        RECT 2717.290 3501.700 2717.610 3501.760 ;
      LAYER via ;
        RECT 1220.940 3501.700 1221.200 3501.960 ;
        RECT 2717.320 3501.700 2717.580 3501.960 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.990 2717.520 3517.600 ;
        RECT 1220.940 3501.670 1221.200 3501.990 ;
        RECT 2717.320 3501.670 2717.580 3501.990 ;
        RECT 1216.840 3218.850 1217.120 3220.000 ;
        RECT 1221.000 3218.850 1221.140 3501.670 ;
        RECT 1216.840 3218.710 1221.140 3218.850 ;
        RECT 1216.840 3216.000 1217.120 3218.710 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.010 3503.600 1283.330 3503.660 ;
        RECT 2392.530 3503.600 2392.850 3503.660 ;
        RECT 1283.010 3503.460 2392.850 3503.600 ;
        RECT 1283.010 3503.400 1283.330 3503.460 ;
        RECT 2392.530 3503.400 2392.850 3503.460 ;
      LAYER via ;
        RECT 1283.040 3503.400 1283.300 3503.660 ;
        RECT 2392.560 3503.400 2392.820 3503.660 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3503.690 2392.760 3517.600 ;
        RECT 1283.040 3503.370 1283.300 3503.690 ;
        RECT 2392.560 3503.370 2392.820 3503.690 ;
        RECT 1280.320 3218.850 1280.600 3220.000 ;
        RECT 1283.100 3218.850 1283.240 3503.370 ;
        RECT 1280.320 3218.710 1283.240 3218.850 ;
        RECT 1280.320 3216.000 1280.600 3218.710 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1345.110 3501.220 1345.430 3501.280 ;
        RECT 2068.230 3501.220 2068.550 3501.280 ;
        RECT 1345.110 3501.080 2068.550 3501.220 ;
        RECT 1345.110 3501.020 1345.430 3501.080 ;
        RECT 2068.230 3501.020 2068.550 3501.080 ;
      LAYER via ;
        RECT 1345.140 3501.020 1345.400 3501.280 ;
        RECT 2068.260 3501.020 2068.520 3501.280 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3501.310 2068.460 3517.600 ;
        RECT 1345.140 3500.990 1345.400 3501.310 ;
        RECT 2068.260 3500.990 2068.520 3501.310 ;
        RECT 1343.340 3219.530 1343.620 3220.000 ;
        RECT 1345.200 3219.530 1345.340 3500.990 ;
        RECT 1343.340 3219.390 1345.340 3219.530 ;
        RECT 1343.340 3216.000 1343.620 3219.390 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1407.210 3499.520 1407.530 3499.580 ;
        RECT 1743.930 3499.520 1744.250 3499.580 ;
        RECT 1407.210 3499.380 1744.250 3499.520 ;
        RECT 1407.210 3499.320 1407.530 3499.380 ;
        RECT 1743.930 3499.320 1744.250 3499.380 ;
      LAYER via ;
        RECT 1407.240 3499.320 1407.500 3499.580 ;
        RECT 1743.960 3499.320 1744.220 3499.580 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3499.610 1744.160 3517.600 ;
        RECT 1407.240 3499.290 1407.500 3499.610 ;
        RECT 1743.960 3499.290 1744.220 3499.610 ;
        RECT 1406.360 3219.530 1406.640 3220.000 ;
        RECT 1407.300 3219.530 1407.440 3499.290 ;
        RECT 1406.360 3219.390 1407.440 3219.530 ;
        RECT 1406.360 3216.000 1406.640 3219.390 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.170 3498.500 1419.490 3498.560 ;
        RECT 1469.770 3498.500 1470.090 3498.560 ;
        RECT 1419.170 3498.360 1470.090 3498.500 ;
        RECT 1419.170 3498.300 1419.490 3498.360 ;
        RECT 1469.770 3498.300 1470.090 3498.360 ;
      LAYER via ;
        RECT 1419.200 3498.300 1419.460 3498.560 ;
        RECT 1469.800 3498.300 1470.060 3498.560 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3498.590 1419.400 3517.600 ;
        RECT 1419.200 3498.270 1419.460 3498.590 ;
        RECT 1469.800 3498.270 1470.060 3498.590 ;
        RECT 1469.860 3220.000 1470.000 3498.270 ;
        RECT 1469.840 3216.000 1470.120 3220.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 628.965 3208.665 629.135 3218.695 ;
      LAYER mcon ;
        RECT 628.965 3218.525 629.135 3218.695 ;
      LAYER met1 ;
        RECT 628.890 3218.680 629.210 3218.740 ;
        RECT 628.695 3218.540 629.210 3218.680 ;
        RECT 628.890 3218.480 629.210 3218.540 ;
        RECT 628.905 3208.820 629.195 3208.865 ;
        RECT 2901.750 3208.820 2902.070 3208.880 ;
        RECT 628.905 3208.680 2902.070 3208.820 ;
        RECT 628.905 3208.635 629.195 3208.680 ;
        RECT 2901.750 3208.620 2902.070 3208.680 ;
      LAYER via ;
        RECT 628.920 3218.480 629.180 3218.740 ;
        RECT 2901.780 3208.620 2902.040 3208.880 ;
      LAYER met2 ;
        RECT 332.670 3232.195 332.950 3232.565 ;
        RECT 332.740 3220.000 332.880 3232.195 ;
        RECT 332.720 3216.000 333.000 3220.000 ;
        RECT 628.910 3218.595 629.190 3218.965 ;
        RECT 628.920 3218.450 629.180 3218.595 ;
        RECT 2901.780 3208.590 2902.040 3208.910 ;
        RECT 2901.840 381.325 2901.980 3208.590 ;
        RECT 2901.770 380.955 2902.050 381.325 ;
      LAYER via2 ;
        RECT 332.670 3232.240 332.950 3232.520 ;
        RECT 628.910 3218.640 629.190 3218.920 ;
        RECT 2901.770 381.000 2902.050 381.280 ;
      LAYER met3 ;
        RECT 332.645 3232.530 332.975 3232.545 ;
        RECT 628.630 3232.530 629.010 3232.540 ;
        RECT 332.645 3232.230 629.010 3232.530 ;
        RECT 332.645 3232.215 332.975 3232.230 ;
        RECT 628.630 3232.220 629.010 3232.230 ;
        RECT 628.885 3218.940 629.215 3218.945 ;
        RECT 628.630 3218.930 629.215 3218.940 ;
        RECT 628.430 3218.630 629.215 3218.930 ;
        RECT 628.630 3218.620 629.215 3218.630 ;
        RECT 628.885 3218.615 629.215 3218.620 ;
        RECT 2901.745 381.290 2902.075 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2901.745 380.990 2924.800 381.290 ;
        RECT 2901.745 380.975 2902.075 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
      LAYER via3 ;
        RECT 628.660 3232.220 628.980 3232.540 ;
        RECT 628.660 3218.620 628.980 3218.940 ;
      LAYER met4 ;
        RECT 628.655 3232.215 628.985 3232.545 ;
        RECT 628.670 3218.945 628.970 3232.215 ;
        RECT 628.655 3218.615 628.985 3218.945 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1094.870 3499.860 1095.190 3499.920 ;
        RECT 1531.870 3499.860 1532.190 3499.920 ;
        RECT 1094.870 3499.720 1532.190 3499.860 ;
        RECT 1094.870 3499.660 1095.190 3499.720 ;
        RECT 1531.870 3499.660 1532.190 3499.720 ;
      LAYER via ;
        RECT 1094.900 3499.660 1095.160 3499.920 ;
        RECT 1531.900 3499.660 1532.160 3499.920 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3499.950 1095.100 3517.600 ;
        RECT 1094.900 3499.630 1095.160 3499.950 ;
        RECT 1531.900 3499.630 1532.160 3499.950 ;
        RECT 1531.960 3219.530 1532.100 3499.630 ;
        RECT 1532.860 3219.530 1533.140 3220.000 ;
        RECT 1531.960 3219.390 1533.140 3219.530 ;
        RECT 1532.860 3216.000 1533.140 3219.390 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 770.570 3504.960 770.890 3505.020 ;
        RECT 1593.970 3504.960 1594.290 3505.020 ;
        RECT 770.570 3504.820 1594.290 3504.960 ;
        RECT 770.570 3504.760 770.890 3504.820 ;
        RECT 1593.970 3504.760 1594.290 3504.820 ;
      LAYER via ;
        RECT 770.600 3504.760 770.860 3505.020 ;
        RECT 1594.000 3504.760 1594.260 3505.020 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3505.050 770.800 3517.600 ;
        RECT 770.600 3504.730 770.860 3505.050 ;
        RECT 1594.000 3504.730 1594.260 3505.050 ;
        RECT 1594.060 3219.530 1594.200 3504.730 ;
        RECT 1595.880 3219.530 1596.160 3220.000 ;
        RECT 1594.060 3219.390 1596.160 3219.530 ;
        RECT 1595.880 3216.000 1596.160 3219.390 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3503.260 446.130 3503.320 ;
        RECT 1656.070 3503.260 1656.390 3503.320 ;
        RECT 445.810 3503.120 1656.390 3503.260 ;
        RECT 445.810 3503.060 446.130 3503.120 ;
        RECT 1656.070 3503.060 1656.390 3503.120 ;
      LAYER via ;
        RECT 445.840 3503.060 446.100 3503.320 ;
        RECT 1656.100 3503.060 1656.360 3503.320 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3503.350 446.040 3517.600 ;
        RECT 445.840 3503.030 446.100 3503.350 ;
        RECT 1656.100 3503.030 1656.360 3503.350 ;
        RECT 1656.160 3218.850 1656.300 3503.030 ;
        RECT 1658.900 3218.850 1659.180 3220.000 ;
        RECT 1656.160 3218.710 1659.180 3218.850 ;
        RECT 1658.900 3216.000 1659.180 3218.710 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3501.560 121.830 3501.620 ;
        RECT 1718.170 3501.560 1718.490 3501.620 ;
        RECT 121.510 3501.420 1718.490 3501.560 ;
        RECT 121.510 3501.360 121.830 3501.420 ;
        RECT 1718.170 3501.360 1718.490 3501.420 ;
      LAYER via ;
        RECT 121.540 3501.360 121.800 3501.620 ;
        RECT 1718.200 3501.360 1718.460 3501.620 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3501.650 121.740 3517.600 ;
        RECT 121.540 3501.330 121.800 3501.650 ;
        RECT 1718.200 3501.330 1718.460 3501.650 ;
        RECT 1718.260 3218.850 1718.400 3501.330 ;
        RECT 1722.380 3218.850 1722.660 3220.000 ;
        RECT 1718.260 3218.710 1722.660 3218.850 ;
        RECT 1722.380 3216.000 1722.660 3218.710 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 1780.270 3339.720 1780.590 3339.780 ;
        RECT 17.090 3339.580 1780.590 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 1780.270 3339.520 1780.590 3339.580 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 1780.300 3339.520 1780.560 3339.780 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 1780.300 3339.490 1780.560 3339.810 ;
        RECT 1780.360 3218.850 1780.500 3339.490 ;
        RECT 1785.400 3218.850 1785.680 3220.000 ;
        RECT 1780.360 3218.710 1785.680 3218.850 ;
        RECT 1785.400 3216.000 1785.680 3218.710 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 3056.500 16.950 3056.560 ;
        RECT 52.050 3056.500 52.370 3056.560 ;
        RECT 16.630 3056.360 52.370 3056.500 ;
        RECT 16.630 3056.300 16.950 3056.360 ;
        RECT 52.050 3056.300 52.370 3056.360 ;
      LAYER via ;
        RECT 16.660 3056.300 16.920 3056.560 ;
        RECT 52.080 3056.300 52.340 3056.560 ;
      LAYER met2 ;
        RECT 1846.990 3216.810 1847.270 3216.925 ;
        RECT 1848.420 3216.810 1848.700 3220.000 ;
        RECT 1846.990 3216.670 1848.700 3216.810 ;
        RECT 1846.990 3216.555 1847.270 3216.670 ;
        RECT 1848.420 3216.000 1848.700 3216.670 ;
        RECT 52.070 3210.435 52.350 3210.805 ;
        RECT 52.140 3056.590 52.280 3210.435 ;
        RECT 16.660 3056.270 16.920 3056.590 ;
        RECT 52.080 3056.270 52.340 3056.590 ;
        RECT 16.720 3052.365 16.860 3056.270 ;
        RECT 16.650 3051.995 16.930 3052.365 ;
      LAYER via2 ;
        RECT 1846.990 3216.600 1847.270 3216.880 ;
        RECT 52.070 3210.480 52.350 3210.760 ;
        RECT 16.650 3052.040 16.930 3052.320 ;
      LAYER met3 ;
        RECT 1846.965 3216.900 1847.295 3216.905 ;
        RECT 1846.710 3216.890 1847.295 3216.900 ;
        RECT 1846.510 3216.590 1847.295 3216.890 ;
        RECT 1846.710 3216.580 1847.295 3216.590 ;
        RECT 1846.965 3216.575 1847.295 3216.580 ;
        RECT 52.045 3210.770 52.375 3210.785 ;
        RECT 1846.710 3210.770 1847.090 3210.780 ;
        RECT 52.045 3210.470 1847.090 3210.770 ;
        RECT 52.045 3210.455 52.375 3210.470 ;
        RECT 1846.710 3210.460 1847.090 3210.470 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 16.625 3052.330 16.955 3052.345 ;
        RECT -4.800 3052.030 16.955 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 16.625 3052.015 16.955 3052.030 ;
      LAYER via3 ;
        RECT 1846.740 3216.580 1847.060 3216.900 ;
        RECT 1846.740 3210.460 1847.060 3210.780 ;
      LAYER met4 ;
        RECT 1846.735 3216.575 1847.065 3216.905 ;
        RECT 1846.750 3210.785 1847.050 3216.575 ;
        RECT 1846.735 3210.455 1847.065 3210.785 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 25.370 3234.320 25.690 3234.380 ;
        RECT 1911.830 3234.320 1912.150 3234.380 ;
        RECT 25.370 3234.180 1912.150 3234.320 ;
        RECT 25.370 3234.120 25.690 3234.180 ;
        RECT 1911.830 3234.120 1912.150 3234.180 ;
        RECT 13.870 2765.460 14.190 2765.520 ;
        RECT 25.370 2765.460 25.690 2765.520 ;
        RECT 13.870 2765.320 25.690 2765.460 ;
        RECT 13.870 2765.260 14.190 2765.320 ;
        RECT 25.370 2765.260 25.690 2765.320 ;
      LAYER via ;
        RECT 25.400 3234.120 25.660 3234.380 ;
        RECT 1911.860 3234.120 1912.120 3234.380 ;
        RECT 13.900 2765.260 14.160 2765.520 ;
        RECT 25.400 2765.260 25.660 2765.520 ;
      LAYER met2 ;
        RECT 25.400 3234.090 25.660 3234.410 ;
        RECT 1911.860 3234.090 1912.120 3234.410 ;
        RECT 25.460 2765.550 25.600 3234.090 ;
        RECT 1911.920 3220.000 1912.060 3234.090 ;
        RECT 1911.900 3216.000 1912.180 3220.000 ;
        RECT 13.900 2765.405 14.160 2765.550 ;
        RECT 13.890 2765.035 14.170 2765.405 ;
        RECT 25.400 2765.230 25.660 2765.550 ;
      LAYER via2 ;
        RECT 13.890 2765.080 14.170 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 13.865 2765.370 14.195 2765.385 ;
        RECT -4.800 2765.070 14.195 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 13.865 2765.055 14.195 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2477.820 16.950 2477.880 ;
        RECT 44.230 2477.820 44.550 2477.880 ;
        RECT 16.630 2477.680 44.550 2477.820 ;
        RECT 16.630 2477.620 16.950 2477.680 ;
        RECT 44.230 2477.620 44.550 2477.680 ;
      LAYER via ;
        RECT 16.660 2477.620 16.920 2477.880 ;
        RECT 44.260 2477.620 44.520 2477.880 ;
      LAYER met2 ;
        RECT 1973.950 3216.810 1974.230 3216.925 ;
        RECT 1974.920 3216.810 1975.200 3220.000 ;
        RECT 1973.950 3216.670 1975.200 3216.810 ;
        RECT 1973.950 3216.555 1974.230 3216.670 ;
        RECT 1974.920 3216.000 1975.200 3216.670 ;
        RECT 44.250 3208.395 44.530 3208.765 ;
        RECT 44.320 2477.910 44.460 3208.395 ;
        RECT 16.660 2477.765 16.920 2477.910 ;
        RECT 16.650 2477.395 16.930 2477.765 ;
        RECT 44.260 2477.590 44.520 2477.910 ;
      LAYER via2 ;
        RECT 1973.950 3216.600 1974.230 3216.880 ;
        RECT 44.250 3208.440 44.530 3208.720 ;
        RECT 16.650 2477.440 16.930 2477.720 ;
      LAYER met3 ;
        RECT 1973.925 3216.900 1974.255 3216.905 ;
        RECT 1973.670 3216.890 1974.255 3216.900 ;
        RECT 1973.470 3216.590 1974.255 3216.890 ;
        RECT 1973.670 3216.580 1974.255 3216.590 ;
        RECT 1973.925 3216.575 1974.255 3216.580 ;
        RECT 44.225 3208.730 44.555 3208.745 ;
        RECT 1973.670 3208.730 1974.050 3208.740 ;
        RECT 44.225 3208.430 1974.050 3208.730 ;
        RECT 44.225 3208.415 44.555 3208.430 ;
        RECT 1973.670 3208.420 1974.050 3208.430 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 16.625 2477.730 16.955 2477.745 ;
        RECT -4.800 2477.430 16.955 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 16.625 2477.415 16.955 2477.430 ;
      LAYER via3 ;
        RECT 1973.700 3216.580 1974.020 3216.900 ;
        RECT 1973.700 3208.420 1974.020 3208.740 ;
      LAYER met4 ;
        RECT 1973.695 3216.575 1974.025 3216.905 ;
        RECT 1973.710 3208.745 1974.010 3216.575 ;
        RECT 1973.695 3208.415 1974.025 3208.745 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 959.170 3235.680 959.490 3235.740 ;
        RECT 2037.870 3235.680 2038.190 3235.740 ;
        RECT 959.170 3235.540 2038.190 3235.680 ;
        RECT 959.170 3235.480 959.490 3235.540 ;
        RECT 2037.870 3235.480 2038.190 3235.540 ;
        RECT 19.390 3221.740 19.710 3221.800 ;
        RECT 959.170 3221.740 959.490 3221.800 ;
        RECT 19.390 3221.600 959.490 3221.740 ;
        RECT 19.390 3221.540 19.710 3221.600 ;
        RECT 959.170 3221.540 959.490 3221.600 ;
      LAYER via ;
        RECT 959.200 3235.480 959.460 3235.740 ;
        RECT 2037.900 3235.480 2038.160 3235.740 ;
        RECT 19.420 3221.540 19.680 3221.800 ;
        RECT 959.200 3221.540 959.460 3221.800 ;
      LAYER met2 ;
        RECT 959.200 3235.450 959.460 3235.770 ;
        RECT 2037.900 3235.450 2038.160 3235.770 ;
        RECT 959.260 3221.830 959.400 3235.450 ;
        RECT 19.420 3221.510 19.680 3221.830 ;
        RECT 959.200 3221.510 959.460 3221.830 ;
        RECT 19.480 2190.125 19.620 3221.510 ;
        RECT 2037.960 3220.000 2038.100 3235.450 ;
        RECT 2037.940 3216.000 2038.220 3220.000 ;
        RECT 19.410 2189.755 19.690 2190.125 ;
      LAYER via2 ;
        RECT 19.410 2189.800 19.690 2190.080 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 19.385 2190.090 19.715 2190.105 ;
        RECT -4.800 2189.790 19.715 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 19.385 2189.775 19.715 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.930 3218.000 19.250 3218.060 ;
        RECT 2099.510 3218.000 2099.830 3218.060 ;
        RECT 18.930 3217.860 2099.830 3218.000 ;
        RECT 18.930 3217.800 19.250 3217.860 ;
        RECT 2099.510 3217.800 2099.830 3217.860 ;
      LAYER via ;
        RECT 18.960 3217.800 19.220 3218.060 ;
        RECT 2099.540 3217.800 2099.800 3218.060 ;
      LAYER met2 ;
        RECT 2100.960 3218.170 2101.240 3220.000 ;
        RECT 2099.600 3218.090 2101.240 3218.170 ;
        RECT 18.960 3217.770 19.220 3218.090 ;
        RECT 2099.540 3218.030 2101.240 3218.090 ;
        RECT 2099.540 3217.770 2099.800 3218.030 ;
        RECT 19.020 1903.165 19.160 3217.770 ;
        RECT 2100.960 3216.000 2101.240 3218.030 ;
        RECT 18.950 1902.795 19.230 1903.165 ;
      LAYER via2 ;
        RECT 18.950 1902.840 19.230 1903.120 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 18.925 1903.130 19.255 1903.145 ;
        RECT -4.800 1902.830 19.255 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 18.925 1902.815 19.255 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 398.045 3215.465 398.215 3216.995 ;
      LAYER mcon ;
        RECT 398.045 3216.825 398.215 3216.995 ;
      LAYER met1 ;
        RECT 397.970 3216.980 398.290 3217.040 ;
        RECT 397.775 3216.840 398.290 3216.980 ;
        RECT 397.970 3216.780 398.290 3216.840 ;
        RECT 397.985 3215.620 398.275 3215.665 ;
        RECT 2902.210 3215.620 2902.530 3215.680 ;
        RECT 397.985 3215.480 2902.530 3215.620 ;
        RECT 397.985 3215.435 398.275 3215.480 ;
        RECT 2902.210 3215.420 2902.530 3215.480 ;
      LAYER via ;
        RECT 398.000 3216.780 398.260 3217.040 ;
        RECT 2902.240 3215.420 2902.500 3215.680 ;
      LAYER met2 ;
        RECT 396.200 3216.810 396.480 3220.000 ;
        RECT 398.000 3216.810 398.260 3217.070 ;
        RECT 396.200 3216.750 398.260 3216.810 ;
        RECT 396.200 3216.670 398.200 3216.750 ;
        RECT 396.200 3216.000 396.480 3216.670 ;
        RECT 2902.240 3215.390 2902.500 3215.710 ;
        RECT 2902.300 615.925 2902.440 3215.390 ;
        RECT 2902.230 615.555 2902.510 615.925 ;
      LAYER via2 ;
        RECT 2902.230 615.600 2902.510 615.880 ;
      LAYER met3 ;
        RECT 2902.205 615.890 2902.535 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2902.205 615.590 2924.800 615.890 ;
        RECT 2902.205 615.575 2902.535 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 3232.620 18.330 3232.680 ;
        RECT 2164.370 3232.620 2164.690 3232.680 ;
        RECT 18.010 3232.480 2164.690 3232.620 ;
        RECT 18.010 3232.420 18.330 3232.480 ;
        RECT 2164.370 3232.420 2164.690 3232.480 ;
      LAYER via ;
        RECT 18.040 3232.420 18.300 3232.680 ;
        RECT 2164.400 3232.420 2164.660 3232.680 ;
      LAYER met2 ;
        RECT 18.040 3232.390 18.300 3232.710 ;
        RECT 2164.400 3232.390 2164.660 3232.710 ;
        RECT 18.100 1615.525 18.240 3232.390 ;
        RECT 2164.460 3220.000 2164.600 3232.390 ;
        RECT 2164.440 3216.000 2164.720 3220.000 ;
        RECT 18.030 1615.155 18.310 1615.525 ;
      LAYER via2 ;
        RECT 18.030 1615.200 18.310 1615.480 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 18.005 1615.490 18.335 1615.505 ;
        RECT -4.800 1615.190 18.335 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 18.005 1615.175 18.335 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 32.270 3231.940 32.590 3232.000 ;
        RECT 2227.390 3231.940 2227.710 3232.000 ;
        RECT 32.270 3231.800 2227.710 3231.940 ;
        RECT 32.270 3231.740 32.590 3231.800 ;
        RECT 2227.390 3231.740 2227.710 3231.800 ;
        RECT 16.170 1400.700 16.490 1400.760 ;
        RECT 32.270 1400.700 32.590 1400.760 ;
        RECT 16.170 1400.560 32.590 1400.700 ;
        RECT 16.170 1400.500 16.490 1400.560 ;
        RECT 32.270 1400.500 32.590 1400.560 ;
      LAYER via ;
        RECT 32.300 3231.740 32.560 3232.000 ;
        RECT 2227.420 3231.740 2227.680 3232.000 ;
        RECT 16.200 1400.500 16.460 1400.760 ;
        RECT 32.300 1400.500 32.560 1400.760 ;
      LAYER met2 ;
        RECT 32.300 3231.710 32.560 3232.030 ;
        RECT 2227.420 3231.710 2227.680 3232.030 ;
        RECT 32.360 1400.790 32.500 3231.710 ;
        RECT 2227.480 3220.000 2227.620 3231.710 ;
        RECT 2227.460 3216.000 2227.740 3220.000 ;
        RECT 16.200 1400.645 16.460 1400.790 ;
        RECT 16.190 1400.275 16.470 1400.645 ;
        RECT 32.300 1400.470 32.560 1400.790 ;
      LAYER via2 ;
        RECT 16.190 1400.320 16.470 1400.600 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 16.165 1400.610 16.495 1400.625 ;
        RECT -4.800 1400.310 16.495 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 16.165 1400.295 16.495 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 31.350 3231.600 31.670 3231.660 ;
        RECT 2290.410 3231.600 2290.730 3231.660 ;
        RECT 31.350 3231.460 2290.730 3231.600 ;
        RECT 31.350 3231.400 31.670 3231.460 ;
        RECT 2290.410 3231.400 2290.730 3231.460 ;
        RECT 15.710 1185.480 16.030 1185.540 ;
        RECT 31.350 1185.480 31.670 1185.540 ;
        RECT 15.710 1185.340 31.670 1185.480 ;
        RECT 15.710 1185.280 16.030 1185.340 ;
        RECT 31.350 1185.280 31.670 1185.340 ;
      LAYER via ;
        RECT 31.380 3231.400 31.640 3231.660 ;
        RECT 2290.440 3231.400 2290.700 3231.660 ;
        RECT 15.740 1185.280 16.000 1185.540 ;
        RECT 31.380 1185.280 31.640 1185.540 ;
      LAYER met2 ;
        RECT 31.380 3231.370 31.640 3231.690 ;
        RECT 2290.440 3231.370 2290.700 3231.690 ;
        RECT 31.440 1185.570 31.580 3231.370 ;
        RECT 2290.500 3220.000 2290.640 3231.370 ;
        RECT 2290.480 3216.000 2290.760 3220.000 ;
        RECT 15.740 1185.250 16.000 1185.570 ;
        RECT 31.380 1185.250 31.640 1185.570 ;
        RECT 15.800 1185.085 15.940 1185.250 ;
        RECT 15.730 1184.715 16.010 1185.085 ;
      LAYER via2 ;
        RECT 15.730 1184.760 16.010 1185.040 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 15.705 1185.050 16.035 1185.065 ;
        RECT -4.800 1184.750 16.035 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 15.705 1184.735 16.035 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 30.890 3230.920 31.210 3230.980 ;
        RECT 2353.890 3230.920 2354.210 3230.980 ;
        RECT 30.890 3230.780 2354.210 3230.920 ;
        RECT 30.890 3230.720 31.210 3230.780 ;
        RECT 2353.890 3230.720 2354.210 3230.780 ;
        RECT 15.250 969.920 15.570 969.980 ;
        RECT 30.890 969.920 31.210 969.980 ;
        RECT 15.250 969.780 31.210 969.920 ;
        RECT 15.250 969.720 15.570 969.780 ;
        RECT 30.890 969.720 31.210 969.780 ;
      LAYER via ;
        RECT 30.920 3230.720 31.180 3230.980 ;
        RECT 2353.920 3230.720 2354.180 3230.980 ;
        RECT 15.280 969.720 15.540 969.980 ;
        RECT 30.920 969.720 31.180 969.980 ;
      LAYER met2 ;
        RECT 30.920 3230.690 31.180 3231.010 ;
        RECT 2353.920 3230.690 2354.180 3231.010 ;
        RECT 30.980 970.010 31.120 3230.690 ;
        RECT 2353.980 3220.000 2354.120 3230.690 ;
        RECT 2353.960 3216.000 2354.240 3220.000 ;
        RECT 15.280 969.690 15.540 970.010 ;
        RECT 30.920 969.690 31.180 970.010 ;
        RECT 15.340 969.525 15.480 969.690 ;
        RECT 15.270 969.155 15.550 969.525 ;
      LAYER via2 ;
        RECT 15.270 969.200 15.550 969.480 ;
      LAYER met3 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 15.245 969.490 15.575 969.505 ;
        RECT -4.800 969.190 15.575 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 15.245 969.175 15.575 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 51.590 3230.580 51.910 3230.640 ;
        RECT 2416.910 3230.580 2417.230 3230.640 ;
        RECT 51.590 3230.440 2417.230 3230.580 ;
        RECT 51.590 3230.380 51.910 3230.440 ;
        RECT 2416.910 3230.380 2417.230 3230.440 ;
        RECT 16.630 758.780 16.950 758.840 ;
        RECT 51.590 758.780 51.910 758.840 ;
        RECT 16.630 758.640 51.910 758.780 ;
        RECT 16.630 758.580 16.950 758.640 ;
        RECT 51.590 758.580 51.910 758.640 ;
      LAYER via ;
        RECT 51.620 3230.380 51.880 3230.640 ;
        RECT 2416.940 3230.380 2417.200 3230.640 ;
        RECT 16.660 758.580 16.920 758.840 ;
        RECT 51.620 758.580 51.880 758.840 ;
      LAYER met2 ;
        RECT 51.620 3230.350 51.880 3230.670 ;
        RECT 2416.940 3230.350 2417.200 3230.670 ;
        RECT 51.680 758.870 51.820 3230.350 ;
        RECT 2417.000 3220.000 2417.140 3230.350 ;
        RECT 2416.980 3216.000 2417.260 3220.000 ;
        RECT 16.660 758.550 16.920 758.870 ;
        RECT 51.620 758.550 51.880 758.870 ;
        RECT 16.720 753.965 16.860 758.550 ;
        RECT 16.650 753.595 16.930 753.965 ;
      LAYER via2 ;
        RECT 16.650 753.640 16.930 753.920 ;
      LAYER met3 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 16.625 753.930 16.955 753.945 ;
        RECT -4.800 753.630 16.955 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 16.625 753.615 16.955 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 65.390 3230.240 65.710 3230.300 ;
        RECT 2479.930 3230.240 2480.250 3230.300 ;
        RECT 65.390 3230.100 2480.250 3230.240 ;
        RECT 65.390 3230.040 65.710 3230.100 ;
        RECT 2479.930 3230.040 2480.250 3230.100 ;
        RECT 16.170 544.920 16.490 544.980 ;
        RECT 65.390 544.920 65.710 544.980 ;
        RECT 16.170 544.780 65.710 544.920 ;
        RECT 16.170 544.720 16.490 544.780 ;
        RECT 65.390 544.720 65.710 544.780 ;
      LAYER via ;
        RECT 65.420 3230.040 65.680 3230.300 ;
        RECT 2479.960 3230.040 2480.220 3230.300 ;
        RECT 16.200 544.720 16.460 544.980 ;
        RECT 65.420 544.720 65.680 544.980 ;
      LAYER met2 ;
        RECT 65.420 3230.010 65.680 3230.330 ;
        RECT 2479.960 3230.010 2480.220 3230.330 ;
        RECT 65.480 545.010 65.620 3230.010 ;
        RECT 2480.020 3220.000 2480.160 3230.010 ;
        RECT 2480.000 3216.000 2480.280 3220.000 ;
        RECT 16.200 544.690 16.460 545.010 ;
        RECT 65.420 544.690 65.680 545.010 ;
        RECT 16.260 538.405 16.400 544.690 ;
        RECT 16.190 538.035 16.470 538.405 ;
      LAYER via2 ;
        RECT 16.190 538.080 16.470 538.360 ;
      LAYER met3 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 16.165 538.370 16.495 538.385 ;
        RECT -4.800 538.070 16.495 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 16.165 538.055 16.495 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 72.290 3229.560 72.610 3229.620 ;
        RECT 2542.950 3229.560 2543.270 3229.620 ;
        RECT 72.290 3229.420 2543.270 3229.560 ;
        RECT 72.290 3229.360 72.610 3229.420 ;
        RECT 2542.950 3229.360 2543.270 3229.420 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 72.290 324.260 72.610 324.320 ;
        RECT 16.630 324.120 72.610 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 72.290 324.060 72.610 324.120 ;
      LAYER via ;
        RECT 72.320 3229.360 72.580 3229.620 ;
        RECT 2542.980 3229.360 2543.240 3229.620 ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 72.320 324.060 72.580 324.320 ;
      LAYER met2 ;
        RECT 72.320 3229.330 72.580 3229.650 ;
        RECT 2542.980 3229.330 2543.240 3229.650 ;
        RECT 72.380 324.350 72.520 3229.330 ;
        RECT 2543.040 3220.000 2543.180 3229.330 ;
        RECT 2543.020 3216.000 2543.300 3220.000 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 72.320 324.030 72.580 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2604.610 3216.810 2604.890 3216.925 ;
        RECT 2606.500 3216.810 2606.780 3220.000 ;
        RECT 2604.610 3216.670 2606.780 3216.810 ;
        RECT 2604.610 3216.555 2604.890 3216.670 ;
        RECT 2606.500 3216.000 2606.780 3216.670 ;
      LAYER via2 ;
        RECT 2604.610 3216.600 2604.890 3216.880 ;
      LAYER met3 ;
        RECT 2590.070 3216.890 2590.450 3216.900 ;
        RECT 2604.585 3216.890 2604.915 3216.905 ;
        RECT 2590.070 3216.590 2604.915 3216.890 ;
        RECT 2590.070 3216.580 2590.450 3216.590 ;
        RECT 2604.585 3216.575 2604.915 3216.590 ;
        RECT 2590.070 109.970 2590.450 109.980 ;
        RECT 3.070 109.670 2590.450 109.970 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 3.070 107.250 3.370 109.670 ;
        RECT 2590.070 109.660 2590.450 109.670 ;
        RECT -4.800 106.950 3.370 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
      LAYER via3 ;
        RECT 2590.100 3216.580 2590.420 3216.900 ;
        RECT 2590.100 109.660 2590.420 109.980 ;
      LAYER met4 ;
        RECT 2590.095 3216.575 2590.425 3216.905 ;
        RECT 2590.110 109.985 2590.410 3216.575 ;
        RECT 2590.095 109.655 2590.425 109.985 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 460.530 3217.320 460.850 3217.380 ;
        RECT 2625.290 3217.320 2625.610 3217.380 ;
        RECT 460.530 3217.180 2625.610 3217.320 ;
        RECT 460.530 3217.120 460.850 3217.180 ;
        RECT 2625.290 3217.120 2625.610 3217.180 ;
        RECT 2625.290 855.340 2625.610 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 2625.290 855.200 2901.150 855.340 ;
        RECT 2625.290 855.140 2625.610 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 460.560 3217.120 460.820 3217.380 ;
        RECT 2625.320 3217.120 2625.580 3217.380 ;
        RECT 2625.320 855.140 2625.580 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 459.220 3217.490 459.500 3220.000 ;
        RECT 459.220 3217.410 460.760 3217.490 ;
        RECT 459.220 3217.350 460.820 3217.410 ;
        RECT 459.220 3216.000 459.500 3217.350 ;
        RECT 460.560 3217.090 460.820 3217.350 ;
        RECT 2625.320 3217.090 2625.580 3217.410 ;
        RECT 2625.380 855.430 2625.520 3217.090 ;
        RECT 2625.320 855.110 2625.580 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 522.170 3233.640 522.490 3233.700 ;
        RECT 700.190 3233.640 700.510 3233.700 ;
        RECT 522.170 3233.500 700.510 3233.640 ;
        RECT 522.170 3233.440 522.490 3233.500 ;
        RECT 700.190 3233.440 700.510 3233.500 ;
        RECT 700.190 3219.700 700.510 3219.760 ;
        RECT 2902.670 3219.700 2902.990 3219.760 ;
        RECT 700.190 3219.560 2902.990 3219.700 ;
        RECT 700.190 3219.500 700.510 3219.560 ;
        RECT 2902.670 3219.500 2902.990 3219.560 ;
      LAYER via ;
        RECT 522.200 3233.440 522.460 3233.700 ;
        RECT 700.220 3233.440 700.480 3233.700 ;
        RECT 700.220 3219.500 700.480 3219.760 ;
        RECT 2902.700 3219.500 2902.960 3219.760 ;
      LAYER met2 ;
        RECT 522.200 3233.410 522.460 3233.730 ;
        RECT 700.220 3233.410 700.480 3233.730 ;
        RECT 522.260 3220.000 522.400 3233.410 ;
        RECT 522.240 3216.000 522.520 3220.000 ;
        RECT 700.280 3219.790 700.420 3233.410 ;
        RECT 700.220 3219.470 700.480 3219.790 ;
        RECT 2902.700 3219.470 2902.960 3219.790 ;
        RECT 2902.760 1085.125 2902.900 3219.470 ;
        RECT 2902.690 1084.755 2902.970 1085.125 ;
      LAYER via2 ;
        RECT 2902.690 1084.800 2902.970 1085.080 ;
      LAYER met3 ;
        RECT 2902.665 1085.090 2902.995 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2902.665 1084.790 2924.800 1085.090 ;
        RECT 2902.665 1084.775 2902.995 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 586.185 3216.145 586.355 3218.355 ;
      LAYER mcon ;
        RECT 586.185 3218.185 586.355 3218.355 ;
      LAYER met1 ;
        RECT 586.110 3218.340 586.430 3218.400 ;
        RECT 585.915 3218.200 586.430 3218.340 ;
        RECT 586.110 3218.140 586.430 3218.200 ;
        RECT 586.125 3216.300 586.415 3216.345 ;
        RECT 2903.130 3216.300 2903.450 3216.360 ;
        RECT 586.125 3216.160 2903.450 3216.300 ;
        RECT 586.125 3216.115 586.415 3216.160 ;
        RECT 2903.130 3216.100 2903.450 3216.160 ;
      LAYER via ;
        RECT 586.140 3218.140 586.400 3218.400 ;
        RECT 2903.160 3216.100 2903.420 3216.360 ;
      LAYER met2 ;
        RECT 585.260 3218.170 585.540 3220.000 ;
        RECT 586.140 3218.170 586.400 3218.430 ;
        RECT 585.260 3218.110 586.400 3218.170 ;
        RECT 585.260 3218.030 586.340 3218.110 ;
        RECT 585.260 3216.000 585.540 3218.030 ;
        RECT 2903.160 3216.070 2903.420 3216.390 ;
        RECT 2903.220 1319.725 2903.360 3216.070 ;
        RECT 2903.150 1319.355 2903.430 1319.725 ;
      LAYER via2 ;
        RECT 2903.150 1319.400 2903.430 1319.680 ;
      LAYER met3 ;
        RECT 2903.125 1319.690 2903.455 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2903.125 1319.390 2924.800 1319.690 ;
        RECT 2903.125 1319.375 2903.455 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 648.670 3232.960 648.990 3233.020 ;
        RECT 2626.210 3232.960 2626.530 3233.020 ;
        RECT 648.670 3232.820 2626.530 3232.960 ;
        RECT 648.670 3232.760 648.990 3232.820 ;
        RECT 2626.210 3232.760 2626.530 3232.820 ;
        RECT 2626.210 1559.140 2626.530 1559.200 ;
        RECT 2900.830 1559.140 2901.150 1559.200 ;
        RECT 2626.210 1559.000 2901.150 1559.140 ;
        RECT 2626.210 1558.940 2626.530 1559.000 ;
        RECT 2900.830 1558.940 2901.150 1559.000 ;
      LAYER via ;
        RECT 648.700 3232.760 648.960 3233.020 ;
        RECT 2626.240 3232.760 2626.500 3233.020 ;
        RECT 2626.240 1558.940 2626.500 1559.200 ;
        RECT 2900.860 1558.940 2901.120 1559.200 ;
      LAYER met2 ;
        RECT 648.700 3232.730 648.960 3233.050 ;
        RECT 2626.240 3232.730 2626.500 3233.050 ;
        RECT 648.760 3220.000 648.900 3232.730 ;
        RECT 648.740 3216.000 649.020 3220.000 ;
        RECT 2626.300 1559.230 2626.440 3232.730 ;
        RECT 2626.240 1558.910 2626.500 1559.230 ;
        RECT 2900.860 1558.910 2901.120 1559.230 ;
        RECT 2900.920 1554.325 2901.060 1558.910 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
      LAYER via2 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
      LAYER met3 ;
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 711.690 3233.640 712.010 3233.700 ;
        RECT 2626.670 3233.640 2626.990 3233.700 ;
        RECT 711.690 3233.500 2626.990 3233.640 ;
        RECT 711.690 3233.440 712.010 3233.500 ;
        RECT 2626.670 3233.440 2626.990 3233.500 ;
        RECT 2626.670 1793.740 2626.990 1793.800 ;
        RECT 2899.910 1793.740 2900.230 1793.800 ;
        RECT 2626.670 1793.600 2900.230 1793.740 ;
        RECT 2626.670 1793.540 2626.990 1793.600 ;
        RECT 2899.910 1793.540 2900.230 1793.600 ;
      LAYER via ;
        RECT 711.720 3233.440 711.980 3233.700 ;
        RECT 2626.700 3233.440 2626.960 3233.700 ;
        RECT 2626.700 1793.540 2626.960 1793.800 ;
        RECT 2899.940 1793.540 2900.200 1793.800 ;
      LAYER met2 ;
        RECT 711.720 3233.410 711.980 3233.730 ;
        RECT 2626.700 3233.410 2626.960 3233.730 ;
        RECT 711.780 3220.000 711.920 3233.410 ;
        RECT 711.760 3216.000 712.040 3220.000 ;
        RECT 2626.760 1793.830 2626.900 3233.410 ;
        RECT 2626.700 1793.510 2626.960 1793.830 ;
        RECT 2899.940 1793.510 2900.200 1793.830 ;
        RECT 2900.000 1789.605 2900.140 1793.510 ;
        RECT 2899.930 1789.235 2900.210 1789.605 ;
      LAYER via2 ;
        RECT 2899.930 1789.280 2900.210 1789.560 ;
      LAYER met3 ;
        RECT 2899.905 1789.570 2900.235 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2899.905 1789.270 2924.800 1789.570 ;
        RECT 2899.905 1789.255 2900.235 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 774.710 3233.980 775.030 3234.040 ;
        RECT 2687.390 3233.980 2687.710 3234.040 ;
        RECT 774.710 3233.840 2687.710 3233.980 ;
        RECT 774.710 3233.780 775.030 3233.840 ;
        RECT 2687.390 3233.780 2687.710 3233.840 ;
        RECT 2687.390 2028.340 2687.710 2028.400 ;
        RECT 2899.910 2028.340 2900.230 2028.400 ;
        RECT 2687.390 2028.200 2900.230 2028.340 ;
        RECT 2687.390 2028.140 2687.710 2028.200 ;
        RECT 2899.910 2028.140 2900.230 2028.200 ;
      LAYER via ;
        RECT 774.740 3233.780 775.000 3234.040 ;
        RECT 2687.420 3233.780 2687.680 3234.040 ;
        RECT 2687.420 2028.140 2687.680 2028.400 ;
        RECT 2899.940 2028.140 2900.200 2028.400 ;
      LAYER met2 ;
        RECT 774.740 3233.750 775.000 3234.070 ;
        RECT 2687.420 3233.750 2687.680 3234.070 ;
        RECT 774.800 3220.000 774.940 3233.750 ;
        RECT 774.780 3216.000 775.060 3220.000 ;
        RECT 2687.480 2028.430 2687.620 3233.750 ;
        RECT 2687.420 2028.110 2687.680 2028.430 ;
        RECT 2899.940 2028.110 2900.200 2028.430 ;
        RECT 2900.000 2024.205 2900.140 2028.110 ;
        RECT 2899.930 2023.835 2900.210 2024.205 ;
      LAYER via2 ;
        RECT 2899.930 2023.880 2900.210 2024.160 ;
      LAYER met3 ;
        RECT 2899.905 2024.170 2900.235 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2899.905 2023.870 2924.800 2024.170 ;
        RECT 2899.905 2023.855 2900.235 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 838.190 3235.340 838.510 3235.400 ;
        RECT 2613.330 3235.340 2613.650 3235.400 ;
        RECT 838.190 3235.200 2613.650 3235.340 ;
        RECT 838.190 3235.140 838.510 3235.200 ;
        RECT 2613.330 3235.140 2613.650 3235.200 ;
        RECT 2613.330 2262.940 2613.650 2263.000 ;
        RECT 2899.910 2262.940 2900.230 2263.000 ;
        RECT 2613.330 2262.800 2900.230 2262.940 ;
        RECT 2613.330 2262.740 2613.650 2262.800 ;
        RECT 2899.910 2262.740 2900.230 2262.800 ;
      LAYER via ;
        RECT 838.220 3235.140 838.480 3235.400 ;
        RECT 2613.360 3235.140 2613.620 3235.400 ;
        RECT 2613.360 2262.740 2613.620 2263.000 ;
        RECT 2899.940 2262.740 2900.200 2263.000 ;
      LAYER met2 ;
        RECT 838.220 3235.110 838.480 3235.430 ;
        RECT 2613.360 3235.110 2613.620 3235.430 ;
        RECT 838.280 3220.000 838.420 3235.110 ;
        RECT 838.260 3216.000 838.540 3220.000 ;
        RECT 2613.420 2263.030 2613.560 3235.110 ;
        RECT 2613.360 2262.710 2613.620 2263.030 ;
        RECT 2899.940 2262.710 2900.200 2263.030 ;
        RECT 2900.000 2258.805 2900.140 2262.710 ;
        RECT 2899.930 2258.435 2900.210 2258.805 ;
      LAYER via2 ;
        RECT 2899.930 2258.480 2900.210 2258.760 ;
      LAYER met3 ;
        RECT 2899.905 2258.770 2900.235 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2899.905 2258.470 2924.800 2258.770 ;
        RECT 2899.905 2258.455 2900.235 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 633.030 17.240 633.350 17.300 ;
        RECT 738.830 17.240 739.150 17.300 ;
        RECT 633.030 17.100 739.150 17.240 ;
        RECT 633.030 17.040 633.350 17.100 ;
        RECT 738.830 17.040 739.150 17.100 ;
      LAYER via ;
        RECT 633.060 17.040 633.320 17.300 ;
        RECT 738.860 17.040 739.120 17.300 ;
      LAYER met2 ;
        RECT 738.900 220.000 739.180 224.000 ;
        RECT 738.920 17.330 739.060 220.000 ;
        RECT 633.060 17.010 633.320 17.330 ;
        RECT 738.860 17.010 739.120 17.330 ;
        RECT 633.120 2.400 633.260 17.010 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2208.070 207.300 2208.390 207.360 ;
        RECT 2214.050 207.300 2214.370 207.360 ;
        RECT 2208.070 207.160 2214.370 207.300 ;
        RECT 2208.070 207.100 2208.390 207.160 ;
        RECT 2214.050 207.100 2214.370 207.160 ;
        RECT 2214.050 25.740 2214.370 25.800 ;
        RECT 2417.370 25.740 2417.690 25.800 ;
        RECT 2214.050 25.600 2417.690 25.740 ;
        RECT 2214.050 25.540 2214.370 25.600 ;
        RECT 2417.370 25.540 2417.690 25.600 ;
      LAYER via ;
        RECT 2208.100 207.100 2208.360 207.360 ;
        RECT 2214.080 207.100 2214.340 207.360 ;
        RECT 2214.080 25.540 2214.340 25.800 ;
        RECT 2417.400 25.540 2417.660 25.800 ;
      LAYER met2 ;
        RECT 2208.140 220.000 2208.420 224.000 ;
        RECT 2208.160 207.390 2208.300 220.000 ;
        RECT 2208.100 207.070 2208.360 207.390 ;
        RECT 2214.080 207.070 2214.340 207.390 ;
        RECT 2214.140 25.830 2214.280 207.070 ;
        RECT 2214.080 25.510 2214.340 25.830 ;
        RECT 2417.400 25.510 2417.660 25.830 ;
        RECT 2417.460 2.400 2417.600 25.510 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2222.790 207.300 2223.110 207.360 ;
        RECT 2228.310 207.300 2228.630 207.360 ;
        RECT 2222.790 207.160 2228.630 207.300 ;
        RECT 2222.790 207.100 2223.110 207.160 ;
        RECT 2228.310 207.100 2228.630 207.160 ;
        RECT 2228.310 26.080 2228.630 26.140 ;
        RECT 2434.850 26.080 2435.170 26.140 ;
        RECT 2228.310 25.940 2435.170 26.080 ;
        RECT 2228.310 25.880 2228.630 25.940 ;
        RECT 2434.850 25.880 2435.170 25.940 ;
      LAYER via ;
        RECT 2222.820 207.100 2223.080 207.360 ;
        RECT 2228.340 207.100 2228.600 207.360 ;
        RECT 2228.340 25.880 2228.600 26.140 ;
        RECT 2434.880 25.880 2435.140 26.140 ;
      LAYER met2 ;
        RECT 2222.860 220.000 2223.140 224.000 ;
        RECT 2222.880 207.390 2223.020 220.000 ;
        RECT 2222.820 207.070 2223.080 207.390 ;
        RECT 2228.340 207.070 2228.600 207.390 ;
        RECT 2228.400 26.170 2228.540 207.070 ;
        RECT 2228.340 25.850 2228.600 26.170 ;
        RECT 2434.880 25.850 2435.140 26.170 ;
        RECT 2434.940 2.400 2435.080 25.850 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2237.510 207.300 2237.830 207.360 ;
        RECT 2242.110 207.300 2242.430 207.360 ;
        RECT 2237.510 207.160 2242.430 207.300 ;
        RECT 2237.510 207.100 2237.830 207.160 ;
        RECT 2242.110 207.100 2242.430 207.160 ;
        RECT 2242.110 25.400 2242.430 25.460 ;
        RECT 2452.790 25.400 2453.110 25.460 ;
        RECT 2242.110 25.260 2453.110 25.400 ;
        RECT 2242.110 25.200 2242.430 25.260 ;
        RECT 2452.790 25.200 2453.110 25.260 ;
      LAYER via ;
        RECT 2237.540 207.100 2237.800 207.360 ;
        RECT 2242.140 207.100 2242.400 207.360 ;
        RECT 2242.140 25.200 2242.400 25.460 ;
        RECT 2452.820 25.200 2453.080 25.460 ;
      LAYER met2 ;
        RECT 2237.580 220.000 2237.860 224.000 ;
        RECT 2237.600 207.390 2237.740 220.000 ;
        RECT 2237.540 207.070 2237.800 207.390 ;
        RECT 2242.140 207.070 2242.400 207.390 ;
        RECT 2242.200 25.490 2242.340 207.070 ;
        RECT 2242.140 25.170 2242.400 25.490 ;
        RECT 2452.820 25.170 2453.080 25.490 ;
        RECT 2452.880 2.400 2453.020 25.170 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2252.230 207.300 2252.550 207.360 ;
        RECT 2255.910 207.300 2256.230 207.360 ;
        RECT 2252.230 207.160 2256.230 207.300 ;
        RECT 2252.230 207.100 2252.550 207.160 ;
        RECT 2255.910 207.100 2256.230 207.160 ;
        RECT 2255.910 24.380 2256.230 24.440 ;
        RECT 2470.730 24.380 2471.050 24.440 ;
        RECT 2255.910 24.240 2471.050 24.380 ;
        RECT 2255.910 24.180 2256.230 24.240 ;
        RECT 2470.730 24.180 2471.050 24.240 ;
      LAYER via ;
        RECT 2252.260 207.100 2252.520 207.360 ;
        RECT 2255.940 207.100 2256.200 207.360 ;
        RECT 2255.940 24.180 2256.200 24.440 ;
        RECT 2470.760 24.180 2471.020 24.440 ;
      LAYER met2 ;
        RECT 2252.300 220.000 2252.580 224.000 ;
        RECT 2252.320 207.390 2252.460 220.000 ;
        RECT 2252.260 207.070 2252.520 207.390 ;
        RECT 2255.940 207.070 2256.200 207.390 ;
        RECT 2256.000 24.470 2256.140 207.070 ;
        RECT 2255.940 24.150 2256.200 24.470 ;
        RECT 2470.760 24.150 2471.020 24.470 ;
        RECT 2470.820 2.400 2470.960 24.150 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 25.060 2270.030 25.120 ;
        RECT 2488.670 25.060 2488.990 25.120 ;
        RECT 2269.710 24.920 2488.990 25.060 ;
        RECT 2269.710 24.860 2270.030 24.920 ;
        RECT 2488.670 24.860 2488.990 24.920 ;
      LAYER via ;
        RECT 2269.740 24.860 2270.000 25.120 ;
        RECT 2488.700 24.860 2488.960 25.120 ;
      LAYER met2 ;
        RECT 2267.020 220.730 2267.300 224.000 ;
        RECT 2267.020 220.590 2269.940 220.730 ;
        RECT 2267.020 220.000 2267.300 220.590 ;
        RECT 2269.800 25.150 2269.940 220.590 ;
        RECT 2269.740 24.830 2270.000 25.150 ;
        RECT 2488.700 24.830 2488.960 25.150 ;
        RECT 2488.760 2.400 2488.900 24.830 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2311.645 24.565 2311.815 26.435 ;
      LAYER mcon ;
        RECT 2311.645 26.265 2311.815 26.435 ;
      LAYER met1 ;
        RECT 2283.510 26.420 2283.830 26.480 ;
        RECT 2311.585 26.420 2311.875 26.465 ;
        RECT 2283.510 26.280 2311.875 26.420 ;
        RECT 2283.510 26.220 2283.830 26.280 ;
        RECT 2311.585 26.235 2311.875 26.280 ;
        RECT 2311.585 24.720 2311.875 24.765 ;
        RECT 2506.150 24.720 2506.470 24.780 ;
        RECT 2311.585 24.580 2506.470 24.720 ;
        RECT 2311.585 24.535 2311.875 24.580 ;
        RECT 2506.150 24.520 2506.470 24.580 ;
      LAYER via ;
        RECT 2283.540 26.220 2283.800 26.480 ;
        RECT 2506.180 24.520 2506.440 24.780 ;
      LAYER met2 ;
        RECT 2281.740 220.730 2282.020 224.000 ;
        RECT 2281.740 220.590 2283.740 220.730 ;
        RECT 2281.740 220.000 2282.020 220.590 ;
        RECT 2283.600 26.510 2283.740 220.590 ;
        RECT 2283.540 26.190 2283.800 26.510 ;
        RECT 2506.180 24.490 2506.440 24.810 ;
        RECT 2506.240 2.400 2506.380 24.490 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2297.310 23.700 2297.630 23.760 ;
        RECT 2524.090 23.700 2524.410 23.760 ;
        RECT 2297.310 23.560 2524.410 23.700 ;
        RECT 2297.310 23.500 2297.630 23.560 ;
        RECT 2524.090 23.500 2524.410 23.560 ;
      LAYER via ;
        RECT 2297.340 23.500 2297.600 23.760 ;
        RECT 2524.120 23.500 2524.380 23.760 ;
      LAYER met2 ;
        RECT 2296.460 220.730 2296.740 224.000 ;
        RECT 2296.460 220.590 2297.540 220.730 ;
        RECT 2296.460 220.000 2296.740 220.590 ;
        RECT 2297.400 23.790 2297.540 220.590 ;
        RECT 2297.340 23.470 2297.600 23.790 ;
        RECT 2524.120 23.470 2524.380 23.790 ;
        RECT 2524.180 2.400 2524.320 23.470 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2311.110 24.040 2311.430 24.100 ;
        RECT 2542.030 24.040 2542.350 24.100 ;
        RECT 2311.110 23.900 2542.350 24.040 ;
        RECT 2311.110 23.840 2311.430 23.900 ;
        RECT 2542.030 23.840 2542.350 23.900 ;
      LAYER via ;
        RECT 2311.140 23.840 2311.400 24.100 ;
        RECT 2542.060 23.840 2542.320 24.100 ;
      LAYER met2 ;
        RECT 2311.180 220.000 2311.460 224.000 ;
        RECT 2311.200 24.130 2311.340 220.000 ;
        RECT 2311.140 23.810 2311.400 24.130 ;
        RECT 2542.060 23.810 2542.320 24.130 ;
        RECT 2542.120 2.400 2542.260 23.810 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2325.830 207.300 2326.150 207.360 ;
        RECT 2331.350 207.300 2331.670 207.360 ;
        RECT 2325.830 207.160 2331.670 207.300 ;
        RECT 2325.830 207.100 2326.150 207.160 ;
        RECT 2331.350 207.100 2331.670 207.160 ;
        RECT 2331.350 27.440 2331.670 27.500 ;
        RECT 2559.970 27.440 2560.290 27.500 ;
        RECT 2331.350 27.300 2560.290 27.440 ;
        RECT 2331.350 27.240 2331.670 27.300 ;
        RECT 2559.970 27.240 2560.290 27.300 ;
      LAYER via ;
        RECT 2325.860 207.100 2326.120 207.360 ;
        RECT 2331.380 207.100 2331.640 207.360 ;
        RECT 2331.380 27.240 2331.640 27.500 ;
        RECT 2560.000 27.240 2560.260 27.500 ;
      LAYER met2 ;
        RECT 2325.900 220.000 2326.180 224.000 ;
        RECT 2325.920 207.390 2326.060 220.000 ;
        RECT 2325.860 207.070 2326.120 207.390 ;
        RECT 2331.380 207.070 2331.640 207.390 ;
        RECT 2331.440 27.530 2331.580 207.070 ;
        RECT 2331.380 27.210 2331.640 27.530 ;
        RECT 2560.000 27.210 2560.260 27.530 ;
        RECT 2560.060 2.400 2560.200 27.210 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2340.550 207.300 2340.870 207.360 ;
        RECT 2345.610 207.300 2345.930 207.360 ;
        RECT 2340.550 207.160 2345.930 207.300 ;
        RECT 2340.550 207.100 2340.870 207.160 ;
        RECT 2345.610 207.100 2345.930 207.160 ;
        RECT 2345.610 30.840 2345.930 30.900 ;
        RECT 2577.910 30.840 2578.230 30.900 ;
        RECT 2345.610 30.700 2578.230 30.840 ;
        RECT 2345.610 30.640 2345.930 30.700 ;
        RECT 2577.910 30.640 2578.230 30.700 ;
      LAYER via ;
        RECT 2340.580 207.100 2340.840 207.360 ;
        RECT 2345.640 207.100 2345.900 207.360 ;
        RECT 2345.640 30.640 2345.900 30.900 ;
        RECT 2577.940 30.640 2578.200 30.900 ;
      LAYER met2 ;
        RECT 2340.620 220.000 2340.900 224.000 ;
        RECT 2340.640 207.390 2340.780 220.000 ;
        RECT 2340.580 207.070 2340.840 207.390 ;
        RECT 2345.640 207.070 2345.900 207.390 ;
        RECT 2345.700 30.930 2345.840 207.070 ;
        RECT 2345.640 30.610 2345.900 30.930 ;
        RECT 2577.940 30.610 2578.200 30.930 ;
        RECT 2578.000 2.400 2578.140 30.610 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 813.810 210.360 814.130 210.420 ;
        RECT 885.570 210.360 885.890 210.420 ;
        RECT 813.810 210.220 885.890 210.360 ;
        RECT 813.810 210.160 814.130 210.220 ;
        RECT 885.570 210.160 885.890 210.220 ;
        RECT 811.510 17.580 811.830 17.640 ;
        RECT 813.810 17.580 814.130 17.640 ;
        RECT 811.510 17.440 814.130 17.580 ;
        RECT 811.510 17.380 811.830 17.440 ;
        RECT 813.810 17.380 814.130 17.440 ;
      LAYER via ;
        RECT 813.840 210.160 814.100 210.420 ;
        RECT 885.600 210.160 885.860 210.420 ;
        RECT 811.540 17.380 811.800 17.640 ;
        RECT 813.840 17.380 814.100 17.640 ;
      LAYER met2 ;
        RECT 885.640 220.000 885.920 224.000 ;
        RECT 885.660 210.450 885.800 220.000 ;
        RECT 813.840 210.130 814.100 210.450 ;
        RECT 885.600 210.130 885.860 210.450 ;
        RECT 813.900 17.670 814.040 210.130 ;
        RECT 811.540 17.350 811.800 17.670 ;
        RECT 813.840 17.350 814.100 17.670 ;
        RECT 811.600 2.400 811.740 17.350 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2355.270 207.300 2355.590 207.360 ;
        RECT 2359.410 207.300 2359.730 207.360 ;
        RECT 2355.270 207.160 2359.730 207.300 ;
        RECT 2355.270 207.100 2355.590 207.160 ;
        RECT 2359.410 207.100 2359.730 207.160 ;
        RECT 2359.410 32.880 2359.730 32.940 ;
        RECT 2595.390 32.880 2595.710 32.940 ;
        RECT 2359.410 32.740 2595.710 32.880 ;
        RECT 2359.410 32.680 2359.730 32.740 ;
        RECT 2595.390 32.680 2595.710 32.740 ;
      LAYER via ;
        RECT 2355.300 207.100 2355.560 207.360 ;
        RECT 2359.440 207.100 2359.700 207.360 ;
        RECT 2359.440 32.680 2359.700 32.940 ;
        RECT 2595.420 32.680 2595.680 32.940 ;
      LAYER met2 ;
        RECT 2355.340 220.000 2355.620 224.000 ;
        RECT 2355.360 207.390 2355.500 220.000 ;
        RECT 2355.300 207.070 2355.560 207.390 ;
        RECT 2359.440 207.070 2359.700 207.390 ;
        RECT 2359.500 32.970 2359.640 207.070 ;
        RECT 2359.440 32.650 2359.700 32.970 ;
        RECT 2595.420 32.650 2595.680 32.970 ;
        RECT 2595.480 2.400 2595.620 32.650 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2373.210 32.540 2373.530 32.600 ;
        RECT 2613.330 32.540 2613.650 32.600 ;
        RECT 2373.210 32.400 2613.650 32.540 ;
        RECT 2373.210 32.340 2373.530 32.400 ;
        RECT 2613.330 32.340 2613.650 32.400 ;
      LAYER via ;
        RECT 2373.240 32.340 2373.500 32.600 ;
        RECT 2613.360 32.340 2613.620 32.600 ;
      LAYER met2 ;
        RECT 2370.060 220.730 2370.340 224.000 ;
        RECT 2370.060 220.590 2373.440 220.730 ;
        RECT 2370.060 220.000 2370.340 220.590 ;
        RECT 2373.300 32.630 2373.440 220.590 ;
        RECT 2373.240 32.310 2373.500 32.630 ;
        RECT 2613.360 32.310 2613.620 32.630 ;
        RECT 2613.420 2.400 2613.560 32.310 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2387.010 32.200 2387.330 32.260 ;
        RECT 2631.270 32.200 2631.590 32.260 ;
        RECT 2387.010 32.060 2631.590 32.200 ;
        RECT 2387.010 32.000 2387.330 32.060 ;
        RECT 2631.270 32.000 2631.590 32.060 ;
      LAYER via ;
        RECT 2387.040 32.000 2387.300 32.260 ;
        RECT 2631.300 32.000 2631.560 32.260 ;
      LAYER met2 ;
        RECT 2384.320 220.730 2384.600 224.000 ;
        RECT 2384.320 220.590 2387.240 220.730 ;
        RECT 2384.320 220.000 2384.600 220.590 ;
        RECT 2387.100 32.290 2387.240 220.590 ;
        RECT 2387.040 31.970 2387.300 32.290 ;
        RECT 2631.300 31.970 2631.560 32.290 ;
        RECT 2631.360 2.400 2631.500 31.970 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2400.810 27.100 2401.130 27.160 ;
        RECT 2649.210 27.100 2649.530 27.160 ;
        RECT 2400.810 26.960 2649.530 27.100 ;
        RECT 2400.810 26.900 2401.130 26.960 ;
        RECT 2649.210 26.900 2649.530 26.960 ;
      LAYER via ;
        RECT 2400.840 26.900 2401.100 27.160 ;
        RECT 2649.240 26.900 2649.500 27.160 ;
      LAYER met2 ;
        RECT 2399.040 220.730 2399.320 224.000 ;
        RECT 2399.040 220.590 2401.040 220.730 ;
        RECT 2399.040 220.000 2399.320 220.590 ;
        RECT 2400.900 27.190 2401.040 220.590 ;
        RECT 2400.840 26.870 2401.100 27.190 ;
        RECT 2649.240 26.870 2649.500 27.190 ;
        RECT 2649.300 2.400 2649.440 26.870 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2414.150 26.420 2414.470 26.480 ;
        RECT 2667.150 26.420 2667.470 26.480 ;
        RECT 2414.150 26.280 2667.470 26.420 ;
        RECT 2414.150 26.220 2414.470 26.280 ;
        RECT 2667.150 26.220 2667.470 26.280 ;
      LAYER via ;
        RECT 2414.180 26.220 2414.440 26.480 ;
        RECT 2667.180 26.220 2667.440 26.480 ;
      LAYER met2 ;
        RECT 2413.760 220.730 2414.040 224.000 ;
        RECT 2413.760 220.590 2414.380 220.730 ;
        RECT 2413.760 220.000 2414.040 220.590 ;
        RECT 2414.240 26.510 2414.380 220.590 ;
        RECT 2414.180 26.190 2414.440 26.510 ;
        RECT 2667.180 26.190 2667.440 26.510 ;
        RECT 2667.240 2.400 2667.380 26.190 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2428.410 25.740 2428.730 25.800 ;
        RECT 2684.630 25.740 2684.950 25.800 ;
        RECT 2428.410 25.600 2684.950 25.740 ;
        RECT 2428.410 25.540 2428.730 25.600 ;
        RECT 2684.630 25.540 2684.950 25.600 ;
      LAYER via ;
        RECT 2428.440 25.540 2428.700 25.800 ;
        RECT 2684.660 25.540 2684.920 25.800 ;
      LAYER met2 ;
        RECT 2428.480 220.000 2428.760 224.000 ;
        RECT 2428.500 25.830 2428.640 220.000 ;
        RECT 2428.440 25.510 2428.700 25.830 ;
        RECT 2684.660 25.510 2684.920 25.830 ;
        RECT 2684.720 2.400 2684.860 25.510 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2443.130 207.300 2443.450 207.360 ;
        RECT 2448.650 207.300 2448.970 207.360 ;
        RECT 2443.130 207.160 2448.970 207.300 ;
        RECT 2443.130 207.100 2443.450 207.160 ;
        RECT 2448.650 207.100 2448.970 207.160 ;
        RECT 2448.650 26.760 2448.970 26.820 ;
        RECT 2702.570 26.760 2702.890 26.820 ;
        RECT 2448.650 26.620 2702.890 26.760 ;
        RECT 2448.650 26.560 2448.970 26.620 ;
        RECT 2702.570 26.560 2702.890 26.620 ;
      LAYER via ;
        RECT 2443.160 207.100 2443.420 207.360 ;
        RECT 2448.680 207.100 2448.940 207.360 ;
        RECT 2448.680 26.560 2448.940 26.820 ;
        RECT 2702.600 26.560 2702.860 26.820 ;
      LAYER met2 ;
        RECT 2443.200 220.000 2443.480 224.000 ;
        RECT 2443.220 207.390 2443.360 220.000 ;
        RECT 2443.160 207.070 2443.420 207.390 ;
        RECT 2448.680 207.070 2448.940 207.390 ;
        RECT 2448.740 26.850 2448.880 207.070 ;
        RECT 2448.680 26.530 2448.940 26.850 ;
        RECT 2702.600 26.530 2702.860 26.850 ;
        RECT 2702.660 2.400 2702.800 26.530 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2457.850 207.300 2458.170 207.360 ;
        RECT 2462.450 207.300 2462.770 207.360 ;
        RECT 2457.850 207.160 2462.770 207.300 ;
        RECT 2457.850 207.100 2458.170 207.160 ;
        RECT 2462.450 207.100 2462.770 207.160 ;
        RECT 2462.450 25.400 2462.770 25.460 ;
        RECT 2720.510 25.400 2720.830 25.460 ;
        RECT 2462.450 25.260 2720.830 25.400 ;
        RECT 2462.450 25.200 2462.770 25.260 ;
        RECT 2720.510 25.200 2720.830 25.260 ;
      LAYER via ;
        RECT 2457.880 207.100 2458.140 207.360 ;
        RECT 2462.480 207.100 2462.740 207.360 ;
        RECT 2462.480 25.200 2462.740 25.460 ;
        RECT 2720.540 25.200 2720.800 25.460 ;
      LAYER met2 ;
        RECT 2457.920 220.000 2458.200 224.000 ;
        RECT 2457.940 207.390 2458.080 220.000 ;
        RECT 2457.880 207.070 2458.140 207.390 ;
        RECT 2462.480 207.070 2462.740 207.390 ;
        RECT 2462.540 25.490 2462.680 207.070 ;
        RECT 2462.480 25.170 2462.740 25.490 ;
        RECT 2720.540 25.170 2720.800 25.490 ;
        RECT 2720.600 2.400 2720.740 25.170 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2472.570 207.300 2472.890 207.360 ;
        RECT 2476.710 207.300 2477.030 207.360 ;
        RECT 2472.570 207.160 2477.030 207.300 ;
        RECT 2472.570 207.100 2472.890 207.160 ;
        RECT 2476.710 207.100 2477.030 207.160 ;
        RECT 2476.710 26.080 2477.030 26.140 ;
        RECT 2738.450 26.080 2738.770 26.140 ;
        RECT 2476.710 25.940 2738.770 26.080 ;
        RECT 2476.710 25.880 2477.030 25.940 ;
        RECT 2738.450 25.880 2738.770 25.940 ;
      LAYER via ;
        RECT 2472.600 207.100 2472.860 207.360 ;
        RECT 2476.740 207.100 2477.000 207.360 ;
        RECT 2476.740 25.880 2477.000 26.140 ;
        RECT 2738.480 25.880 2738.740 26.140 ;
      LAYER met2 ;
        RECT 2472.640 220.000 2472.920 224.000 ;
        RECT 2472.660 207.390 2472.800 220.000 ;
        RECT 2472.600 207.070 2472.860 207.390 ;
        RECT 2476.740 207.070 2477.000 207.390 ;
        RECT 2476.800 26.170 2476.940 207.070 ;
        RECT 2476.740 25.850 2477.000 26.170 ;
        RECT 2738.480 25.850 2738.740 26.170 ;
        RECT 2738.540 2.400 2738.680 25.850 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2490.510 25.060 2490.830 25.120 ;
        RECT 2755.930 25.060 2756.250 25.120 ;
        RECT 2490.510 24.920 2756.250 25.060 ;
        RECT 2490.510 24.860 2490.830 24.920 ;
        RECT 2755.930 24.860 2756.250 24.920 ;
      LAYER via ;
        RECT 2490.540 24.860 2490.800 25.120 ;
        RECT 2755.960 24.860 2756.220 25.120 ;
      LAYER met2 ;
        RECT 2487.360 220.730 2487.640 224.000 ;
        RECT 2487.360 220.590 2490.740 220.730 ;
        RECT 2487.360 220.000 2487.640 220.590 ;
        RECT 2490.600 25.150 2490.740 220.590 ;
        RECT 2490.540 24.830 2490.800 25.150 ;
        RECT 2755.960 24.830 2756.220 25.150 ;
        RECT 2756.020 2.400 2756.160 24.830 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 834.510 209.000 834.830 209.060 ;
        RECT 900.290 209.000 900.610 209.060 ;
        RECT 834.510 208.860 900.610 209.000 ;
        RECT 834.510 208.800 834.830 208.860 ;
        RECT 900.290 208.800 900.610 208.860 ;
        RECT 829.450 17.580 829.770 17.640 ;
        RECT 834.510 17.580 834.830 17.640 ;
        RECT 829.450 17.440 834.830 17.580 ;
        RECT 829.450 17.380 829.770 17.440 ;
        RECT 834.510 17.380 834.830 17.440 ;
      LAYER via ;
        RECT 834.540 208.800 834.800 209.060 ;
        RECT 900.320 208.800 900.580 209.060 ;
        RECT 829.480 17.380 829.740 17.640 ;
        RECT 834.540 17.380 834.800 17.640 ;
      LAYER met2 ;
        RECT 900.360 220.000 900.640 224.000 ;
        RECT 900.380 209.090 900.520 220.000 ;
        RECT 834.540 208.770 834.800 209.090 ;
        RECT 900.320 208.770 900.580 209.090 ;
        RECT 834.600 17.670 834.740 208.770 ;
        RECT 829.480 17.350 829.740 17.670 ;
        RECT 834.540 17.350 834.800 17.670 ;
        RECT 829.540 2.400 829.680 17.350 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2504.310 24.380 2504.630 24.440 ;
        RECT 2773.870 24.380 2774.190 24.440 ;
        RECT 2504.310 24.240 2774.190 24.380 ;
        RECT 2504.310 24.180 2504.630 24.240 ;
        RECT 2773.870 24.180 2774.190 24.240 ;
      LAYER via ;
        RECT 2504.340 24.180 2504.600 24.440 ;
        RECT 2773.900 24.180 2774.160 24.440 ;
      LAYER met2 ;
        RECT 2502.080 220.730 2502.360 224.000 ;
        RECT 2502.080 220.590 2504.540 220.730 ;
        RECT 2502.080 220.000 2502.360 220.590 ;
        RECT 2504.400 24.470 2504.540 220.590 ;
        RECT 2504.340 24.150 2504.600 24.470 ;
        RECT 2773.900 24.150 2774.160 24.470 ;
        RECT 2773.960 2.400 2774.100 24.150 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2518.110 24.720 2518.430 24.780 ;
        RECT 2791.810 24.720 2792.130 24.780 ;
        RECT 2518.110 24.580 2792.130 24.720 ;
        RECT 2518.110 24.520 2518.430 24.580 ;
        RECT 2791.810 24.520 2792.130 24.580 ;
      LAYER via ;
        RECT 2518.140 24.520 2518.400 24.780 ;
        RECT 2791.840 24.520 2792.100 24.780 ;
      LAYER met2 ;
        RECT 2516.800 220.730 2517.080 224.000 ;
        RECT 2516.800 220.590 2518.340 220.730 ;
        RECT 2516.800 220.000 2517.080 220.590 ;
        RECT 2518.200 24.810 2518.340 220.590 ;
        RECT 2518.140 24.490 2518.400 24.810 ;
        RECT 2791.840 24.490 2792.100 24.810 ;
        RECT 2791.900 2.400 2792.040 24.490 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2531.450 31.180 2531.770 31.240 ;
        RECT 2809.750 31.180 2810.070 31.240 ;
        RECT 2531.450 31.040 2810.070 31.180 ;
        RECT 2531.450 30.980 2531.770 31.040 ;
        RECT 2809.750 30.980 2810.070 31.040 ;
      LAYER via ;
        RECT 2531.480 30.980 2531.740 31.240 ;
        RECT 2809.780 30.980 2810.040 31.240 ;
      LAYER met2 ;
        RECT 2531.520 220.000 2531.800 224.000 ;
        RECT 2531.540 31.270 2531.680 220.000 ;
        RECT 2531.480 30.950 2531.740 31.270 ;
        RECT 2809.780 30.950 2810.040 31.270 ;
        RECT 2809.840 2.400 2809.980 30.950 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2546.170 207.300 2546.490 207.360 ;
        RECT 2552.150 207.300 2552.470 207.360 ;
        RECT 2546.170 207.160 2552.470 207.300 ;
        RECT 2546.170 207.100 2546.490 207.160 ;
        RECT 2552.150 207.100 2552.470 207.160 ;
        RECT 2552.150 24.040 2552.470 24.100 ;
        RECT 2827.690 24.040 2828.010 24.100 ;
        RECT 2552.150 23.900 2828.010 24.040 ;
        RECT 2552.150 23.840 2552.470 23.900 ;
        RECT 2827.690 23.840 2828.010 23.900 ;
      LAYER via ;
        RECT 2546.200 207.100 2546.460 207.360 ;
        RECT 2552.180 207.100 2552.440 207.360 ;
        RECT 2552.180 23.840 2552.440 24.100 ;
        RECT 2827.720 23.840 2827.980 24.100 ;
      LAYER met2 ;
        RECT 2546.240 220.000 2546.520 224.000 ;
        RECT 2546.260 207.390 2546.400 220.000 ;
        RECT 2546.200 207.070 2546.460 207.390 ;
        RECT 2552.180 207.070 2552.440 207.390 ;
        RECT 2552.240 24.130 2552.380 207.070 ;
        RECT 2552.180 23.810 2552.440 24.130 ;
        RECT 2827.720 23.810 2827.980 24.130 ;
        RECT 2827.780 2.400 2827.920 23.810 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2560.890 207.300 2561.210 207.360 ;
        RECT 2566.410 207.300 2566.730 207.360 ;
        RECT 2560.890 207.160 2566.730 207.300 ;
        RECT 2560.890 207.100 2561.210 207.160 ;
        RECT 2566.410 207.100 2566.730 207.160 ;
        RECT 2566.410 31.860 2566.730 31.920 ;
        RECT 2845.170 31.860 2845.490 31.920 ;
        RECT 2566.410 31.720 2845.490 31.860 ;
        RECT 2566.410 31.660 2566.730 31.720 ;
        RECT 2845.170 31.660 2845.490 31.720 ;
      LAYER via ;
        RECT 2560.920 207.100 2561.180 207.360 ;
        RECT 2566.440 207.100 2566.700 207.360 ;
        RECT 2566.440 31.660 2566.700 31.920 ;
        RECT 2845.200 31.660 2845.460 31.920 ;
      LAYER met2 ;
        RECT 2560.960 220.000 2561.240 224.000 ;
        RECT 2560.980 207.390 2561.120 220.000 ;
        RECT 2560.920 207.070 2561.180 207.390 ;
        RECT 2566.440 207.070 2566.700 207.390 ;
        RECT 2566.500 31.950 2566.640 207.070 ;
        RECT 2566.440 31.630 2566.700 31.950 ;
        RECT 2845.200 31.630 2845.460 31.950 ;
        RECT 2845.260 2.400 2845.400 31.630 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2575.610 207.300 2575.930 207.360 ;
        RECT 2579.750 207.300 2580.070 207.360 ;
        RECT 2575.610 207.160 2580.070 207.300 ;
        RECT 2575.610 207.100 2575.930 207.160 ;
        RECT 2579.750 207.100 2580.070 207.160 ;
        RECT 2579.750 31.520 2580.070 31.580 ;
        RECT 2863.110 31.520 2863.430 31.580 ;
        RECT 2579.750 31.380 2863.430 31.520 ;
        RECT 2579.750 31.320 2580.070 31.380 ;
        RECT 2863.110 31.320 2863.430 31.380 ;
      LAYER via ;
        RECT 2575.640 207.100 2575.900 207.360 ;
        RECT 2579.780 207.100 2580.040 207.360 ;
        RECT 2579.780 31.320 2580.040 31.580 ;
        RECT 2863.140 31.320 2863.400 31.580 ;
      LAYER met2 ;
        RECT 2575.680 220.000 2575.960 224.000 ;
        RECT 2575.700 207.390 2575.840 220.000 ;
        RECT 2575.640 207.070 2575.900 207.390 ;
        RECT 2579.780 207.070 2580.040 207.390 ;
        RECT 2579.840 31.610 2579.980 207.070 ;
        RECT 2579.780 31.290 2580.040 31.610 ;
        RECT 2863.140 31.290 2863.400 31.610 ;
        RECT 2863.200 2.400 2863.340 31.290 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2594.010 30.840 2594.330 30.900 ;
        RECT 2881.050 30.840 2881.370 30.900 ;
        RECT 2594.010 30.700 2881.370 30.840 ;
        RECT 2594.010 30.640 2594.330 30.700 ;
        RECT 2881.050 30.640 2881.370 30.700 ;
      LAYER via ;
        RECT 2594.040 30.640 2594.300 30.900 ;
        RECT 2881.080 30.640 2881.340 30.900 ;
      LAYER met2 ;
        RECT 2590.400 220.730 2590.680 224.000 ;
        RECT 2590.400 220.590 2594.240 220.730 ;
        RECT 2590.400 220.000 2590.680 220.590 ;
        RECT 2594.100 30.930 2594.240 220.590 ;
        RECT 2594.040 30.610 2594.300 30.930 ;
        RECT 2881.080 30.610 2881.340 30.930 ;
        RECT 2881.140 2.400 2881.280 30.610 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2673.205 15.045 2673.375 16.575 ;
      LAYER mcon ;
        RECT 2673.205 16.405 2673.375 16.575 ;
      LAYER met1 ;
        RECT 2605.050 207.980 2605.370 208.040 ;
        RECT 2645.990 207.980 2646.310 208.040 ;
        RECT 2605.050 207.840 2646.310 207.980 ;
        RECT 2605.050 207.780 2605.370 207.840 ;
        RECT 2645.990 207.780 2646.310 207.840 ;
        RECT 2673.145 16.560 2673.435 16.605 ;
        RECT 2898.990 16.560 2899.310 16.620 ;
        RECT 2673.145 16.420 2899.310 16.560 ;
        RECT 2673.145 16.375 2673.435 16.420 ;
        RECT 2898.990 16.360 2899.310 16.420 ;
        RECT 2645.990 15.200 2646.310 15.260 ;
        RECT 2673.145 15.200 2673.435 15.245 ;
        RECT 2645.990 15.060 2673.435 15.200 ;
        RECT 2645.990 15.000 2646.310 15.060 ;
        RECT 2673.145 15.015 2673.435 15.060 ;
      LAYER via ;
        RECT 2605.080 207.780 2605.340 208.040 ;
        RECT 2646.020 207.780 2646.280 208.040 ;
        RECT 2899.020 16.360 2899.280 16.620 ;
        RECT 2646.020 15.000 2646.280 15.260 ;
      LAYER met2 ;
        RECT 2605.120 220.000 2605.400 224.000 ;
        RECT 2605.140 208.070 2605.280 220.000 ;
        RECT 2605.080 207.750 2605.340 208.070 ;
        RECT 2646.020 207.750 2646.280 208.070 ;
        RECT 2646.080 15.290 2646.220 207.750 ;
        RECT 2899.020 16.330 2899.280 16.650 ;
        RECT 2646.020 14.970 2646.280 15.290 ;
        RECT 2899.080 2.400 2899.220 16.330 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 848.310 213.420 848.630 213.480 ;
        RECT 915.010 213.420 915.330 213.480 ;
        RECT 848.310 213.280 915.330 213.420 ;
        RECT 848.310 213.220 848.630 213.280 ;
        RECT 915.010 213.220 915.330 213.280 ;
        RECT 846.930 14.180 847.250 14.240 ;
        RECT 848.310 14.180 848.630 14.240 ;
        RECT 846.930 14.040 848.630 14.180 ;
        RECT 846.930 13.980 847.250 14.040 ;
        RECT 848.310 13.980 848.630 14.040 ;
      LAYER via ;
        RECT 848.340 213.220 848.600 213.480 ;
        RECT 915.040 213.220 915.300 213.480 ;
        RECT 846.960 13.980 847.220 14.240 ;
        RECT 848.340 13.980 848.600 14.240 ;
      LAYER met2 ;
        RECT 915.080 220.000 915.360 224.000 ;
        RECT 915.100 213.510 915.240 220.000 ;
        RECT 848.340 213.190 848.600 213.510 ;
        RECT 915.040 213.190 915.300 213.510 ;
        RECT 848.400 14.270 848.540 213.190 ;
        RECT 846.960 13.950 847.220 14.270 ;
        RECT 848.340 13.950 848.600 14.270 ;
        RECT 847.020 2.400 847.160 13.950 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 869.010 213.760 869.330 213.820 ;
        RECT 929.730 213.760 930.050 213.820 ;
        RECT 869.010 213.620 930.050 213.760 ;
        RECT 869.010 213.560 869.330 213.620 ;
        RECT 929.730 213.560 930.050 213.620 ;
        RECT 864.870 17.580 865.190 17.640 ;
        RECT 869.010 17.580 869.330 17.640 ;
        RECT 864.870 17.440 869.330 17.580 ;
        RECT 864.870 17.380 865.190 17.440 ;
        RECT 869.010 17.380 869.330 17.440 ;
      LAYER via ;
        RECT 869.040 213.560 869.300 213.820 ;
        RECT 929.760 213.560 930.020 213.820 ;
        RECT 864.900 17.380 865.160 17.640 ;
        RECT 869.040 17.380 869.300 17.640 ;
      LAYER met2 ;
        RECT 929.800 220.000 930.080 224.000 ;
        RECT 929.820 213.850 929.960 220.000 ;
        RECT 869.040 213.530 869.300 213.850 ;
        RECT 929.760 213.530 930.020 213.850 ;
        RECT 869.100 17.670 869.240 213.530 ;
        RECT 864.900 17.350 865.160 17.670 ;
        RECT 869.040 17.350 869.300 17.670 ;
        RECT 864.960 2.400 865.100 17.350 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.810 210.020 883.130 210.080 ;
        RECT 944.450 210.020 944.770 210.080 ;
        RECT 882.810 209.880 944.770 210.020 ;
        RECT 882.810 209.820 883.130 209.880 ;
        RECT 944.450 209.820 944.770 209.880 ;
      LAYER via ;
        RECT 882.840 209.820 883.100 210.080 ;
        RECT 944.480 209.820 944.740 210.080 ;
      LAYER met2 ;
        RECT 944.520 220.000 944.800 224.000 ;
        RECT 944.540 210.110 944.680 220.000 ;
        RECT 882.840 209.790 883.100 210.110 ;
        RECT 944.480 209.790 944.740 210.110 ;
        RECT 882.900 2.400 883.040 209.790 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 903.510 211.380 903.830 211.440 ;
        RECT 959.170 211.380 959.490 211.440 ;
        RECT 903.510 211.240 959.490 211.380 ;
        RECT 903.510 211.180 903.830 211.240 ;
        RECT 959.170 211.180 959.490 211.240 ;
        RECT 900.750 17.580 901.070 17.640 ;
        RECT 903.510 17.580 903.830 17.640 ;
        RECT 900.750 17.440 903.830 17.580 ;
        RECT 900.750 17.380 901.070 17.440 ;
        RECT 903.510 17.380 903.830 17.440 ;
      LAYER via ;
        RECT 903.540 211.180 903.800 211.440 ;
        RECT 959.200 211.180 959.460 211.440 ;
        RECT 900.780 17.380 901.040 17.640 ;
        RECT 903.540 17.380 903.800 17.640 ;
      LAYER met2 ;
        RECT 959.240 220.000 959.520 224.000 ;
        RECT 959.260 211.470 959.400 220.000 ;
        RECT 903.540 211.150 903.800 211.470 ;
        RECT 959.200 211.150 959.460 211.470 ;
        RECT 903.600 17.670 903.740 211.150 ;
        RECT 900.780 17.350 901.040 17.670 ;
        RECT 903.540 17.350 903.800 17.670 ;
        RECT 900.840 2.400 900.980 17.350 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 924.210 209.680 924.530 209.740 ;
        RECT 973.890 209.680 974.210 209.740 ;
        RECT 924.210 209.540 974.210 209.680 ;
        RECT 924.210 209.480 924.530 209.540 ;
        RECT 973.890 209.480 974.210 209.540 ;
        RECT 918.690 17.920 919.010 17.980 ;
        RECT 924.210 17.920 924.530 17.980 ;
        RECT 918.690 17.780 924.530 17.920 ;
        RECT 918.690 17.720 919.010 17.780 ;
        RECT 924.210 17.720 924.530 17.780 ;
      LAYER via ;
        RECT 924.240 209.480 924.500 209.740 ;
        RECT 973.920 209.480 974.180 209.740 ;
        RECT 918.720 17.720 918.980 17.980 ;
        RECT 924.240 17.720 924.500 17.980 ;
      LAYER met2 ;
        RECT 973.960 220.000 974.240 224.000 ;
        RECT 973.980 209.770 974.120 220.000 ;
        RECT 924.240 209.450 924.500 209.770 ;
        RECT 973.920 209.450 974.180 209.770 ;
        RECT 924.300 18.010 924.440 209.450 ;
        RECT 918.720 17.690 918.980 18.010 ;
        RECT 924.240 17.690 924.500 18.010 ;
        RECT 918.780 2.400 918.920 17.690 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 938.010 212.400 938.330 212.460 ;
        RECT 988.610 212.400 988.930 212.460 ;
        RECT 938.010 212.260 988.930 212.400 ;
        RECT 938.010 212.200 938.330 212.260 ;
        RECT 988.610 212.200 988.930 212.260 ;
      LAYER via ;
        RECT 938.040 212.200 938.300 212.460 ;
        RECT 988.640 212.200 988.900 212.460 ;
      LAYER met2 ;
        RECT 988.680 220.000 988.960 224.000 ;
        RECT 988.700 212.490 988.840 220.000 ;
        RECT 938.040 212.170 938.300 212.490 ;
        RECT 988.640 212.170 988.900 212.490 ;
        RECT 938.100 17.410 938.240 212.170 ;
        RECT 936.260 17.270 938.240 17.410 ;
        RECT 936.260 2.400 936.400 17.270 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 958.710 212.060 959.030 212.120 ;
        RECT 1003.330 212.060 1003.650 212.120 ;
        RECT 958.710 211.920 1003.650 212.060 ;
        RECT 958.710 211.860 959.030 211.920 ;
        RECT 1003.330 211.860 1003.650 211.920 ;
        RECT 954.110 15.200 954.430 15.260 ;
        RECT 958.710 15.200 959.030 15.260 ;
        RECT 954.110 15.060 959.030 15.200 ;
        RECT 954.110 15.000 954.430 15.060 ;
        RECT 958.710 15.000 959.030 15.060 ;
      LAYER via ;
        RECT 958.740 211.860 959.000 212.120 ;
        RECT 1003.360 211.860 1003.620 212.120 ;
        RECT 954.140 15.000 954.400 15.260 ;
        RECT 958.740 15.000 959.000 15.260 ;
      LAYER met2 ;
        RECT 1003.400 220.000 1003.680 224.000 ;
        RECT 1003.420 212.150 1003.560 220.000 ;
        RECT 958.740 211.830 959.000 212.150 ;
        RECT 1003.360 211.830 1003.620 212.150 ;
        RECT 958.800 15.290 958.940 211.830 ;
        RECT 954.140 14.970 954.400 15.290 ;
        RECT 958.740 14.970 959.000 15.290 ;
        RECT 954.200 2.400 954.340 14.970 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.050 210.360 972.370 210.420 ;
        RECT 1018.050 210.360 1018.370 210.420 ;
        RECT 972.050 210.220 1018.370 210.360 ;
        RECT 972.050 210.160 972.370 210.220 ;
        RECT 1018.050 210.160 1018.370 210.220 ;
      LAYER via ;
        RECT 972.080 210.160 972.340 210.420 ;
        RECT 1018.080 210.160 1018.340 210.420 ;
      LAYER met2 ;
        RECT 1018.120 220.000 1018.400 224.000 ;
        RECT 1018.140 210.450 1018.280 220.000 ;
        RECT 972.080 210.130 972.340 210.450 ;
        RECT 1018.080 210.130 1018.340 210.450 ;
        RECT 972.140 2.400 972.280 210.130 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 655.110 209.680 655.430 209.740 ;
        RECT 753.550 209.680 753.870 209.740 ;
        RECT 655.110 209.540 753.870 209.680 ;
        RECT 655.110 209.480 655.430 209.540 ;
        RECT 753.550 209.480 753.870 209.540 ;
        RECT 650.970 17.580 651.290 17.640 ;
        RECT 655.110 17.580 655.430 17.640 ;
        RECT 650.970 17.440 655.430 17.580 ;
        RECT 650.970 17.380 651.290 17.440 ;
        RECT 655.110 17.380 655.430 17.440 ;
      LAYER via ;
        RECT 655.140 209.480 655.400 209.740 ;
        RECT 753.580 209.480 753.840 209.740 ;
        RECT 651.000 17.380 651.260 17.640 ;
        RECT 655.140 17.380 655.400 17.640 ;
      LAYER met2 ;
        RECT 753.620 220.000 753.900 224.000 ;
        RECT 753.640 209.770 753.780 220.000 ;
        RECT 655.140 209.450 655.400 209.770 ;
        RECT 753.580 209.450 753.840 209.770 ;
        RECT 655.200 17.670 655.340 209.450 ;
        RECT 651.000 17.350 651.260 17.670 ;
        RECT 655.140 17.350 655.400 17.670 ;
        RECT 651.060 2.400 651.200 17.350 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 993.210 212.400 993.530 212.460 ;
        RECT 1032.770 212.400 1033.090 212.460 ;
        RECT 993.210 212.260 1033.090 212.400 ;
        RECT 993.210 212.200 993.530 212.260 ;
        RECT 1032.770 212.200 1033.090 212.260 ;
        RECT 989.990 17.580 990.310 17.640 ;
        RECT 993.210 17.580 993.530 17.640 ;
        RECT 989.990 17.440 993.530 17.580 ;
        RECT 989.990 17.380 990.310 17.440 ;
        RECT 993.210 17.380 993.530 17.440 ;
      LAYER via ;
        RECT 993.240 212.200 993.500 212.460 ;
        RECT 1032.800 212.200 1033.060 212.460 ;
        RECT 990.020 17.380 990.280 17.640 ;
        RECT 993.240 17.380 993.500 17.640 ;
      LAYER met2 ;
        RECT 1032.840 220.000 1033.120 224.000 ;
        RECT 1032.860 212.490 1033.000 220.000 ;
        RECT 993.240 212.170 993.500 212.490 ;
        RECT 1032.800 212.170 1033.060 212.490 ;
        RECT 993.300 17.670 993.440 212.170 ;
        RECT 990.020 17.350 990.280 17.670 ;
        RECT 993.240 17.350 993.500 17.670 ;
        RECT 990.080 2.400 990.220 17.350 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1013.450 207.980 1013.770 208.040 ;
        RECT 1047.490 207.980 1047.810 208.040 ;
        RECT 1013.450 207.840 1047.810 207.980 ;
        RECT 1013.450 207.780 1013.770 207.840 ;
        RECT 1047.490 207.780 1047.810 207.840 ;
        RECT 1007.470 17.920 1007.790 17.980 ;
        RECT 1013.450 17.920 1013.770 17.980 ;
        RECT 1007.470 17.780 1013.770 17.920 ;
        RECT 1007.470 17.720 1007.790 17.780 ;
        RECT 1013.450 17.720 1013.770 17.780 ;
      LAYER via ;
        RECT 1013.480 207.780 1013.740 208.040 ;
        RECT 1047.520 207.780 1047.780 208.040 ;
        RECT 1007.500 17.720 1007.760 17.980 ;
        RECT 1013.480 17.720 1013.740 17.980 ;
      LAYER met2 ;
        RECT 1047.560 220.000 1047.840 224.000 ;
        RECT 1047.580 208.070 1047.720 220.000 ;
        RECT 1013.480 207.750 1013.740 208.070 ;
        RECT 1047.520 207.750 1047.780 208.070 ;
        RECT 1013.540 18.010 1013.680 207.750 ;
        RECT 1007.500 17.690 1007.760 18.010 ;
        RECT 1013.480 17.690 1013.740 18.010 ;
        RECT 1007.560 2.400 1007.700 17.690 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1027.710 207.300 1028.030 207.360 ;
        RECT 1062.210 207.300 1062.530 207.360 ;
        RECT 1027.710 207.160 1062.530 207.300 ;
        RECT 1027.710 207.100 1028.030 207.160 ;
        RECT 1062.210 207.100 1062.530 207.160 ;
        RECT 1025.410 17.580 1025.730 17.640 ;
        RECT 1027.710 17.580 1028.030 17.640 ;
        RECT 1025.410 17.440 1028.030 17.580 ;
        RECT 1025.410 17.380 1025.730 17.440 ;
        RECT 1027.710 17.380 1028.030 17.440 ;
      LAYER via ;
        RECT 1027.740 207.100 1028.000 207.360 ;
        RECT 1062.240 207.100 1062.500 207.360 ;
        RECT 1025.440 17.380 1025.700 17.640 ;
        RECT 1027.740 17.380 1028.000 17.640 ;
      LAYER met2 ;
        RECT 1062.280 220.000 1062.560 224.000 ;
        RECT 1062.300 207.390 1062.440 220.000 ;
        RECT 1027.740 207.070 1028.000 207.390 ;
        RECT 1062.240 207.070 1062.500 207.390 ;
        RECT 1027.800 17.670 1027.940 207.070 ;
        RECT 1025.440 17.350 1025.700 17.670 ;
        RECT 1027.740 17.350 1028.000 17.670 ;
        RECT 1025.500 2.400 1025.640 17.350 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1048.410 211.380 1048.730 211.440 ;
        RECT 1076.930 211.380 1077.250 211.440 ;
        RECT 1048.410 211.240 1077.250 211.380 ;
        RECT 1048.410 211.180 1048.730 211.240 ;
        RECT 1076.930 211.180 1077.250 211.240 ;
        RECT 1043.350 17.580 1043.670 17.640 ;
        RECT 1048.410 17.580 1048.730 17.640 ;
        RECT 1043.350 17.440 1048.730 17.580 ;
        RECT 1043.350 17.380 1043.670 17.440 ;
        RECT 1048.410 17.380 1048.730 17.440 ;
      LAYER via ;
        RECT 1048.440 211.180 1048.700 211.440 ;
        RECT 1076.960 211.180 1077.220 211.440 ;
        RECT 1043.380 17.380 1043.640 17.640 ;
        RECT 1048.440 17.380 1048.700 17.640 ;
      LAYER met2 ;
        RECT 1077.000 220.000 1077.280 224.000 ;
        RECT 1077.020 211.470 1077.160 220.000 ;
        RECT 1048.440 211.150 1048.700 211.470 ;
        RECT 1076.960 211.150 1077.220 211.470 ;
        RECT 1048.500 17.670 1048.640 211.150 ;
        RECT 1043.380 17.350 1043.640 17.670 ;
        RECT 1048.440 17.350 1048.700 17.670 ;
        RECT 1043.440 2.400 1043.580 17.350 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1062.670 208.320 1062.990 208.380 ;
        RECT 1091.650 208.320 1091.970 208.380 ;
        RECT 1062.670 208.180 1091.970 208.320 ;
        RECT 1062.670 208.120 1062.990 208.180 ;
        RECT 1091.650 208.120 1091.970 208.180 ;
      LAYER via ;
        RECT 1062.700 208.120 1062.960 208.380 ;
        RECT 1091.680 208.120 1091.940 208.380 ;
      LAYER met2 ;
        RECT 1091.720 220.000 1092.000 224.000 ;
        RECT 1091.740 208.410 1091.880 220.000 ;
        RECT 1062.700 208.090 1062.960 208.410 ;
        RECT 1091.680 208.090 1091.940 208.410 ;
        RECT 1062.760 206.450 1062.900 208.090 ;
        RECT 1062.300 206.310 1062.900 206.450 ;
        RECT 1062.300 17.410 1062.440 206.310 ;
        RECT 1061.380 17.270 1062.440 17.410 ;
        RECT 1061.380 2.400 1061.520 17.270 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1082.910 207.300 1083.230 207.360 ;
        RECT 1106.370 207.300 1106.690 207.360 ;
        RECT 1082.910 207.160 1106.690 207.300 ;
        RECT 1082.910 207.100 1083.230 207.160 ;
        RECT 1106.370 207.100 1106.690 207.160 ;
        RECT 1079.230 17.580 1079.550 17.640 ;
        RECT 1082.910 17.580 1083.230 17.640 ;
        RECT 1079.230 17.440 1083.230 17.580 ;
        RECT 1079.230 17.380 1079.550 17.440 ;
        RECT 1082.910 17.380 1083.230 17.440 ;
      LAYER via ;
        RECT 1082.940 207.100 1083.200 207.360 ;
        RECT 1106.400 207.100 1106.660 207.360 ;
        RECT 1079.260 17.380 1079.520 17.640 ;
        RECT 1082.940 17.380 1083.200 17.640 ;
      LAYER met2 ;
        RECT 1106.440 220.000 1106.720 224.000 ;
        RECT 1106.460 207.390 1106.600 220.000 ;
        RECT 1082.940 207.070 1083.200 207.390 ;
        RECT 1106.400 207.070 1106.660 207.390 ;
        RECT 1083.000 17.670 1083.140 207.070 ;
        RECT 1079.260 17.350 1079.520 17.670 ;
        RECT 1082.940 17.350 1083.200 17.670 ;
        RECT 1079.320 2.400 1079.460 17.350 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.250 210.360 1096.570 210.420 ;
        RECT 1121.090 210.360 1121.410 210.420 ;
        RECT 1096.250 210.220 1121.410 210.360 ;
        RECT 1096.250 210.160 1096.570 210.220 ;
        RECT 1121.090 210.160 1121.410 210.220 ;
      LAYER via ;
        RECT 1096.280 210.160 1096.540 210.420 ;
        RECT 1121.120 210.160 1121.380 210.420 ;
      LAYER met2 ;
        RECT 1121.160 220.000 1121.440 224.000 ;
        RECT 1121.180 210.450 1121.320 220.000 ;
        RECT 1096.280 210.130 1096.540 210.450 ;
        RECT 1121.120 210.130 1121.380 210.450 ;
        RECT 1096.340 7.890 1096.480 210.130 ;
        RECT 1096.340 7.750 1096.940 7.890 ;
        RECT 1096.800 2.400 1096.940 7.750 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1117.410 207.300 1117.730 207.360 ;
        RECT 1135.350 207.300 1135.670 207.360 ;
        RECT 1117.410 207.160 1135.670 207.300 ;
        RECT 1117.410 207.100 1117.730 207.160 ;
        RECT 1135.350 207.100 1135.670 207.160 ;
        RECT 1114.650 17.580 1114.970 17.640 ;
        RECT 1117.410 17.580 1117.730 17.640 ;
        RECT 1114.650 17.440 1117.730 17.580 ;
        RECT 1114.650 17.380 1114.970 17.440 ;
        RECT 1117.410 17.380 1117.730 17.440 ;
      LAYER via ;
        RECT 1117.440 207.100 1117.700 207.360 ;
        RECT 1135.380 207.100 1135.640 207.360 ;
        RECT 1114.680 17.380 1114.940 17.640 ;
        RECT 1117.440 17.380 1117.700 17.640 ;
      LAYER met2 ;
        RECT 1135.420 220.000 1135.700 224.000 ;
        RECT 1135.440 207.390 1135.580 220.000 ;
        RECT 1117.440 207.070 1117.700 207.390 ;
        RECT 1135.380 207.070 1135.640 207.390 ;
        RECT 1117.500 17.670 1117.640 207.070 ;
        RECT 1114.680 17.350 1114.940 17.670 ;
        RECT 1117.440 17.350 1117.700 17.670 ;
        RECT 1114.740 2.400 1114.880 17.350 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1138.110 207.300 1138.430 207.360 ;
        RECT 1150.070 207.300 1150.390 207.360 ;
        RECT 1138.110 207.160 1150.390 207.300 ;
        RECT 1138.110 207.100 1138.430 207.160 ;
        RECT 1150.070 207.100 1150.390 207.160 ;
        RECT 1132.590 16.560 1132.910 16.620 ;
        RECT 1138.110 16.560 1138.430 16.620 ;
        RECT 1132.590 16.420 1138.430 16.560 ;
        RECT 1132.590 16.360 1132.910 16.420 ;
        RECT 1138.110 16.360 1138.430 16.420 ;
      LAYER via ;
        RECT 1138.140 207.100 1138.400 207.360 ;
        RECT 1150.100 207.100 1150.360 207.360 ;
        RECT 1132.620 16.360 1132.880 16.620 ;
        RECT 1138.140 16.360 1138.400 16.620 ;
      LAYER met2 ;
        RECT 1150.140 220.000 1150.420 224.000 ;
        RECT 1150.160 207.390 1150.300 220.000 ;
        RECT 1138.140 207.070 1138.400 207.390 ;
        RECT 1150.100 207.070 1150.360 207.390 ;
        RECT 1138.200 16.650 1138.340 207.070 ;
        RECT 1132.620 16.330 1132.880 16.650 ;
        RECT 1138.140 16.330 1138.400 16.650 ;
        RECT 1132.680 2.400 1132.820 16.330 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1151.910 207.640 1152.230 207.700 ;
        RECT 1164.790 207.640 1165.110 207.700 ;
        RECT 1151.910 207.500 1165.110 207.640 ;
        RECT 1151.910 207.440 1152.230 207.500 ;
        RECT 1164.790 207.440 1165.110 207.500 ;
      LAYER via ;
        RECT 1151.940 207.440 1152.200 207.700 ;
        RECT 1164.820 207.440 1165.080 207.700 ;
      LAYER met2 ;
        RECT 1164.860 220.000 1165.140 224.000 ;
        RECT 1164.880 207.730 1165.020 220.000 ;
        RECT 1151.940 207.410 1152.200 207.730 ;
        RECT 1164.820 207.410 1165.080 207.730 ;
        RECT 1152.000 17.410 1152.140 207.410 ;
        RECT 1150.620 17.270 1152.140 17.410 ;
        RECT 1150.620 2.400 1150.760 17.270 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 675.440 213.960 680.640 214.100 ;
        RECT 668.910 213.760 669.230 213.820 ;
        RECT 675.440 213.760 675.580 213.960 ;
        RECT 668.910 213.620 675.580 213.760 ;
        RECT 680.500 213.760 680.640 213.960 ;
        RECT 768.270 213.760 768.590 213.820 ;
        RECT 680.500 213.620 768.590 213.760 ;
        RECT 668.910 213.560 669.230 213.620 ;
        RECT 768.270 213.560 768.590 213.620 ;
      LAYER via ;
        RECT 668.940 213.560 669.200 213.820 ;
        RECT 768.300 213.560 768.560 213.820 ;
      LAYER met2 ;
        RECT 768.340 220.000 768.620 224.000 ;
        RECT 768.360 213.850 768.500 220.000 ;
        RECT 668.940 213.530 669.200 213.850 ;
        RECT 768.300 213.530 768.560 213.850 ;
        RECT 669.000 2.400 669.140 213.530 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1172.610 207.300 1172.930 207.360 ;
        RECT 1179.510 207.300 1179.830 207.360 ;
        RECT 1172.610 207.160 1179.830 207.300 ;
        RECT 1172.610 207.100 1172.930 207.160 ;
        RECT 1179.510 207.100 1179.830 207.160 ;
        RECT 1168.470 17.580 1168.790 17.640 ;
        RECT 1172.610 17.580 1172.930 17.640 ;
        RECT 1168.470 17.440 1172.930 17.580 ;
        RECT 1168.470 17.380 1168.790 17.440 ;
        RECT 1172.610 17.380 1172.930 17.440 ;
      LAYER via ;
        RECT 1172.640 207.100 1172.900 207.360 ;
        RECT 1179.540 207.100 1179.800 207.360 ;
        RECT 1168.500 17.380 1168.760 17.640 ;
        RECT 1172.640 17.380 1172.900 17.640 ;
      LAYER met2 ;
        RECT 1179.580 220.000 1179.860 224.000 ;
        RECT 1179.600 207.390 1179.740 220.000 ;
        RECT 1172.640 207.070 1172.900 207.390 ;
        RECT 1179.540 207.070 1179.800 207.390 ;
        RECT 1172.700 17.670 1172.840 207.070 ;
        RECT 1168.500 17.350 1168.760 17.670 ;
        RECT 1172.640 17.350 1172.900 17.670 ;
        RECT 1168.560 2.400 1168.700 17.350 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 213.760 1186.730 213.820 ;
        RECT 1194.230 213.760 1194.550 213.820 ;
        RECT 1186.410 213.620 1194.550 213.760 ;
        RECT 1186.410 213.560 1186.730 213.620 ;
        RECT 1194.230 213.560 1194.550 213.620 ;
      LAYER via ;
        RECT 1186.440 213.560 1186.700 213.820 ;
        RECT 1194.260 213.560 1194.520 213.820 ;
      LAYER met2 ;
        RECT 1194.300 220.000 1194.580 224.000 ;
        RECT 1194.320 213.850 1194.460 220.000 ;
        RECT 1186.440 213.530 1186.700 213.850 ;
        RECT 1194.260 213.530 1194.520 213.850 ;
        RECT 1186.500 17.410 1186.640 213.530 ;
        RECT 1186.040 17.270 1186.640 17.410 ;
        RECT 1186.040 2.400 1186.180 17.270 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1203.890 20.640 1204.210 20.700 ;
        RECT 1207.110 20.640 1207.430 20.700 ;
        RECT 1203.890 20.500 1207.430 20.640 ;
        RECT 1203.890 20.440 1204.210 20.500 ;
        RECT 1207.110 20.440 1207.430 20.500 ;
      LAYER via ;
        RECT 1203.920 20.440 1204.180 20.700 ;
        RECT 1207.140 20.440 1207.400 20.700 ;
      LAYER met2 ;
        RECT 1209.020 220.730 1209.300 224.000 ;
        RECT 1208.120 220.590 1209.300 220.730 ;
        RECT 1208.120 213.930 1208.260 220.590 ;
        RECT 1209.020 220.000 1209.300 220.590 ;
        RECT 1207.200 213.790 1208.260 213.930 ;
        RECT 1207.200 20.730 1207.340 213.790 ;
        RECT 1203.920 20.410 1204.180 20.730 ;
        RECT 1207.140 20.410 1207.400 20.730 ;
        RECT 1203.980 2.400 1204.120 20.410 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1221.905 138.125 1222.075 186.235 ;
        RECT 1221.445 48.365 1221.615 113.815 ;
      LAYER mcon ;
        RECT 1221.905 186.065 1222.075 186.235 ;
        RECT 1221.445 113.645 1221.615 113.815 ;
      LAYER met1 ;
        RECT 1221.370 193.020 1221.690 193.080 ;
        RECT 1221.830 193.020 1222.150 193.080 ;
        RECT 1221.370 192.880 1222.150 193.020 ;
        RECT 1221.370 192.820 1221.690 192.880 ;
        RECT 1221.830 192.820 1222.150 192.880 ;
        RECT 1221.830 186.220 1222.150 186.280 ;
        RECT 1221.635 186.080 1222.150 186.220 ;
        RECT 1221.830 186.020 1222.150 186.080 ;
        RECT 1221.370 138.280 1221.690 138.340 ;
        RECT 1221.845 138.280 1222.135 138.325 ;
        RECT 1221.370 138.140 1222.135 138.280 ;
        RECT 1221.370 138.080 1221.690 138.140 ;
        RECT 1221.845 138.095 1222.135 138.140 ;
        RECT 1221.370 113.800 1221.690 113.860 ;
        RECT 1221.175 113.660 1221.690 113.800 ;
        RECT 1221.370 113.600 1221.690 113.660 ;
        RECT 1221.385 48.520 1221.675 48.565 ;
        RECT 1221.830 48.520 1222.150 48.580 ;
        RECT 1221.385 48.380 1222.150 48.520 ;
        RECT 1221.385 48.335 1221.675 48.380 ;
        RECT 1221.830 48.320 1222.150 48.380 ;
      LAYER via ;
        RECT 1221.400 192.820 1221.660 193.080 ;
        RECT 1221.860 192.820 1222.120 193.080 ;
        RECT 1221.860 186.020 1222.120 186.280 ;
        RECT 1221.400 138.080 1221.660 138.340 ;
        RECT 1221.400 113.600 1221.660 113.860 ;
        RECT 1221.860 48.320 1222.120 48.580 ;
      LAYER met2 ;
        RECT 1223.740 220.730 1224.020 224.000 ;
        RECT 1221.460 220.590 1224.020 220.730 ;
        RECT 1221.460 193.110 1221.600 220.590 ;
        RECT 1223.740 220.000 1224.020 220.590 ;
        RECT 1221.400 192.790 1221.660 193.110 ;
        RECT 1221.860 192.790 1222.120 193.110 ;
        RECT 1221.920 186.310 1222.060 192.790 ;
        RECT 1221.860 185.990 1222.120 186.310 ;
        RECT 1221.400 138.050 1221.660 138.370 ;
        RECT 1221.460 113.890 1221.600 138.050 ;
        RECT 1221.400 113.570 1221.660 113.890 ;
        RECT 1221.860 48.290 1222.120 48.610 ;
        RECT 1221.920 2.400 1222.060 48.290 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1235.170 20.640 1235.490 20.700 ;
        RECT 1239.770 20.640 1240.090 20.700 ;
        RECT 1235.170 20.500 1240.090 20.640 ;
        RECT 1235.170 20.440 1235.490 20.500 ;
        RECT 1239.770 20.440 1240.090 20.500 ;
      LAYER via ;
        RECT 1235.200 20.440 1235.460 20.700 ;
        RECT 1239.800 20.440 1240.060 20.700 ;
      LAYER met2 ;
        RECT 1238.460 220.730 1238.740 224.000 ;
        RECT 1235.260 220.590 1238.740 220.730 ;
        RECT 1235.260 20.730 1235.400 220.590 ;
        RECT 1238.460 220.000 1238.740 220.590 ;
        RECT 1235.200 20.410 1235.460 20.730 ;
        RECT 1239.800 20.410 1240.060 20.730 ;
        RECT 1239.860 2.400 1240.000 20.410 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1253.180 220.730 1253.460 224.000 ;
        RECT 1253.180 220.590 1255.640 220.730 ;
        RECT 1253.180 220.000 1253.460 220.590 ;
        RECT 1255.500 20.130 1255.640 220.590 ;
        RECT 1255.500 19.990 1257.480 20.130 ;
        RECT 1257.340 2.400 1257.480 19.990 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1270.130 2.960 1270.450 3.020 ;
        RECT 1275.190 2.960 1275.510 3.020 ;
        RECT 1270.130 2.820 1275.510 2.960 ;
        RECT 1270.130 2.760 1270.450 2.820 ;
        RECT 1275.190 2.760 1275.510 2.820 ;
      LAYER via ;
        RECT 1270.160 2.760 1270.420 3.020 ;
        RECT 1275.220 2.760 1275.480 3.020 ;
      LAYER met2 ;
        RECT 1267.900 220.730 1268.180 224.000 ;
        RECT 1267.900 220.590 1269.440 220.730 ;
        RECT 1267.900 220.000 1268.180 220.590 ;
        RECT 1269.300 207.130 1269.440 220.590 ;
        RECT 1269.300 206.990 1270.360 207.130 ;
        RECT 1270.220 3.050 1270.360 206.990 ;
        RECT 1270.160 2.730 1270.420 3.050 ;
        RECT 1275.220 2.730 1275.480 3.050 ;
        RECT 1275.280 2.400 1275.420 2.730 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1283.010 16.560 1283.330 16.620 ;
        RECT 1293.130 16.560 1293.450 16.620 ;
        RECT 1283.010 16.420 1293.450 16.560 ;
        RECT 1283.010 16.360 1283.330 16.420 ;
        RECT 1293.130 16.360 1293.450 16.420 ;
      LAYER via ;
        RECT 1283.040 16.360 1283.300 16.620 ;
        RECT 1293.160 16.360 1293.420 16.620 ;
      LAYER met2 ;
        RECT 1282.620 220.730 1282.900 224.000 ;
        RECT 1282.620 220.590 1283.240 220.730 ;
        RECT 1282.620 220.000 1282.900 220.590 ;
        RECT 1283.100 16.650 1283.240 220.590 ;
        RECT 1283.040 16.330 1283.300 16.650 ;
        RECT 1293.160 16.330 1293.420 16.650 ;
        RECT 1293.220 2.400 1293.360 16.330 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1297.270 207.300 1297.590 207.360 ;
        RECT 1307.390 207.300 1307.710 207.360 ;
        RECT 1297.270 207.160 1307.710 207.300 ;
        RECT 1297.270 207.100 1297.590 207.160 ;
        RECT 1307.390 207.100 1307.710 207.160 ;
        RECT 1307.390 17.580 1307.710 17.640 ;
        RECT 1311.070 17.580 1311.390 17.640 ;
        RECT 1307.390 17.440 1311.390 17.580 ;
        RECT 1307.390 17.380 1307.710 17.440 ;
        RECT 1311.070 17.380 1311.390 17.440 ;
      LAYER via ;
        RECT 1297.300 207.100 1297.560 207.360 ;
        RECT 1307.420 207.100 1307.680 207.360 ;
        RECT 1307.420 17.380 1307.680 17.640 ;
        RECT 1311.100 17.380 1311.360 17.640 ;
      LAYER met2 ;
        RECT 1297.340 220.000 1297.620 224.000 ;
        RECT 1297.360 207.390 1297.500 220.000 ;
        RECT 1297.300 207.070 1297.560 207.390 ;
        RECT 1307.420 207.070 1307.680 207.390 ;
        RECT 1307.480 17.670 1307.620 207.070 ;
        RECT 1307.420 17.350 1307.680 17.670 ;
        RECT 1311.100 17.350 1311.360 17.670 ;
        RECT 1311.160 2.400 1311.300 17.350 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.990 207.300 1312.310 207.360 ;
        RECT 1317.050 207.300 1317.370 207.360 ;
        RECT 1311.990 207.160 1317.370 207.300 ;
        RECT 1311.990 207.100 1312.310 207.160 ;
        RECT 1317.050 207.100 1317.370 207.160 ;
        RECT 1317.050 17.580 1317.370 17.640 ;
        RECT 1329.010 17.580 1329.330 17.640 ;
        RECT 1317.050 17.440 1329.330 17.580 ;
        RECT 1317.050 17.380 1317.370 17.440 ;
        RECT 1329.010 17.380 1329.330 17.440 ;
      LAYER via ;
        RECT 1312.020 207.100 1312.280 207.360 ;
        RECT 1317.080 207.100 1317.340 207.360 ;
        RECT 1317.080 17.380 1317.340 17.640 ;
        RECT 1329.040 17.380 1329.300 17.640 ;
      LAYER met2 ;
        RECT 1312.060 220.000 1312.340 224.000 ;
        RECT 1312.080 207.390 1312.220 220.000 ;
        RECT 1312.020 207.070 1312.280 207.390 ;
        RECT 1317.080 207.070 1317.340 207.390 ;
        RECT 1317.140 17.670 1317.280 207.070 ;
        RECT 1317.080 17.350 1317.340 17.670 ;
        RECT 1329.040 17.350 1329.300 17.670 ;
        RECT 1329.100 2.400 1329.240 17.350 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 689.610 209.340 689.930 209.400 ;
        RECT 782.990 209.340 783.310 209.400 ;
        RECT 689.610 209.200 783.310 209.340 ;
        RECT 689.610 209.140 689.930 209.200 ;
        RECT 782.990 209.140 783.310 209.200 ;
        RECT 686.390 17.580 686.710 17.640 ;
        RECT 689.610 17.580 689.930 17.640 ;
        RECT 686.390 17.440 689.930 17.580 ;
        RECT 686.390 17.380 686.710 17.440 ;
        RECT 689.610 17.380 689.930 17.440 ;
      LAYER via ;
        RECT 689.640 209.140 689.900 209.400 ;
        RECT 783.020 209.140 783.280 209.400 ;
        RECT 686.420 17.380 686.680 17.640 ;
        RECT 689.640 17.380 689.900 17.640 ;
      LAYER met2 ;
        RECT 783.060 220.000 783.340 224.000 ;
        RECT 783.080 209.430 783.220 220.000 ;
        RECT 689.640 209.110 689.900 209.430 ;
        RECT 783.020 209.110 783.280 209.430 ;
        RECT 689.700 17.670 689.840 209.110 ;
        RECT 686.420 17.350 686.680 17.670 ;
        RECT 689.640 17.350 689.900 17.670 ;
        RECT 686.480 2.400 686.620 17.350 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1326.710 207.300 1327.030 207.360 ;
        RECT 1330.850 207.300 1331.170 207.360 ;
        RECT 1326.710 207.160 1331.170 207.300 ;
        RECT 1326.710 207.100 1327.030 207.160 ;
        RECT 1330.850 207.100 1331.170 207.160 ;
        RECT 1330.850 17.240 1331.170 17.300 ;
        RECT 1346.490 17.240 1346.810 17.300 ;
        RECT 1330.850 17.100 1346.810 17.240 ;
        RECT 1330.850 17.040 1331.170 17.100 ;
        RECT 1346.490 17.040 1346.810 17.100 ;
      LAYER via ;
        RECT 1326.740 207.100 1327.000 207.360 ;
        RECT 1330.880 207.100 1331.140 207.360 ;
        RECT 1330.880 17.040 1331.140 17.300 ;
        RECT 1346.520 17.040 1346.780 17.300 ;
      LAYER met2 ;
        RECT 1326.780 220.000 1327.060 224.000 ;
        RECT 1326.800 207.390 1326.940 220.000 ;
        RECT 1326.740 207.070 1327.000 207.390 ;
        RECT 1330.880 207.070 1331.140 207.390 ;
        RECT 1330.940 17.330 1331.080 207.070 ;
        RECT 1330.880 17.010 1331.140 17.330 ;
        RECT 1346.520 17.010 1346.780 17.330 ;
        RECT 1346.580 2.400 1346.720 17.010 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1341.430 207.300 1341.750 207.360 ;
        RECT 1345.110 207.300 1345.430 207.360 ;
        RECT 1341.430 207.160 1345.430 207.300 ;
        RECT 1341.430 207.100 1341.750 207.160 ;
        RECT 1345.110 207.100 1345.430 207.160 ;
        RECT 1345.110 15.880 1345.430 15.940 ;
        RECT 1364.430 15.880 1364.750 15.940 ;
        RECT 1345.110 15.740 1364.750 15.880 ;
        RECT 1345.110 15.680 1345.430 15.740 ;
        RECT 1364.430 15.680 1364.750 15.740 ;
      LAYER via ;
        RECT 1341.460 207.100 1341.720 207.360 ;
        RECT 1345.140 207.100 1345.400 207.360 ;
        RECT 1345.140 15.680 1345.400 15.940 ;
        RECT 1364.460 15.680 1364.720 15.940 ;
      LAYER met2 ;
        RECT 1341.500 220.000 1341.780 224.000 ;
        RECT 1341.520 207.390 1341.660 220.000 ;
        RECT 1341.460 207.070 1341.720 207.390 ;
        RECT 1345.140 207.070 1345.400 207.390 ;
        RECT 1345.200 15.970 1345.340 207.070 ;
        RECT 1345.140 15.650 1345.400 15.970 ;
        RECT 1364.460 15.650 1364.720 15.970 ;
        RECT 1364.520 2.400 1364.660 15.650 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1356.150 207.640 1356.470 207.700 ;
        RECT 1362.590 207.640 1362.910 207.700 ;
        RECT 1356.150 207.500 1362.910 207.640 ;
        RECT 1356.150 207.440 1356.470 207.500 ;
        RECT 1362.590 207.440 1362.910 207.500 ;
        RECT 1362.590 16.560 1362.910 16.620 ;
        RECT 1382.370 16.560 1382.690 16.620 ;
        RECT 1362.590 16.420 1382.690 16.560 ;
        RECT 1362.590 16.360 1362.910 16.420 ;
        RECT 1382.370 16.360 1382.690 16.420 ;
      LAYER via ;
        RECT 1356.180 207.440 1356.440 207.700 ;
        RECT 1362.620 207.440 1362.880 207.700 ;
        RECT 1362.620 16.360 1362.880 16.620 ;
        RECT 1382.400 16.360 1382.660 16.620 ;
      LAYER met2 ;
        RECT 1356.220 220.000 1356.500 224.000 ;
        RECT 1356.240 207.730 1356.380 220.000 ;
        RECT 1356.180 207.410 1356.440 207.730 ;
        RECT 1362.620 207.410 1362.880 207.730 ;
        RECT 1362.680 16.650 1362.820 207.410 ;
        RECT 1362.620 16.330 1362.880 16.650 ;
        RECT 1382.400 16.330 1382.660 16.650 ;
        RECT 1382.460 2.400 1382.600 16.330 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1372.710 14.860 1373.030 14.920 ;
        RECT 1400.310 14.860 1400.630 14.920 ;
        RECT 1372.710 14.720 1400.630 14.860 ;
        RECT 1372.710 14.660 1373.030 14.720 ;
        RECT 1400.310 14.660 1400.630 14.720 ;
      LAYER via ;
        RECT 1372.740 14.660 1373.000 14.920 ;
        RECT 1400.340 14.660 1400.600 14.920 ;
      LAYER met2 ;
        RECT 1370.940 220.730 1371.220 224.000 ;
        RECT 1370.940 220.590 1372.940 220.730 ;
        RECT 1370.940 220.000 1371.220 220.590 ;
        RECT 1372.800 14.950 1372.940 220.590 ;
        RECT 1372.740 14.630 1373.000 14.950 ;
        RECT 1400.340 14.630 1400.600 14.950 ;
        RECT 1400.400 2.400 1400.540 14.630 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1386.050 17.240 1386.370 17.300 ;
        RECT 1418.250 17.240 1418.570 17.300 ;
        RECT 1386.050 17.100 1418.570 17.240 ;
        RECT 1386.050 17.040 1386.370 17.100 ;
        RECT 1418.250 17.040 1418.570 17.100 ;
      LAYER via ;
        RECT 1386.080 17.040 1386.340 17.300 ;
        RECT 1418.280 17.040 1418.540 17.300 ;
      LAYER met2 ;
        RECT 1385.200 220.730 1385.480 224.000 ;
        RECT 1385.200 220.590 1386.280 220.730 ;
        RECT 1385.200 220.000 1385.480 220.590 ;
        RECT 1386.140 17.330 1386.280 220.590 ;
        RECT 1386.080 17.010 1386.340 17.330 ;
        RECT 1418.280 17.010 1418.540 17.330 ;
        RECT 1418.340 2.400 1418.480 17.010 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1399.850 17.920 1400.170 17.980 ;
        RECT 1399.850 17.780 1430.440 17.920 ;
        RECT 1399.850 17.720 1400.170 17.780 ;
        RECT 1430.300 17.580 1430.440 17.780 ;
        RECT 1435.730 17.580 1436.050 17.640 ;
        RECT 1430.300 17.440 1436.050 17.580 ;
        RECT 1435.730 17.380 1436.050 17.440 ;
      LAYER via ;
        RECT 1399.880 17.720 1400.140 17.980 ;
        RECT 1435.760 17.380 1436.020 17.640 ;
      LAYER met2 ;
        RECT 1399.920 220.000 1400.200 224.000 ;
        RECT 1399.940 18.010 1400.080 220.000 ;
        RECT 1399.880 17.690 1400.140 18.010 ;
        RECT 1435.760 17.350 1436.020 17.670 ;
        RECT 1435.820 2.400 1435.960 17.350 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1414.570 207.300 1414.890 207.360 ;
        RECT 1420.550 207.300 1420.870 207.360 ;
        RECT 1414.570 207.160 1420.870 207.300 ;
        RECT 1414.570 207.100 1414.890 207.160 ;
        RECT 1420.550 207.100 1420.870 207.160 ;
        RECT 1420.550 18.260 1420.870 18.320 ;
        RECT 1453.670 18.260 1453.990 18.320 ;
        RECT 1420.550 18.120 1453.990 18.260 ;
        RECT 1420.550 18.060 1420.870 18.120 ;
        RECT 1453.670 18.060 1453.990 18.120 ;
      LAYER via ;
        RECT 1414.600 207.100 1414.860 207.360 ;
        RECT 1420.580 207.100 1420.840 207.360 ;
        RECT 1420.580 18.060 1420.840 18.320 ;
        RECT 1453.700 18.060 1453.960 18.320 ;
      LAYER met2 ;
        RECT 1414.640 220.000 1414.920 224.000 ;
        RECT 1414.660 207.390 1414.800 220.000 ;
        RECT 1414.600 207.070 1414.860 207.390 ;
        RECT 1420.580 207.070 1420.840 207.390 ;
        RECT 1420.640 18.350 1420.780 207.070 ;
        RECT 1420.580 18.030 1420.840 18.350 ;
        RECT 1453.700 18.030 1453.960 18.350 ;
        RECT 1453.760 2.400 1453.900 18.030 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1429.290 207.300 1429.610 207.360 ;
        RECT 1434.350 207.300 1434.670 207.360 ;
        RECT 1429.290 207.160 1434.670 207.300 ;
        RECT 1429.290 207.100 1429.610 207.160 ;
        RECT 1434.350 207.100 1434.670 207.160 ;
        RECT 1434.350 17.920 1434.670 17.980 ;
        RECT 1471.610 17.920 1471.930 17.980 ;
        RECT 1434.350 17.780 1471.930 17.920 ;
        RECT 1434.350 17.720 1434.670 17.780 ;
        RECT 1471.610 17.720 1471.930 17.780 ;
      LAYER via ;
        RECT 1429.320 207.100 1429.580 207.360 ;
        RECT 1434.380 207.100 1434.640 207.360 ;
        RECT 1434.380 17.720 1434.640 17.980 ;
        RECT 1471.640 17.720 1471.900 17.980 ;
      LAYER met2 ;
        RECT 1429.360 220.000 1429.640 224.000 ;
        RECT 1429.380 207.390 1429.520 220.000 ;
        RECT 1429.320 207.070 1429.580 207.390 ;
        RECT 1434.380 207.070 1434.640 207.390 ;
        RECT 1434.440 18.010 1434.580 207.070 ;
        RECT 1434.380 17.690 1434.640 18.010 ;
        RECT 1471.640 17.690 1471.900 18.010 ;
        RECT 1471.700 2.400 1471.840 17.690 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1444.010 207.300 1444.330 207.360 ;
        RECT 1448.610 207.300 1448.930 207.360 ;
        RECT 1444.010 207.160 1448.930 207.300 ;
        RECT 1444.010 207.100 1444.330 207.160 ;
        RECT 1448.610 207.100 1448.930 207.160 ;
        RECT 1448.610 20.300 1448.930 20.360 ;
        RECT 1489.550 20.300 1489.870 20.360 ;
        RECT 1448.610 20.160 1489.870 20.300 ;
        RECT 1448.610 20.100 1448.930 20.160 ;
        RECT 1489.550 20.100 1489.870 20.160 ;
      LAYER via ;
        RECT 1444.040 207.100 1444.300 207.360 ;
        RECT 1448.640 207.100 1448.900 207.360 ;
        RECT 1448.640 20.100 1448.900 20.360 ;
        RECT 1489.580 20.100 1489.840 20.360 ;
      LAYER met2 ;
        RECT 1444.080 220.000 1444.360 224.000 ;
        RECT 1444.100 207.390 1444.240 220.000 ;
        RECT 1444.040 207.070 1444.300 207.390 ;
        RECT 1448.640 207.070 1448.900 207.390 ;
        RECT 1448.700 20.390 1448.840 207.070 ;
        RECT 1448.640 20.070 1448.900 20.390 ;
        RECT 1489.580 20.070 1489.840 20.390 ;
        RECT 1489.640 2.400 1489.780 20.070 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1462.410 18.940 1462.730 19.000 ;
        RECT 1507.030 18.940 1507.350 19.000 ;
        RECT 1462.410 18.800 1507.350 18.940 ;
        RECT 1462.410 18.740 1462.730 18.800 ;
        RECT 1507.030 18.740 1507.350 18.800 ;
      LAYER via ;
        RECT 1462.440 18.740 1462.700 19.000 ;
        RECT 1507.060 18.740 1507.320 19.000 ;
      LAYER met2 ;
        RECT 1458.800 220.730 1459.080 224.000 ;
        RECT 1458.800 220.590 1462.640 220.730 ;
        RECT 1458.800 220.000 1459.080 220.590 ;
        RECT 1462.500 19.030 1462.640 220.590 ;
        RECT 1462.440 18.710 1462.700 19.030 ;
        RECT 1507.060 18.710 1507.320 19.030 ;
        RECT 1507.120 2.400 1507.260 18.710 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 709.850 212.060 710.170 212.120 ;
        RECT 797.710 212.060 798.030 212.120 ;
        RECT 709.850 211.920 798.030 212.060 ;
        RECT 709.850 211.860 710.170 211.920 ;
        RECT 797.710 211.860 798.030 211.920 ;
        RECT 704.330 17.580 704.650 17.640 ;
        RECT 709.850 17.580 710.170 17.640 ;
        RECT 704.330 17.440 710.170 17.580 ;
        RECT 704.330 17.380 704.650 17.440 ;
        RECT 709.850 17.380 710.170 17.440 ;
      LAYER via ;
        RECT 709.880 211.860 710.140 212.120 ;
        RECT 797.740 211.860 798.000 212.120 ;
        RECT 704.360 17.380 704.620 17.640 ;
        RECT 709.880 17.380 710.140 17.640 ;
      LAYER met2 ;
        RECT 797.780 220.000 798.060 224.000 ;
        RECT 797.800 212.150 797.940 220.000 ;
        RECT 709.880 211.830 710.140 212.150 ;
        RECT 797.740 211.830 798.000 212.150 ;
        RECT 709.940 17.670 710.080 211.830 ;
        RECT 704.360 17.350 704.620 17.670 ;
        RECT 709.880 17.350 710.140 17.670 ;
        RECT 704.420 2.400 704.560 17.350 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1476.210 19.960 1476.530 20.020 ;
        RECT 1524.970 19.960 1525.290 20.020 ;
        RECT 1476.210 19.820 1525.290 19.960 ;
        RECT 1476.210 19.760 1476.530 19.820 ;
        RECT 1524.970 19.760 1525.290 19.820 ;
      LAYER via ;
        RECT 1476.240 19.760 1476.500 20.020 ;
        RECT 1525.000 19.760 1525.260 20.020 ;
      LAYER met2 ;
        RECT 1473.520 220.730 1473.800 224.000 ;
        RECT 1473.520 220.590 1476.440 220.730 ;
        RECT 1473.520 220.000 1473.800 220.590 ;
        RECT 1476.300 20.050 1476.440 220.590 ;
        RECT 1476.240 19.730 1476.500 20.050 ;
        RECT 1525.000 19.730 1525.260 20.050 ;
        RECT 1525.060 2.400 1525.200 19.730 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1490.010 17.920 1490.330 17.980 ;
        RECT 1542.910 17.920 1543.230 17.980 ;
        RECT 1490.010 17.780 1543.230 17.920 ;
        RECT 1490.010 17.720 1490.330 17.780 ;
        RECT 1542.910 17.720 1543.230 17.780 ;
      LAYER via ;
        RECT 1490.040 17.720 1490.300 17.980 ;
        RECT 1542.940 17.720 1543.200 17.980 ;
      LAYER met2 ;
        RECT 1488.240 220.730 1488.520 224.000 ;
        RECT 1488.240 220.590 1490.240 220.730 ;
        RECT 1488.240 220.000 1488.520 220.590 ;
        RECT 1490.100 18.010 1490.240 220.590 ;
        RECT 1490.040 17.690 1490.300 18.010 ;
        RECT 1542.940 17.690 1543.200 18.010 ;
        RECT 1543.000 2.400 1543.140 17.690 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1503.350 18.600 1503.670 18.660 ;
        RECT 1560.850 18.600 1561.170 18.660 ;
        RECT 1503.350 18.460 1561.170 18.600 ;
        RECT 1503.350 18.400 1503.670 18.460 ;
        RECT 1560.850 18.400 1561.170 18.460 ;
      LAYER via ;
        RECT 1503.380 18.400 1503.640 18.660 ;
        RECT 1560.880 18.400 1561.140 18.660 ;
      LAYER met2 ;
        RECT 1502.960 220.730 1503.240 224.000 ;
        RECT 1502.960 220.590 1503.580 220.730 ;
        RECT 1502.960 220.000 1503.240 220.590 ;
        RECT 1503.440 18.690 1503.580 220.590 ;
        RECT 1503.380 18.370 1503.640 18.690 ;
        RECT 1560.880 18.370 1561.140 18.690 ;
        RECT 1560.940 2.400 1561.080 18.370 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1517.150 19.280 1517.470 19.340 ;
        RECT 1578.790 19.280 1579.110 19.340 ;
        RECT 1517.150 19.140 1579.110 19.280 ;
        RECT 1517.150 19.080 1517.470 19.140 ;
        RECT 1578.790 19.080 1579.110 19.140 ;
      LAYER via ;
        RECT 1517.180 19.080 1517.440 19.340 ;
        RECT 1578.820 19.080 1579.080 19.340 ;
      LAYER met2 ;
        RECT 1517.680 220.730 1517.960 224.000 ;
        RECT 1517.240 220.590 1517.960 220.730 ;
        RECT 1517.240 19.370 1517.380 220.590 ;
        RECT 1517.680 220.000 1517.960 220.590 ;
        RECT 1517.180 19.050 1517.440 19.370 ;
        RECT 1578.820 19.050 1579.080 19.370 ;
        RECT 1578.880 2.400 1579.020 19.050 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1532.330 207.300 1532.650 207.360 ;
        RECT 1537.850 207.300 1538.170 207.360 ;
        RECT 1532.330 207.160 1538.170 207.300 ;
        RECT 1532.330 207.100 1532.650 207.160 ;
        RECT 1537.850 207.100 1538.170 207.160 ;
        RECT 1537.850 19.960 1538.170 20.020 ;
        RECT 1596.270 19.960 1596.590 20.020 ;
        RECT 1537.850 19.820 1596.590 19.960 ;
        RECT 1537.850 19.760 1538.170 19.820 ;
        RECT 1596.270 19.760 1596.590 19.820 ;
      LAYER via ;
        RECT 1532.360 207.100 1532.620 207.360 ;
        RECT 1537.880 207.100 1538.140 207.360 ;
        RECT 1537.880 19.760 1538.140 20.020 ;
        RECT 1596.300 19.760 1596.560 20.020 ;
      LAYER met2 ;
        RECT 1532.400 220.000 1532.680 224.000 ;
        RECT 1532.420 207.390 1532.560 220.000 ;
        RECT 1532.360 207.070 1532.620 207.390 ;
        RECT 1537.880 207.070 1538.140 207.390 ;
        RECT 1537.940 20.050 1538.080 207.070 ;
        RECT 1537.880 19.730 1538.140 20.050 ;
        RECT 1596.300 19.730 1596.560 20.050 ;
        RECT 1596.360 2.400 1596.500 19.730 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1547.050 207.300 1547.370 207.360 ;
        RECT 1551.650 207.300 1551.970 207.360 ;
        RECT 1547.050 207.160 1551.970 207.300 ;
        RECT 1547.050 207.100 1547.370 207.160 ;
        RECT 1551.650 207.100 1551.970 207.160 ;
        RECT 1551.650 20.300 1551.970 20.360 ;
        RECT 1613.750 20.300 1614.070 20.360 ;
        RECT 1551.650 20.160 1614.070 20.300 ;
        RECT 1551.650 20.100 1551.970 20.160 ;
        RECT 1613.750 20.100 1614.070 20.160 ;
      LAYER via ;
        RECT 1547.080 207.100 1547.340 207.360 ;
        RECT 1551.680 207.100 1551.940 207.360 ;
        RECT 1551.680 20.100 1551.940 20.360 ;
        RECT 1613.780 20.100 1614.040 20.360 ;
      LAYER met2 ;
        RECT 1547.120 220.000 1547.400 224.000 ;
        RECT 1547.140 207.390 1547.280 220.000 ;
        RECT 1547.080 207.070 1547.340 207.390 ;
        RECT 1551.680 207.070 1551.940 207.390 ;
        RECT 1551.740 20.390 1551.880 207.070 ;
        RECT 1551.680 20.070 1551.940 20.390 ;
        RECT 1613.780 20.070 1614.040 20.390 ;
        RECT 1613.840 17.410 1613.980 20.070 ;
        RECT 1613.840 17.270 1614.440 17.410 ;
        RECT 1614.300 2.400 1614.440 17.270 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1561.770 207.300 1562.090 207.360 ;
        RECT 1565.910 207.300 1566.230 207.360 ;
        RECT 1561.770 207.160 1566.230 207.300 ;
        RECT 1561.770 207.100 1562.090 207.160 ;
        RECT 1565.910 207.100 1566.230 207.160 ;
        RECT 1565.910 19.620 1566.230 19.680 ;
        RECT 1632.150 19.620 1632.470 19.680 ;
        RECT 1565.910 19.480 1632.470 19.620 ;
        RECT 1565.910 19.420 1566.230 19.480 ;
        RECT 1632.150 19.420 1632.470 19.480 ;
      LAYER via ;
        RECT 1561.800 207.100 1562.060 207.360 ;
        RECT 1565.940 207.100 1566.200 207.360 ;
        RECT 1565.940 19.420 1566.200 19.680 ;
        RECT 1632.180 19.420 1632.440 19.680 ;
      LAYER met2 ;
        RECT 1561.840 220.000 1562.120 224.000 ;
        RECT 1561.860 207.390 1562.000 220.000 ;
        RECT 1561.800 207.070 1562.060 207.390 ;
        RECT 1565.940 207.070 1566.200 207.390 ;
        RECT 1566.000 19.710 1566.140 207.070 ;
        RECT 1565.940 19.390 1566.200 19.710 ;
        RECT 1632.180 19.390 1632.440 19.710 ;
        RECT 1632.240 2.400 1632.380 19.390 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1579.710 19.280 1580.030 19.340 ;
        RECT 1650.090 19.280 1650.410 19.340 ;
        RECT 1579.710 19.140 1650.410 19.280 ;
        RECT 1579.710 19.080 1580.030 19.140 ;
        RECT 1650.090 19.080 1650.410 19.140 ;
      LAYER via ;
        RECT 1579.740 19.080 1580.000 19.340 ;
        RECT 1650.120 19.080 1650.380 19.340 ;
      LAYER met2 ;
        RECT 1576.560 220.730 1576.840 224.000 ;
        RECT 1576.560 220.590 1579.940 220.730 ;
        RECT 1576.560 220.000 1576.840 220.590 ;
        RECT 1579.800 19.370 1579.940 220.590 ;
        RECT 1579.740 19.050 1580.000 19.370 ;
        RECT 1650.120 19.050 1650.380 19.370 ;
        RECT 1650.180 2.400 1650.320 19.050 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1593.510 15.880 1593.830 15.940 ;
        RECT 1668.030 15.880 1668.350 15.940 ;
        RECT 1593.510 15.740 1668.350 15.880 ;
        RECT 1593.510 15.680 1593.830 15.740 ;
        RECT 1668.030 15.680 1668.350 15.740 ;
      LAYER via ;
        RECT 1593.540 15.680 1593.800 15.940 ;
        RECT 1668.060 15.680 1668.320 15.940 ;
      LAYER met2 ;
        RECT 1591.280 220.730 1591.560 224.000 ;
        RECT 1591.280 220.590 1593.740 220.730 ;
        RECT 1591.280 220.000 1591.560 220.590 ;
        RECT 1593.600 15.970 1593.740 220.590 ;
        RECT 1593.540 15.650 1593.800 15.970 ;
        RECT 1668.060 15.650 1668.320 15.970 ;
        RECT 1668.120 2.400 1668.260 15.650 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1606.850 17.240 1607.170 17.300 ;
        RECT 1685.510 17.240 1685.830 17.300 ;
        RECT 1606.850 17.100 1685.830 17.240 ;
        RECT 1606.850 17.040 1607.170 17.100 ;
        RECT 1685.510 17.040 1685.830 17.100 ;
      LAYER via ;
        RECT 1606.880 17.040 1607.140 17.300 ;
        RECT 1685.540 17.040 1685.800 17.300 ;
      LAYER met2 ;
        RECT 1606.000 220.730 1606.280 224.000 ;
        RECT 1606.000 220.590 1607.080 220.730 ;
        RECT 1606.000 220.000 1606.280 220.590 ;
        RECT 1606.940 17.330 1607.080 220.590 ;
        RECT 1606.880 17.010 1607.140 17.330 ;
        RECT 1685.540 17.010 1685.800 17.330 ;
        RECT 1685.600 2.400 1685.740 17.010 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 723.190 212.740 723.510 212.800 ;
        RECT 812.430 212.740 812.750 212.800 ;
        RECT 723.190 212.600 812.750 212.740 ;
        RECT 723.190 212.540 723.510 212.600 ;
        RECT 812.430 212.540 812.750 212.600 ;
      LAYER via ;
        RECT 723.220 212.540 723.480 212.800 ;
        RECT 812.460 212.540 812.720 212.800 ;
      LAYER met2 ;
        RECT 812.500 220.000 812.780 224.000 ;
        RECT 812.520 212.830 812.660 220.000 ;
        RECT 723.220 212.510 723.480 212.830 ;
        RECT 812.460 212.510 812.720 212.830 ;
        RECT 723.280 196.250 723.420 212.510 ;
        RECT 723.280 196.110 724.340 196.250 ;
        RECT 724.200 16.730 724.340 196.110 ;
        RECT 722.360 16.590 724.340 16.730 ;
        RECT 722.360 2.400 722.500 16.590 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1620.650 17.580 1620.970 17.640 ;
        RECT 1703.450 17.580 1703.770 17.640 ;
        RECT 1620.650 17.440 1703.770 17.580 ;
        RECT 1620.650 17.380 1620.970 17.440 ;
        RECT 1703.450 17.380 1703.770 17.440 ;
      LAYER via ;
        RECT 1620.680 17.380 1620.940 17.640 ;
        RECT 1703.480 17.380 1703.740 17.640 ;
      LAYER met2 ;
        RECT 1620.720 220.000 1621.000 224.000 ;
        RECT 1620.740 17.670 1620.880 220.000 ;
        RECT 1620.680 17.350 1620.940 17.670 ;
        RECT 1703.480 17.350 1703.740 17.670 ;
        RECT 1703.540 2.400 1703.680 17.350 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1634.910 19.960 1635.230 20.020 ;
        RECT 1721.390 19.960 1721.710 20.020 ;
        RECT 1634.910 19.820 1721.710 19.960 ;
        RECT 1634.910 19.760 1635.230 19.820 ;
        RECT 1721.390 19.760 1721.710 19.820 ;
      LAYER via ;
        RECT 1634.940 19.760 1635.200 20.020 ;
        RECT 1721.420 19.760 1721.680 20.020 ;
      LAYER met2 ;
        RECT 1634.980 220.000 1635.260 224.000 ;
        RECT 1635.000 20.050 1635.140 220.000 ;
        RECT 1634.940 19.730 1635.200 20.050 ;
        RECT 1721.420 19.730 1721.680 20.050 ;
        RECT 1721.480 2.400 1721.620 19.730 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1649.630 207.300 1649.950 207.360 ;
        RECT 1655.150 207.300 1655.470 207.360 ;
        RECT 1649.630 207.160 1655.470 207.300 ;
        RECT 1649.630 207.100 1649.950 207.160 ;
        RECT 1655.150 207.100 1655.470 207.160 ;
        RECT 1655.150 19.620 1655.470 19.680 ;
        RECT 1739.330 19.620 1739.650 19.680 ;
        RECT 1655.150 19.480 1739.650 19.620 ;
        RECT 1655.150 19.420 1655.470 19.480 ;
        RECT 1739.330 19.420 1739.650 19.480 ;
      LAYER via ;
        RECT 1649.660 207.100 1649.920 207.360 ;
        RECT 1655.180 207.100 1655.440 207.360 ;
        RECT 1655.180 19.420 1655.440 19.680 ;
        RECT 1739.360 19.420 1739.620 19.680 ;
      LAYER met2 ;
        RECT 1649.700 220.000 1649.980 224.000 ;
        RECT 1649.720 207.390 1649.860 220.000 ;
        RECT 1649.660 207.070 1649.920 207.390 ;
        RECT 1655.180 207.070 1655.440 207.390 ;
        RECT 1655.240 19.710 1655.380 207.070 ;
        RECT 1655.180 19.390 1655.440 19.710 ;
        RECT 1739.360 19.390 1739.620 19.710 ;
        RECT 1739.420 2.400 1739.560 19.390 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1664.350 207.300 1664.670 207.360 ;
        RECT 1668.950 207.300 1669.270 207.360 ;
        RECT 1664.350 207.160 1669.270 207.300 ;
        RECT 1664.350 207.100 1664.670 207.160 ;
        RECT 1668.950 207.100 1669.270 207.160 ;
        RECT 1668.950 16.560 1669.270 16.620 ;
        RECT 1756.810 16.560 1757.130 16.620 ;
        RECT 1668.950 16.420 1757.130 16.560 ;
        RECT 1668.950 16.360 1669.270 16.420 ;
        RECT 1756.810 16.360 1757.130 16.420 ;
      LAYER via ;
        RECT 1664.380 207.100 1664.640 207.360 ;
        RECT 1668.980 207.100 1669.240 207.360 ;
        RECT 1668.980 16.360 1669.240 16.620 ;
        RECT 1756.840 16.360 1757.100 16.620 ;
      LAYER met2 ;
        RECT 1664.420 220.000 1664.700 224.000 ;
        RECT 1664.440 207.390 1664.580 220.000 ;
        RECT 1664.380 207.070 1664.640 207.390 ;
        RECT 1668.980 207.070 1669.240 207.390 ;
        RECT 1669.040 16.650 1669.180 207.070 ;
        RECT 1668.980 16.330 1669.240 16.650 ;
        RECT 1756.840 16.330 1757.100 16.650 ;
        RECT 1756.900 2.400 1757.040 16.330 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1679.070 207.300 1679.390 207.360 ;
        RECT 1683.210 207.300 1683.530 207.360 ;
        RECT 1679.070 207.160 1683.530 207.300 ;
        RECT 1679.070 207.100 1679.390 207.160 ;
        RECT 1683.210 207.100 1683.530 207.160 ;
        RECT 1683.210 19.280 1683.530 19.340 ;
        RECT 1774.750 19.280 1775.070 19.340 ;
        RECT 1683.210 19.140 1775.070 19.280 ;
        RECT 1683.210 19.080 1683.530 19.140 ;
        RECT 1774.750 19.080 1775.070 19.140 ;
      LAYER via ;
        RECT 1679.100 207.100 1679.360 207.360 ;
        RECT 1683.240 207.100 1683.500 207.360 ;
        RECT 1683.240 19.080 1683.500 19.340 ;
        RECT 1774.780 19.080 1775.040 19.340 ;
      LAYER met2 ;
        RECT 1679.140 220.000 1679.420 224.000 ;
        RECT 1679.160 207.390 1679.300 220.000 ;
        RECT 1679.100 207.070 1679.360 207.390 ;
        RECT 1683.240 207.070 1683.500 207.390 ;
        RECT 1683.300 19.370 1683.440 207.070 ;
        RECT 1683.240 19.050 1683.500 19.370 ;
        RECT 1774.780 19.050 1775.040 19.370 ;
        RECT 1774.840 2.400 1774.980 19.050 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1697.010 17.920 1697.330 17.980 ;
        RECT 1792.690 17.920 1793.010 17.980 ;
        RECT 1697.010 17.780 1793.010 17.920 ;
        RECT 1697.010 17.720 1697.330 17.780 ;
        RECT 1792.690 17.720 1793.010 17.780 ;
      LAYER via ;
        RECT 1697.040 17.720 1697.300 17.980 ;
        RECT 1792.720 17.720 1792.980 17.980 ;
      LAYER met2 ;
        RECT 1693.860 220.730 1694.140 224.000 ;
        RECT 1693.860 220.590 1697.240 220.730 ;
        RECT 1693.860 220.000 1694.140 220.590 ;
        RECT 1697.100 18.010 1697.240 220.590 ;
        RECT 1697.040 17.690 1697.300 18.010 ;
        RECT 1792.720 17.690 1792.980 18.010 ;
        RECT 1792.780 2.400 1792.920 17.690 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1710.810 16.220 1711.130 16.280 ;
        RECT 1810.630 16.220 1810.950 16.280 ;
        RECT 1710.810 16.080 1810.950 16.220 ;
        RECT 1710.810 16.020 1711.130 16.080 ;
        RECT 1810.630 16.020 1810.950 16.080 ;
      LAYER via ;
        RECT 1710.840 16.020 1711.100 16.280 ;
        RECT 1810.660 16.020 1810.920 16.280 ;
      LAYER met2 ;
        RECT 1708.580 220.730 1708.860 224.000 ;
        RECT 1708.580 220.590 1711.040 220.730 ;
        RECT 1708.580 220.000 1708.860 220.590 ;
        RECT 1710.900 16.310 1711.040 220.590 ;
        RECT 1710.840 15.990 1711.100 16.310 ;
        RECT 1810.660 15.990 1810.920 16.310 ;
        RECT 1810.720 2.400 1810.860 15.990 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1723.230 210.700 1723.550 210.760 ;
        RECT 1829.030 210.700 1829.350 210.760 ;
        RECT 1723.230 210.560 1829.350 210.700 ;
        RECT 1723.230 210.500 1723.550 210.560 ;
        RECT 1829.030 210.500 1829.350 210.560 ;
      LAYER via ;
        RECT 1723.260 210.500 1723.520 210.760 ;
        RECT 1829.060 210.500 1829.320 210.760 ;
      LAYER met2 ;
        RECT 1723.300 220.000 1723.580 224.000 ;
        RECT 1723.320 210.790 1723.460 220.000 ;
        RECT 1723.260 210.470 1723.520 210.790 ;
        RECT 1829.060 210.470 1829.320 210.790 ;
        RECT 1829.120 17.410 1829.260 210.470 ;
        RECT 1828.660 17.270 1829.260 17.410 ;
        RECT 1828.660 2.400 1828.800 17.270 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1737.950 212.740 1738.270 212.800 ;
        RECT 1842.830 212.740 1843.150 212.800 ;
        RECT 1737.950 212.600 1843.150 212.740 ;
        RECT 1737.950 212.540 1738.270 212.600 ;
        RECT 1842.830 212.540 1843.150 212.600 ;
        RECT 1842.830 2.960 1843.150 3.020 ;
        RECT 1846.050 2.960 1846.370 3.020 ;
        RECT 1842.830 2.820 1846.370 2.960 ;
        RECT 1842.830 2.760 1843.150 2.820 ;
        RECT 1846.050 2.760 1846.370 2.820 ;
      LAYER via ;
        RECT 1737.980 212.540 1738.240 212.800 ;
        RECT 1842.860 212.540 1843.120 212.800 ;
        RECT 1842.860 2.760 1843.120 3.020 ;
        RECT 1846.080 2.760 1846.340 3.020 ;
      LAYER met2 ;
        RECT 1738.020 220.000 1738.300 224.000 ;
        RECT 1738.040 212.830 1738.180 220.000 ;
        RECT 1737.980 212.510 1738.240 212.830 ;
        RECT 1842.860 212.510 1843.120 212.830 ;
        RECT 1842.920 3.050 1843.060 212.510 ;
        RECT 1842.860 2.730 1843.120 3.050 ;
        RECT 1846.080 2.730 1846.340 3.050 ;
        RECT 1846.140 2.400 1846.280 2.730 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1752.670 210.360 1752.990 210.420 ;
        RECT 1863.530 210.360 1863.850 210.420 ;
        RECT 1752.670 210.220 1863.850 210.360 ;
        RECT 1752.670 210.160 1752.990 210.220 ;
        RECT 1863.530 210.160 1863.850 210.220 ;
      LAYER via ;
        RECT 1752.700 210.160 1752.960 210.420 ;
        RECT 1863.560 210.160 1863.820 210.420 ;
      LAYER met2 ;
        RECT 1752.740 220.000 1753.020 224.000 ;
        RECT 1752.760 210.450 1752.900 220.000 ;
        RECT 1752.700 210.130 1752.960 210.450 ;
        RECT 1863.560 210.130 1863.820 210.450 ;
        RECT 1863.620 17.410 1863.760 210.130 ;
        RECT 1863.620 17.270 1864.220 17.410 ;
        RECT 1864.080 2.400 1864.220 17.270 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 744.810 209.000 745.130 209.060 ;
        RECT 827.150 209.000 827.470 209.060 ;
        RECT 744.810 208.860 827.470 209.000 ;
        RECT 744.810 208.800 745.130 208.860 ;
        RECT 827.150 208.800 827.470 208.860 ;
        RECT 740.210 17.580 740.530 17.640 ;
        RECT 744.810 17.580 745.130 17.640 ;
        RECT 740.210 17.440 745.130 17.580 ;
        RECT 740.210 17.380 740.530 17.440 ;
        RECT 744.810 17.380 745.130 17.440 ;
      LAYER via ;
        RECT 744.840 208.800 745.100 209.060 ;
        RECT 827.180 208.800 827.440 209.060 ;
        RECT 740.240 17.380 740.500 17.640 ;
        RECT 744.840 17.380 745.100 17.640 ;
      LAYER met2 ;
        RECT 827.220 220.000 827.500 224.000 ;
        RECT 827.240 209.090 827.380 220.000 ;
        RECT 744.840 208.770 745.100 209.090 ;
        RECT 827.180 208.770 827.440 209.090 ;
        RECT 744.900 17.670 745.040 208.770 ;
        RECT 740.240 17.350 740.500 17.670 ;
        RECT 744.840 17.350 745.100 17.670 ;
        RECT 740.300 2.400 740.440 17.350 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1767.390 212.060 1767.710 212.120 ;
        RECT 1877.330 212.060 1877.650 212.120 ;
        RECT 1767.390 211.920 1877.650 212.060 ;
        RECT 1767.390 211.860 1767.710 211.920 ;
        RECT 1877.330 211.860 1877.650 211.920 ;
        RECT 1877.330 2.960 1877.650 3.020 ;
        RECT 1881.930 2.960 1882.250 3.020 ;
        RECT 1877.330 2.820 1882.250 2.960 ;
        RECT 1877.330 2.760 1877.650 2.820 ;
        RECT 1881.930 2.760 1882.250 2.820 ;
      LAYER via ;
        RECT 1767.420 211.860 1767.680 212.120 ;
        RECT 1877.360 211.860 1877.620 212.120 ;
        RECT 1877.360 2.760 1877.620 3.020 ;
        RECT 1881.960 2.760 1882.220 3.020 ;
      LAYER met2 ;
        RECT 1767.460 220.000 1767.740 224.000 ;
        RECT 1767.480 212.150 1767.620 220.000 ;
        RECT 1767.420 211.830 1767.680 212.150 ;
        RECT 1877.360 211.830 1877.620 212.150 ;
        RECT 1877.420 3.050 1877.560 211.830 ;
        RECT 1877.360 2.730 1877.620 3.050 ;
        RECT 1881.960 2.730 1882.220 3.050 ;
        RECT 1882.020 2.400 1882.160 2.730 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1782.110 211.720 1782.430 211.780 ;
        RECT 1897.570 211.720 1897.890 211.780 ;
        RECT 1782.110 211.580 1897.890 211.720 ;
        RECT 1782.110 211.520 1782.430 211.580 ;
        RECT 1897.570 211.520 1897.890 211.580 ;
        RECT 1897.570 2.960 1897.890 3.020 ;
        RECT 1899.870 2.960 1900.190 3.020 ;
        RECT 1897.570 2.820 1900.190 2.960 ;
        RECT 1897.570 2.760 1897.890 2.820 ;
        RECT 1899.870 2.760 1900.190 2.820 ;
      LAYER via ;
        RECT 1782.140 211.520 1782.400 211.780 ;
        RECT 1897.600 211.520 1897.860 211.780 ;
        RECT 1897.600 2.760 1897.860 3.020 ;
        RECT 1899.900 2.760 1900.160 3.020 ;
      LAYER met2 ;
        RECT 1782.180 220.000 1782.460 224.000 ;
        RECT 1782.200 211.810 1782.340 220.000 ;
        RECT 1782.140 211.490 1782.400 211.810 ;
        RECT 1897.600 211.490 1897.860 211.810 ;
        RECT 1897.660 3.050 1897.800 211.490 ;
        RECT 1897.600 2.730 1897.860 3.050 ;
        RECT 1899.900 2.730 1900.160 3.050 ;
        RECT 1899.960 2.400 1900.100 2.730 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1796.830 212.400 1797.150 212.460 ;
        RECT 1912.290 212.400 1912.610 212.460 ;
        RECT 1796.830 212.260 1912.610 212.400 ;
        RECT 1796.830 212.200 1797.150 212.260 ;
        RECT 1912.290 212.200 1912.610 212.260 ;
        RECT 1912.290 2.960 1912.610 3.020 ;
        RECT 1917.810 2.960 1918.130 3.020 ;
        RECT 1912.290 2.820 1918.130 2.960 ;
        RECT 1912.290 2.760 1912.610 2.820 ;
        RECT 1917.810 2.760 1918.130 2.820 ;
      LAYER via ;
        RECT 1796.860 212.200 1797.120 212.460 ;
        RECT 1912.320 212.200 1912.580 212.460 ;
        RECT 1912.320 2.760 1912.580 3.020 ;
        RECT 1917.840 2.760 1918.100 3.020 ;
      LAYER met2 ;
        RECT 1796.900 220.000 1797.180 224.000 ;
        RECT 1796.920 212.490 1797.060 220.000 ;
        RECT 1796.860 212.170 1797.120 212.490 ;
        RECT 1912.320 212.170 1912.580 212.490 ;
        RECT 1912.380 3.050 1912.520 212.170 ;
        RECT 1912.320 2.730 1912.580 3.050 ;
        RECT 1917.840 2.730 1918.100 3.050 ;
        RECT 1917.900 2.400 1918.040 2.730 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1811.550 211.380 1811.870 211.440 ;
        RECT 1932.530 211.380 1932.850 211.440 ;
        RECT 1811.550 211.240 1932.850 211.380 ;
        RECT 1811.550 211.180 1811.870 211.240 ;
        RECT 1932.530 211.180 1932.850 211.240 ;
        RECT 1932.530 2.960 1932.850 3.020 ;
        RECT 1935.290 2.960 1935.610 3.020 ;
        RECT 1932.530 2.820 1935.610 2.960 ;
        RECT 1932.530 2.760 1932.850 2.820 ;
        RECT 1935.290 2.760 1935.610 2.820 ;
      LAYER via ;
        RECT 1811.580 211.180 1811.840 211.440 ;
        RECT 1932.560 211.180 1932.820 211.440 ;
        RECT 1932.560 2.760 1932.820 3.020 ;
        RECT 1935.320 2.760 1935.580 3.020 ;
      LAYER met2 ;
        RECT 1811.620 220.000 1811.900 224.000 ;
        RECT 1811.640 211.470 1811.780 220.000 ;
        RECT 1811.580 211.150 1811.840 211.470 ;
        RECT 1932.560 211.150 1932.820 211.470 ;
        RECT 1932.620 3.050 1932.760 211.150 ;
        RECT 1932.560 2.730 1932.820 3.050 ;
        RECT 1935.320 2.730 1935.580 3.050 ;
        RECT 1935.380 2.400 1935.520 2.730 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1826.270 213.080 1826.590 213.140 ;
        RECT 1953.230 213.080 1953.550 213.140 ;
        RECT 1826.270 212.940 1953.550 213.080 ;
        RECT 1826.270 212.880 1826.590 212.940 ;
        RECT 1953.230 212.880 1953.550 212.940 ;
      LAYER via ;
        RECT 1826.300 212.880 1826.560 213.140 ;
        RECT 1953.260 212.880 1953.520 213.140 ;
      LAYER met2 ;
        RECT 1826.340 220.000 1826.620 224.000 ;
        RECT 1826.360 213.170 1826.500 220.000 ;
        RECT 1826.300 212.850 1826.560 213.170 ;
        RECT 1953.260 212.850 1953.520 213.170 ;
        RECT 1953.320 2.400 1953.460 212.850 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1840.990 211.040 1841.310 211.100 ;
        RECT 1967.490 211.040 1967.810 211.100 ;
        RECT 1840.990 210.900 1967.810 211.040 ;
        RECT 1840.990 210.840 1841.310 210.900 ;
        RECT 1967.490 210.840 1967.810 210.900 ;
        RECT 1967.490 2.960 1967.810 3.020 ;
        RECT 1971.170 2.960 1971.490 3.020 ;
        RECT 1967.490 2.820 1971.490 2.960 ;
        RECT 1967.490 2.760 1967.810 2.820 ;
        RECT 1971.170 2.760 1971.490 2.820 ;
      LAYER via ;
        RECT 1841.020 210.840 1841.280 211.100 ;
        RECT 1967.520 210.840 1967.780 211.100 ;
        RECT 1967.520 2.760 1967.780 3.020 ;
        RECT 1971.200 2.760 1971.460 3.020 ;
      LAYER met2 ;
        RECT 1841.060 220.000 1841.340 224.000 ;
        RECT 1841.080 211.130 1841.220 220.000 ;
        RECT 1841.020 210.810 1841.280 211.130 ;
        RECT 1967.520 210.810 1967.780 211.130 ;
        RECT 1967.580 3.050 1967.720 210.810 ;
        RECT 1967.520 2.730 1967.780 3.050 ;
        RECT 1971.200 2.730 1971.460 3.050 ;
        RECT 1971.260 2.400 1971.400 2.730 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1855.710 210.700 1856.030 210.760 ;
        RECT 1988.190 210.700 1988.510 210.760 ;
        RECT 1855.710 210.560 1988.510 210.700 ;
        RECT 1855.710 210.500 1856.030 210.560 ;
        RECT 1988.190 210.500 1988.510 210.560 ;
        RECT 1988.190 2.960 1988.510 3.020 ;
        RECT 1989.110 2.960 1989.430 3.020 ;
        RECT 1988.190 2.820 1989.430 2.960 ;
        RECT 1988.190 2.760 1988.510 2.820 ;
        RECT 1989.110 2.760 1989.430 2.820 ;
      LAYER via ;
        RECT 1855.740 210.500 1856.000 210.760 ;
        RECT 1988.220 210.500 1988.480 210.760 ;
        RECT 1988.220 2.760 1988.480 3.020 ;
        RECT 1989.140 2.760 1989.400 3.020 ;
      LAYER met2 ;
        RECT 1855.780 220.000 1856.060 224.000 ;
        RECT 1855.800 210.790 1855.940 220.000 ;
        RECT 1855.740 210.470 1856.000 210.790 ;
        RECT 1988.220 210.470 1988.480 210.790 ;
        RECT 1988.280 3.050 1988.420 210.470 ;
        RECT 1988.220 2.730 1988.480 3.050 ;
        RECT 1989.140 2.730 1989.400 3.050 ;
        RECT 1989.200 2.400 1989.340 2.730 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1870.430 212.740 1870.750 212.800 ;
        RECT 2001.990 212.740 2002.310 212.800 ;
        RECT 1870.430 212.600 2002.310 212.740 ;
        RECT 1870.430 212.540 1870.750 212.600 ;
        RECT 2001.990 212.540 2002.310 212.600 ;
        RECT 2001.990 2.960 2002.310 3.020 ;
        RECT 2006.590 2.960 2006.910 3.020 ;
        RECT 2001.990 2.820 2006.910 2.960 ;
        RECT 2001.990 2.760 2002.310 2.820 ;
        RECT 2006.590 2.760 2006.910 2.820 ;
      LAYER via ;
        RECT 1870.460 212.540 1870.720 212.800 ;
        RECT 2002.020 212.540 2002.280 212.800 ;
        RECT 2002.020 2.760 2002.280 3.020 ;
        RECT 2006.620 2.760 2006.880 3.020 ;
      LAYER met2 ;
        RECT 1870.500 220.000 1870.780 224.000 ;
        RECT 1870.520 212.830 1870.660 220.000 ;
        RECT 1870.460 212.510 1870.720 212.830 ;
        RECT 2002.020 212.510 2002.280 212.830 ;
        RECT 2002.080 3.050 2002.220 212.510 ;
        RECT 2002.020 2.730 2002.280 3.050 ;
        RECT 2006.620 2.730 2006.880 3.050 ;
        RECT 2006.680 2.400 2006.820 2.730 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2022.305 48.365 2022.475 96.475 ;
      LAYER mcon ;
        RECT 2022.305 96.305 2022.475 96.475 ;
      LAYER met1 ;
        RECT 1884.690 210.360 1885.010 210.420 ;
        RECT 2022.690 210.360 2023.010 210.420 ;
        RECT 1884.690 210.220 2023.010 210.360 ;
        RECT 1884.690 210.160 1885.010 210.220 ;
        RECT 2022.690 210.160 2023.010 210.220 ;
        RECT 2022.245 96.460 2022.535 96.505 ;
        RECT 2023.610 96.460 2023.930 96.520 ;
        RECT 2022.245 96.320 2023.930 96.460 ;
        RECT 2022.245 96.275 2022.535 96.320 ;
        RECT 2023.610 96.260 2023.930 96.320 ;
        RECT 2022.230 48.520 2022.550 48.580 ;
        RECT 2022.035 48.380 2022.550 48.520 ;
        RECT 2022.230 48.320 2022.550 48.380 ;
        RECT 2022.230 3.300 2022.550 3.360 ;
        RECT 2022.230 3.160 2024.760 3.300 ;
        RECT 2022.230 3.100 2022.550 3.160 ;
        RECT 2024.620 3.020 2024.760 3.160 ;
        RECT 2024.530 2.760 2024.850 3.020 ;
      LAYER via ;
        RECT 1884.720 210.160 1884.980 210.420 ;
        RECT 2022.720 210.160 2022.980 210.420 ;
        RECT 2023.640 96.260 2023.900 96.520 ;
        RECT 2022.260 48.320 2022.520 48.580 ;
        RECT 2022.260 3.100 2022.520 3.360 ;
        RECT 2024.560 2.760 2024.820 3.020 ;
      LAYER met2 ;
        RECT 1884.760 220.000 1885.040 224.000 ;
        RECT 1884.780 210.450 1884.920 220.000 ;
        RECT 1884.720 210.130 1884.980 210.450 ;
        RECT 2022.720 210.130 2022.980 210.450 ;
        RECT 2022.780 158.850 2022.920 210.130 ;
        RECT 2022.780 158.710 2023.380 158.850 ;
        RECT 2023.240 122.130 2023.380 158.710 ;
        RECT 2023.240 121.990 2023.840 122.130 ;
        RECT 2023.700 96.550 2023.840 121.990 ;
        RECT 2023.640 96.230 2023.900 96.550 ;
        RECT 2022.260 48.290 2022.520 48.610 ;
        RECT 2022.320 3.390 2022.460 48.290 ;
        RECT 2022.260 3.070 2022.520 3.390 ;
        RECT 2024.560 2.730 2024.820 3.050 ;
        RECT 2024.620 2.400 2024.760 2.730 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1899.410 212.060 1899.730 212.120 ;
        RECT 2042.930 212.060 2043.250 212.120 ;
        RECT 1899.410 211.920 2043.250 212.060 ;
        RECT 1899.410 211.860 1899.730 211.920 ;
        RECT 2042.930 211.860 2043.250 211.920 ;
      LAYER via ;
        RECT 1899.440 211.860 1899.700 212.120 ;
        RECT 2042.960 211.860 2043.220 212.120 ;
      LAYER met2 ;
        RECT 1899.480 220.000 1899.760 224.000 ;
        RECT 1899.500 212.150 1899.640 220.000 ;
        RECT 1899.440 211.830 1899.700 212.150 ;
        RECT 2042.960 211.830 2043.220 212.150 ;
        RECT 2043.020 3.130 2043.160 211.830 ;
        RECT 2042.560 2.990 2043.160 3.130 ;
        RECT 2042.560 2.400 2042.700 2.990 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 758.610 211.720 758.930 211.780 ;
        RECT 841.870 211.720 842.190 211.780 ;
        RECT 758.610 211.580 842.190 211.720 ;
        RECT 758.610 211.520 758.930 211.580 ;
        RECT 841.870 211.520 842.190 211.580 ;
      LAYER via ;
        RECT 758.640 211.520 758.900 211.780 ;
        RECT 841.900 211.520 842.160 211.780 ;
      LAYER met2 ;
        RECT 841.940 220.000 842.220 224.000 ;
        RECT 841.960 211.810 842.100 220.000 ;
        RECT 758.640 211.490 758.900 211.810 ;
        RECT 841.900 211.490 842.160 211.810 ;
        RECT 758.700 17.410 758.840 211.490 ;
        RECT 757.780 17.270 758.840 17.410 ;
        RECT 757.780 2.400 757.920 17.270 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1914.130 213.760 1914.450 213.820 ;
        RECT 2057.190 213.760 2057.510 213.820 ;
        RECT 1914.130 213.620 2057.510 213.760 ;
        RECT 1914.130 213.560 1914.450 213.620 ;
        RECT 2057.190 213.560 2057.510 213.620 ;
        RECT 2057.190 2.960 2057.510 3.020 ;
        RECT 2060.410 2.960 2060.730 3.020 ;
        RECT 2057.190 2.820 2060.730 2.960 ;
        RECT 2057.190 2.760 2057.510 2.820 ;
        RECT 2060.410 2.760 2060.730 2.820 ;
      LAYER via ;
        RECT 1914.160 213.560 1914.420 213.820 ;
        RECT 2057.220 213.560 2057.480 213.820 ;
        RECT 2057.220 2.760 2057.480 3.020 ;
        RECT 2060.440 2.760 2060.700 3.020 ;
      LAYER met2 ;
        RECT 1914.200 220.000 1914.480 224.000 ;
        RECT 1914.220 213.850 1914.360 220.000 ;
        RECT 1914.160 213.530 1914.420 213.850 ;
        RECT 2057.220 213.530 2057.480 213.850 ;
        RECT 2057.280 3.050 2057.420 213.530 ;
        RECT 2057.220 2.730 2057.480 3.050 ;
        RECT 2060.440 2.730 2060.700 3.050 ;
        RECT 2060.500 2.400 2060.640 2.730 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1928.850 211.720 1929.170 211.780 ;
        RECT 2077.430 211.720 2077.750 211.780 ;
        RECT 1928.850 211.580 2077.750 211.720 ;
        RECT 1928.850 211.520 1929.170 211.580 ;
        RECT 2077.430 211.520 2077.750 211.580 ;
        RECT 2077.430 2.960 2077.750 3.020 ;
        RECT 2078.350 2.960 2078.670 3.020 ;
        RECT 2077.430 2.820 2078.670 2.960 ;
        RECT 2077.430 2.760 2077.750 2.820 ;
        RECT 2078.350 2.760 2078.670 2.820 ;
      LAYER via ;
        RECT 1928.880 211.520 1929.140 211.780 ;
        RECT 2077.460 211.520 2077.720 211.780 ;
        RECT 2077.460 2.760 2077.720 3.020 ;
        RECT 2078.380 2.760 2078.640 3.020 ;
      LAYER met2 ;
        RECT 1928.920 220.000 1929.200 224.000 ;
        RECT 1928.940 211.810 1929.080 220.000 ;
        RECT 1928.880 211.490 1929.140 211.810 ;
        RECT 2077.460 211.490 2077.720 211.810 ;
        RECT 2077.520 3.050 2077.660 211.490 ;
        RECT 2077.460 2.730 2077.720 3.050 ;
        RECT 2078.380 2.730 2078.640 3.050 ;
        RECT 2078.440 2.400 2078.580 2.730 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1943.570 211.380 1943.890 211.440 ;
        RECT 2091.230 211.380 2091.550 211.440 ;
        RECT 1943.570 211.240 2091.550 211.380 ;
        RECT 1943.570 211.180 1943.890 211.240 ;
        RECT 2091.230 211.180 2091.550 211.240 ;
        RECT 2091.230 2.960 2091.550 3.020 ;
        RECT 2095.830 2.960 2096.150 3.020 ;
        RECT 2091.230 2.820 2096.150 2.960 ;
        RECT 2091.230 2.760 2091.550 2.820 ;
        RECT 2095.830 2.760 2096.150 2.820 ;
      LAYER via ;
        RECT 1943.600 211.180 1943.860 211.440 ;
        RECT 2091.260 211.180 2091.520 211.440 ;
        RECT 2091.260 2.760 2091.520 3.020 ;
        RECT 2095.860 2.760 2096.120 3.020 ;
      LAYER met2 ;
        RECT 1943.640 220.000 1943.920 224.000 ;
        RECT 1943.660 211.470 1943.800 220.000 ;
        RECT 1943.600 211.150 1943.860 211.470 ;
        RECT 2091.260 211.150 2091.520 211.470 ;
        RECT 2091.320 3.050 2091.460 211.150 ;
        RECT 2091.260 2.730 2091.520 3.050 ;
        RECT 2095.860 2.730 2096.120 3.050 ;
        RECT 2095.920 2.400 2096.060 2.730 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1958.750 24.040 1959.070 24.100 ;
        RECT 2113.770 24.040 2114.090 24.100 ;
        RECT 1958.750 23.900 2114.090 24.040 ;
        RECT 1958.750 23.840 1959.070 23.900 ;
        RECT 2113.770 23.840 2114.090 23.900 ;
      LAYER via ;
        RECT 1958.780 23.840 1959.040 24.100 ;
        RECT 2113.800 23.840 2114.060 24.100 ;
      LAYER met2 ;
        RECT 1958.360 220.730 1958.640 224.000 ;
        RECT 1958.360 220.590 1958.980 220.730 ;
        RECT 1958.360 220.000 1958.640 220.590 ;
        RECT 1958.840 24.130 1958.980 220.590 ;
        RECT 1958.780 23.810 1959.040 24.130 ;
        RECT 2113.800 23.810 2114.060 24.130 ;
        RECT 2113.860 2.400 2114.000 23.810 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1973.010 210.020 1973.330 210.080 ;
        RECT 2126.190 210.020 2126.510 210.080 ;
        RECT 1973.010 209.880 2126.510 210.020 ;
        RECT 1973.010 209.820 1973.330 209.880 ;
        RECT 2126.190 209.820 2126.510 209.880 ;
        RECT 2126.190 2.960 2126.510 3.020 ;
        RECT 2131.710 2.960 2132.030 3.020 ;
        RECT 2126.190 2.820 2132.030 2.960 ;
        RECT 2126.190 2.760 2126.510 2.820 ;
        RECT 2131.710 2.760 2132.030 2.820 ;
      LAYER via ;
        RECT 1973.040 209.820 1973.300 210.080 ;
        RECT 2126.220 209.820 2126.480 210.080 ;
        RECT 2126.220 2.760 2126.480 3.020 ;
        RECT 2131.740 2.760 2132.000 3.020 ;
      LAYER met2 ;
        RECT 1973.080 220.000 1973.360 224.000 ;
        RECT 1973.100 210.110 1973.240 220.000 ;
        RECT 1973.040 209.790 1973.300 210.110 ;
        RECT 2126.220 209.790 2126.480 210.110 ;
        RECT 2126.280 3.050 2126.420 209.790 ;
        RECT 2126.220 2.730 2126.480 3.050 ;
        RECT 2131.740 2.730 2132.000 3.050 ;
        RECT 2131.800 2.400 2131.940 2.730 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1987.730 207.300 1988.050 207.360 ;
        RECT 1993.250 207.300 1993.570 207.360 ;
        RECT 1987.730 207.160 1993.570 207.300 ;
        RECT 1987.730 207.100 1988.050 207.160 ;
        RECT 1993.250 207.100 1993.570 207.160 ;
        RECT 1993.250 26.080 1993.570 26.140 ;
        RECT 2149.650 26.080 2149.970 26.140 ;
        RECT 1993.250 25.940 2149.970 26.080 ;
        RECT 1993.250 25.880 1993.570 25.940 ;
        RECT 2149.650 25.880 2149.970 25.940 ;
      LAYER via ;
        RECT 1987.760 207.100 1988.020 207.360 ;
        RECT 1993.280 207.100 1993.540 207.360 ;
        RECT 1993.280 25.880 1993.540 26.140 ;
        RECT 2149.680 25.880 2149.940 26.140 ;
      LAYER met2 ;
        RECT 1987.800 220.000 1988.080 224.000 ;
        RECT 1987.820 207.390 1987.960 220.000 ;
        RECT 1987.760 207.070 1988.020 207.390 ;
        RECT 1993.280 207.070 1993.540 207.390 ;
        RECT 1993.340 26.170 1993.480 207.070 ;
        RECT 1993.280 25.850 1993.540 26.170 ;
        RECT 2149.680 25.850 2149.940 26.170 ;
        RECT 2149.740 2.400 2149.880 25.850 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2167.205 138.125 2167.375 186.235 ;
        RECT 2167.205 41.905 2167.375 89.675 ;
        RECT 2167.665 2.805 2167.835 41.395 ;
      LAYER mcon ;
        RECT 2167.205 186.065 2167.375 186.235 ;
        RECT 2167.205 89.505 2167.375 89.675 ;
        RECT 2167.665 41.225 2167.835 41.395 ;
      LAYER met1 ;
        RECT 2002.450 210.700 2002.770 210.760 ;
        RECT 2167.130 210.700 2167.450 210.760 ;
        RECT 2002.450 210.560 2167.450 210.700 ;
        RECT 2002.450 210.500 2002.770 210.560 ;
        RECT 2167.130 210.500 2167.450 210.560 ;
        RECT 2167.130 186.220 2167.450 186.280 ;
        RECT 2166.935 186.080 2167.450 186.220 ;
        RECT 2167.130 186.020 2167.450 186.080 ;
        RECT 2167.130 138.280 2167.450 138.340 ;
        RECT 2166.935 138.140 2167.450 138.280 ;
        RECT 2167.130 138.080 2167.450 138.140 ;
        RECT 2167.130 89.660 2167.450 89.720 ;
        RECT 2166.935 89.520 2167.450 89.660 ;
        RECT 2167.130 89.460 2167.450 89.520 ;
        RECT 2167.130 42.060 2167.450 42.120 ;
        RECT 2166.935 41.920 2167.450 42.060 ;
        RECT 2167.130 41.860 2167.450 41.920 ;
        RECT 2167.130 41.380 2167.450 41.440 ;
        RECT 2167.605 41.380 2167.895 41.425 ;
        RECT 2167.130 41.240 2167.895 41.380 ;
        RECT 2167.130 41.180 2167.450 41.240 ;
        RECT 2167.605 41.195 2167.895 41.240 ;
        RECT 2167.590 2.960 2167.910 3.020 ;
        RECT 2167.395 2.820 2167.910 2.960 ;
        RECT 2167.590 2.760 2167.910 2.820 ;
      LAYER via ;
        RECT 2002.480 210.500 2002.740 210.760 ;
        RECT 2167.160 210.500 2167.420 210.760 ;
        RECT 2167.160 186.020 2167.420 186.280 ;
        RECT 2167.160 138.080 2167.420 138.340 ;
        RECT 2167.160 89.460 2167.420 89.720 ;
        RECT 2167.160 41.860 2167.420 42.120 ;
        RECT 2167.160 41.180 2167.420 41.440 ;
        RECT 2167.620 2.760 2167.880 3.020 ;
      LAYER met2 ;
        RECT 2002.520 220.000 2002.800 224.000 ;
        RECT 2002.540 210.790 2002.680 220.000 ;
        RECT 2002.480 210.470 2002.740 210.790 ;
        RECT 2167.160 210.470 2167.420 210.790 ;
        RECT 2167.220 186.310 2167.360 210.470 ;
        RECT 2167.160 185.990 2167.420 186.310 ;
        RECT 2167.160 138.050 2167.420 138.370 ;
        RECT 2167.220 89.750 2167.360 138.050 ;
        RECT 2167.160 89.430 2167.420 89.750 ;
        RECT 2167.160 41.830 2167.420 42.150 ;
        RECT 2167.220 41.470 2167.360 41.830 ;
        RECT 2167.160 41.150 2167.420 41.470 ;
        RECT 2167.620 2.730 2167.880 3.050 ;
        RECT 2167.680 2.400 2167.820 2.730 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2017.170 213.420 2017.490 213.480 ;
        RECT 2021.310 213.420 2021.630 213.480 ;
        RECT 2017.170 213.280 2021.630 213.420 ;
        RECT 2017.170 213.220 2017.490 213.280 ;
        RECT 2021.310 213.220 2021.630 213.280 ;
        RECT 2021.310 25.740 2021.630 25.800 ;
        RECT 2185.070 25.740 2185.390 25.800 ;
        RECT 2021.310 25.600 2185.390 25.740 ;
        RECT 2021.310 25.540 2021.630 25.600 ;
        RECT 2185.070 25.540 2185.390 25.600 ;
      LAYER via ;
        RECT 2017.200 213.220 2017.460 213.480 ;
        RECT 2021.340 213.220 2021.600 213.480 ;
        RECT 2021.340 25.540 2021.600 25.800 ;
        RECT 2185.100 25.540 2185.360 25.800 ;
      LAYER met2 ;
        RECT 2017.240 220.000 2017.520 224.000 ;
        RECT 2017.260 213.510 2017.400 220.000 ;
        RECT 2017.200 213.190 2017.460 213.510 ;
        RECT 2021.340 213.190 2021.600 213.510 ;
        RECT 2021.400 25.830 2021.540 213.190 ;
        RECT 2021.340 25.510 2021.600 25.830 ;
        RECT 2185.100 25.510 2185.360 25.830 ;
        RECT 2185.160 2.400 2185.300 25.510 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2035.110 25.400 2035.430 25.460 ;
        RECT 2203.010 25.400 2203.330 25.460 ;
        RECT 2035.110 25.260 2203.330 25.400 ;
        RECT 2035.110 25.200 2035.430 25.260 ;
        RECT 2203.010 25.200 2203.330 25.260 ;
      LAYER via ;
        RECT 2035.140 25.200 2035.400 25.460 ;
        RECT 2203.040 25.200 2203.300 25.460 ;
      LAYER met2 ;
        RECT 2031.960 220.730 2032.240 224.000 ;
        RECT 2031.960 220.590 2035.340 220.730 ;
        RECT 2031.960 220.000 2032.240 220.590 ;
        RECT 2035.200 25.490 2035.340 220.590 ;
        RECT 2035.140 25.170 2035.400 25.490 ;
        RECT 2203.040 25.170 2203.300 25.490 ;
        RECT 2203.100 2.400 2203.240 25.170 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2048.910 25.060 2049.230 25.120 ;
        RECT 2220.950 25.060 2221.270 25.120 ;
        RECT 2048.910 24.920 2221.270 25.060 ;
        RECT 2048.910 24.860 2049.230 24.920 ;
        RECT 2220.950 24.860 2221.270 24.920 ;
      LAYER via ;
        RECT 2048.940 24.860 2049.200 25.120 ;
        RECT 2220.980 24.860 2221.240 25.120 ;
      LAYER met2 ;
        RECT 2046.680 220.730 2046.960 224.000 ;
        RECT 2046.680 220.590 2049.140 220.730 ;
        RECT 2046.680 220.000 2046.960 220.590 ;
        RECT 2049.000 25.150 2049.140 220.590 ;
        RECT 2048.940 24.830 2049.200 25.150 ;
        RECT 2220.980 24.830 2221.240 25.150 ;
        RECT 2221.040 2.400 2221.180 24.830 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 779.310 213.080 779.630 213.140 ;
        RECT 856.590 213.080 856.910 213.140 ;
        RECT 779.310 212.940 856.910 213.080 ;
        RECT 779.310 212.880 779.630 212.940 ;
        RECT 856.590 212.880 856.910 212.940 ;
        RECT 775.630 17.580 775.950 17.640 ;
        RECT 779.310 17.580 779.630 17.640 ;
        RECT 775.630 17.440 779.630 17.580 ;
        RECT 775.630 17.380 775.950 17.440 ;
        RECT 779.310 17.380 779.630 17.440 ;
      LAYER via ;
        RECT 779.340 212.880 779.600 213.140 ;
        RECT 856.620 212.880 856.880 213.140 ;
        RECT 775.660 17.380 775.920 17.640 ;
        RECT 779.340 17.380 779.600 17.640 ;
      LAYER met2 ;
        RECT 856.660 220.000 856.940 224.000 ;
        RECT 856.680 213.170 856.820 220.000 ;
        RECT 779.340 212.850 779.600 213.170 ;
        RECT 856.620 212.850 856.880 213.170 ;
        RECT 779.400 17.670 779.540 212.850 ;
        RECT 775.660 17.350 775.920 17.670 ;
        RECT 779.340 17.350 779.600 17.670 ;
        RECT 775.720 2.400 775.860 17.350 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2062.710 24.380 2063.030 24.440 ;
        RECT 2238.890 24.380 2239.210 24.440 ;
        RECT 2062.710 24.240 2239.210 24.380 ;
        RECT 2062.710 24.180 2063.030 24.240 ;
        RECT 2238.890 24.180 2239.210 24.240 ;
      LAYER via ;
        RECT 2062.740 24.180 2063.000 24.440 ;
        RECT 2238.920 24.180 2239.180 24.440 ;
      LAYER met2 ;
        RECT 2061.400 220.730 2061.680 224.000 ;
        RECT 2061.400 220.590 2062.940 220.730 ;
        RECT 2061.400 220.000 2061.680 220.590 ;
        RECT 2062.800 24.470 2062.940 220.590 ;
        RECT 2062.740 24.150 2063.000 24.470 ;
        RECT 2238.920 24.150 2239.180 24.470 ;
        RECT 2238.980 2.400 2239.120 24.150 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2076.510 24.720 2076.830 24.780 ;
        RECT 2256.370 24.720 2256.690 24.780 ;
        RECT 2076.510 24.580 2256.690 24.720 ;
        RECT 2076.510 24.520 2076.830 24.580 ;
        RECT 2256.370 24.520 2256.690 24.580 ;
      LAYER via ;
        RECT 2076.540 24.520 2076.800 24.780 ;
        RECT 2256.400 24.520 2256.660 24.780 ;
      LAYER met2 ;
        RECT 2076.120 220.730 2076.400 224.000 ;
        RECT 2076.120 220.590 2076.740 220.730 ;
        RECT 2076.120 220.000 2076.400 220.590 ;
        RECT 2076.600 24.810 2076.740 220.590 ;
        RECT 2076.540 24.490 2076.800 24.810 ;
        RECT 2256.400 24.490 2256.660 24.810 ;
        RECT 2256.460 2.400 2256.600 24.490 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2090.770 212.060 2091.090 212.120 ;
        RECT 2270.630 212.060 2270.950 212.120 ;
        RECT 2090.770 211.920 2270.950 212.060 ;
        RECT 2090.770 211.860 2091.090 211.920 ;
        RECT 2270.630 211.860 2270.950 211.920 ;
        RECT 2270.630 2.960 2270.950 3.020 ;
        RECT 2274.310 2.960 2274.630 3.020 ;
        RECT 2270.630 2.820 2274.630 2.960 ;
        RECT 2270.630 2.760 2270.950 2.820 ;
        RECT 2274.310 2.760 2274.630 2.820 ;
      LAYER via ;
        RECT 2090.800 211.860 2091.060 212.120 ;
        RECT 2270.660 211.860 2270.920 212.120 ;
        RECT 2270.660 2.760 2270.920 3.020 ;
        RECT 2274.340 2.760 2274.600 3.020 ;
      LAYER met2 ;
        RECT 2090.840 220.000 2091.120 224.000 ;
        RECT 2090.860 212.150 2091.000 220.000 ;
        RECT 2090.800 211.830 2091.060 212.150 ;
        RECT 2270.660 211.830 2270.920 212.150 ;
        RECT 2270.720 3.050 2270.860 211.830 ;
        RECT 2270.660 2.730 2270.920 3.050 ;
        RECT 2274.340 2.730 2274.600 3.050 ;
        RECT 2274.400 2.400 2274.540 2.730 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2186.985 26.605 2187.615 26.775 ;
        RECT 2215.045 25.925 2215.215 26.775 ;
        RECT 2227.925 25.925 2228.095 26.775 ;
        RECT 2270.245 24.565 2270.415 26.775 ;
      LAYER mcon ;
        RECT 2187.445 26.605 2187.615 26.775 ;
        RECT 2215.045 26.605 2215.215 26.775 ;
        RECT 2227.925 26.605 2228.095 26.775 ;
        RECT 2270.245 26.605 2270.415 26.775 ;
      LAYER met1 ;
        RECT 2105.490 207.300 2105.810 207.360 ;
        RECT 2110.550 207.300 2110.870 207.360 ;
        RECT 2105.490 207.160 2110.870 207.300 ;
        RECT 2105.490 207.100 2105.810 207.160 ;
        RECT 2110.550 207.100 2110.870 207.160 ;
        RECT 2262.900 26.960 2270.400 27.100 ;
        RECT 2110.550 26.760 2110.870 26.820 ;
        RECT 2186.925 26.760 2187.215 26.805 ;
        RECT 2110.550 26.620 2187.215 26.760 ;
        RECT 2110.550 26.560 2110.870 26.620 ;
        RECT 2186.925 26.575 2187.215 26.620 ;
        RECT 2187.385 26.760 2187.675 26.805 ;
        RECT 2214.985 26.760 2215.275 26.805 ;
        RECT 2187.385 26.620 2215.275 26.760 ;
        RECT 2187.385 26.575 2187.675 26.620 ;
        RECT 2214.985 26.575 2215.275 26.620 ;
        RECT 2227.865 26.760 2228.155 26.805 ;
        RECT 2262.900 26.760 2263.040 26.960 ;
        RECT 2270.260 26.805 2270.400 26.960 ;
        RECT 2227.865 26.620 2263.040 26.760 ;
        RECT 2227.865 26.575 2228.155 26.620 ;
        RECT 2270.185 26.575 2270.475 26.805 ;
        RECT 2214.985 26.080 2215.275 26.125 ;
        RECT 2227.865 26.080 2228.155 26.125 ;
        RECT 2214.985 25.940 2228.155 26.080 ;
        RECT 2214.985 25.895 2215.275 25.940 ;
        RECT 2227.865 25.895 2228.155 25.940 ;
        RECT 2270.185 24.720 2270.475 24.765 ;
        RECT 2292.250 24.720 2292.570 24.780 ;
        RECT 2270.185 24.580 2292.570 24.720 ;
        RECT 2270.185 24.535 2270.475 24.580 ;
        RECT 2292.250 24.520 2292.570 24.580 ;
      LAYER via ;
        RECT 2105.520 207.100 2105.780 207.360 ;
        RECT 2110.580 207.100 2110.840 207.360 ;
        RECT 2110.580 26.560 2110.840 26.820 ;
        RECT 2292.280 24.520 2292.540 24.780 ;
      LAYER met2 ;
        RECT 2105.560 220.000 2105.840 224.000 ;
        RECT 2105.580 207.390 2105.720 220.000 ;
        RECT 2105.520 207.070 2105.780 207.390 ;
        RECT 2110.580 207.070 2110.840 207.390 ;
        RECT 2110.640 26.850 2110.780 207.070 ;
        RECT 2110.580 26.530 2110.840 26.850 ;
        RECT 2292.280 24.490 2292.540 24.810 ;
        RECT 2292.340 2.400 2292.480 24.490 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2120.210 207.300 2120.530 207.360 ;
        RECT 2124.350 207.300 2124.670 207.360 ;
        RECT 2120.210 207.160 2124.670 207.300 ;
        RECT 2120.210 207.100 2120.530 207.160 ;
        RECT 2124.350 207.100 2124.670 207.160 ;
        RECT 2124.350 24.040 2124.670 24.100 ;
        RECT 2310.190 24.040 2310.510 24.100 ;
        RECT 2124.350 23.900 2310.510 24.040 ;
        RECT 2124.350 23.840 2124.670 23.900 ;
        RECT 2310.190 23.840 2310.510 23.900 ;
      LAYER via ;
        RECT 2120.240 207.100 2120.500 207.360 ;
        RECT 2124.380 207.100 2124.640 207.360 ;
        RECT 2124.380 23.840 2124.640 24.100 ;
        RECT 2310.220 23.840 2310.480 24.100 ;
      LAYER met2 ;
        RECT 2120.280 220.000 2120.560 224.000 ;
        RECT 2120.300 207.390 2120.440 220.000 ;
        RECT 2120.240 207.070 2120.500 207.390 ;
        RECT 2124.380 207.070 2124.640 207.390 ;
        RECT 2124.440 24.130 2124.580 207.070 ;
        RECT 2124.380 23.810 2124.640 24.130 ;
        RECT 2310.220 23.810 2310.480 24.130 ;
        RECT 2310.280 2.400 2310.420 23.810 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2200.325 14.365 2200.495 20.315 ;
      LAYER mcon ;
        RECT 2200.325 20.145 2200.495 20.315 ;
      LAYER met1 ;
        RECT 2134.470 207.300 2134.790 207.360 ;
        RECT 2138.610 207.300 2138.930 207.360 ;
        RECT 2134.470 207.160 2138.930 207.300 ;
        RECT 2134.470 207.100 2134.790 207.160 ;
        RECT 2138.610 207.100 2138.930 207.160 ;
        RECT 2138.610 20.640 2138.930 20.700 ;
        RECT 2138.610 20.500 2163.220 20.640 ;
        RECT 2138.610 20.440 2138.930 20.500 ;
        RECT 2163.080 20.300 2163.220 20.500 ;
        RECT 2200.265 20.300 2200.555 20.345 ;
        RECT 2163.080 20.160 2200.555 20.300 ;
        RECT 2200.265 20.115 2200.555 20.160 ;
        RECT 2200.265 14.520 2200.555 14.565 ;
        RECT 2328.130 14.520 2328.450 14.580 ;
        RECT 2200.265 14.380 2328.450 14.520 ;
        RECT 2200.265 14.335 2200.555 14.380 ;
        RECT 2328.130 14.320 2328.450 14.380 ;
      LAYER via ;
        RECT 2134.500 207.100 2134.760 207.360 ;
        RECT 2138.640 207.100 2138.900 207.360 ;
        RECT 2138.640 20.440 2138.900 20.700 ;
        RECT 2328.160 14.320 2328.420 14.580 ;
      LAYER met2 ;
        RECT 2134.540 220.000 2134.820 224.000 ;
        RECT 2134.560 207.390 2134.700 220.000 ;
        RECT 2134.500 207.070 2134.760 207.390 ;
        RECT 2138.640 207.070 2138.900 207.390 ;
        RECT 2138.700 20.730 2138.840 207.070 ;
        RECT 2138.640 20.410 2138.900 20.730 ;
        RECT 2328.160 14.290 2328.420 14.610 ;
        RECT 2328.220 2.400 2328.360 14.290 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2152.410 15.200 2152.730 15.260 ;
        RECT 2207.150 15.200 2207.470 15.260 ;
        RECT 2152.410 15.060 2207.470 15.200 ;
        RECT 2152.410 15.000 2152.730 15.060 ;
        RECT 2207.150 15.000 2207.470 15.060 ;
        RECT 2235.210 14.860 2235.530 14.920 ;
        RECT 2345.610 14.860 2345.930 14.920 ;
        RECT 2235.210 14.720 2345.930 14.860 ;
        RECT 2235.210 14.660 2235.530 14.720 ;
        RECT 2345.610 14.660 2345.930 14.720 ;
      LAYER via ;
        RECT 2152.440 15.000 2152.700 15.260 ;
        RECT 2207.180 15.000 2207.440 15.260 ;
        RECT 2235.240 14.660 2235.500 14.920 ;
        RECT 2345.640 14.660 2345.900 14.920 ;
      LAYER met2 ;
        RECT 2149.260 220.730 2149.540 224.000 ;
        RECT 2149.260 220.590 2152.640 220.730 ;
        RECT 2149.260 220.000 2149.540 220.590 ;
        RECT 2152.500 15.290 2152.640 220.590 ;
        RECT 2152.440 14.970 2152.700 15.290 ;
        RECT 2207.170 15.115 2207.450 15.485 ;
        RECT 2235.230 15.115 2235.510 15.485 ;
        RECT 2207.180 14.970 2207.440 15.115 ;
        RECT 2235.300 14.950 2235.440 15.115 ;
        RECT 2235.240 14.630 2235.500 14.950 ;
        RECT 2345.640 14.630 2345.900 14.950 ;
        RECT 2345.700 2.400 2345.840 14.630 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
      LAYER via2 ;
        RECT 2207.170 15.160 2207.450 15.440 ;
        RECT 2235.230 15.160 2235.510 15.440 ;
      LAYER met3 ;
        RECT 2207.145 15.450 2207.475 15.465 ;
        RECT 2235.205 15.450 2235.535 15.465 ;
        RECT 2207.145 15.150 2235.535 15.450 ;
        RECT 2207.145 15.135 2207.475 15.150 ;
        RECT 2235.205 15.135 2235.535 15.150 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2192.965 16.065 2193.135 19.975 ;
      LAYER mcon ;
        RECT 2192.965 19.805 2193.135 19.975 ;
      LAYER met1 ;
        RECT 2166.210 19.960 2166.530 20.020 ;
        RECT 2192.905 19.960 2193.195 20.005 ;
        RECT 2166.210 19.820 2193.195 19.960 ;
        RECT 2166.210 19.760 2166.530 19.820 ;
        RECT 2192.905 19.775 2193.195 19.820 ;
        RECT 2192.905 16.220 2193.195 16.265 ;
        RECT 2192.905 16.080 2211.980 16.220 ;
        RECT 2192.905 16.035 2193.195 16.080 ;
        RECT 2211.840 15.880 2211.980 16.080 ;
        RECT 2363.550 15.880 2363.870 15.940 ;
        RECT 2211.840 15.740 2363.870 15.880 ;
        RECT 2363.550 15.680 2363.870 15.740 ;
      LAYER via ;
        RECT 2166.240 19.760 2166.500 20.020 ;
        RECT 2363.580 15.680 2363.840 15.940 ;
      LAYER met2 ;
        RECT 2163.980 220.730 2164.260 224.000 ;
        RECT 2163.980 220.590 2166.440 220.730 ;
        RECT 2163.980 220.000 2164.260 220.590 ;
        RECT 2166.300 20.050 2166.440 220.590 ;
        RECT 2166.240 19.730 2166.500 20.050 ;
        RECT 2363.580 15.650 2363.840 15.970 ;
        RECT 2363.640 2.400 2363.780 15.650 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.010 20.640 2180.330 20.700 ;
        RECT 2381.490 20.640 2381.810 20.700 ;
        RECT 2180.010 20.500 2381.810 20.640 ;
        RECT 2180.010 20.440 2180.330 20.500 ;
        RECT 2381.490 20.440 2381.810 20.500 ;
      LAYER via ;
        RECT 2180.040 20.440 2180.300 20.700 ;
        RECT 2381.520 20.440 2381.780 20.700 ;
      LAYER met2 ;
        RECT 2178.700 220.730 2178.980 224.000 ;
        RECT 2178.700 220.590 2180.240 220.730 ;
        RECT 2178.700 220.000 2178.980 220.590 ;
        RECT 2180.100 20.730 2180.240 220.590 ;
        RECT 2180.040 20.410 2180.300 20.730 ;
        RECT 2381.520 20.410 2381.780 20.730 ;
        RECT 2381.580 2.400 2381.720 20.410 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2193.350 19.960 2193.670 20.020 ;
        RECT 2399.430 19.960 2399.750 20.020 ;
        RECT 2193.350 19.820 2399.750 19.960 ;
        RECT 2193.350 19.760 2193.670 19.820 ;
        RECT 2399.430 19.760 2399.750 19.820 ;
      LAYER via ;
        RECT 2193.380 19.760 2193.640 20.020 ;
        RECT 2399.460 19.760 2399.720 20.020 ;
      LAYER met2 ;
        RECT 2193.420 220.000 2193.700 224.000 ;
        RECT 2193.440 20.050 2193.580 220.000 ;
        RECT 2193.380 19.730 2193.640 20.050 ;
        RECT 2399.460 19.730 2399.720 20.050 ;
        RECT 2399.520 2.400 2399.660 19.730 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 799.550 212.060 799.870 212.120 ;
        RECT 871.310 212.060 871.630 212.120 ;
        RECT 799.550 211.920 871.630 212.060 ;
        RECT 799.550 211.860 799.870 211.920 ;
        RECT 871.310 211.860 871.630 211.920 ;
        RECT 793.570 17.920 793.890 17.980 ;
        RECT 799.550 17.920 799.870 17.980 ;
        RECT 793.570 17.780 799.870 17.920 ;
        RECT 793.570 17.720 793.890 17.780 ;
        RECT 799.550 17.720 799.870 17.780 ;
      LAYER via ;
        RECT 799.580 211.860 799.840 212.120 ;
        RECT 871.340 211.860 871.600 212.120 ;
        RECT 793.600 17.720 793.860 17.980 ;
        RECT 799.580 17.720 799.840 17.980 ;
      LAYER met2 ;
        RECT 871.380 220.000 871.660 224.000 ;
        RECT 871.400 212.150 871.540 220.000 ;
        RECT 799.580 211.830 799.840 212.150 ;
        RECT 871.340 211.830 871.600 212.150 ;
        RECT 799.640 18.010 799.780 211.830 ;
        RECT 793.600 17.690 793.860 18.010 ;
        RECT 799.580 17.690 799.840 18.010 ;
        RECT 793.660 2.400 793.800 17.690 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 641.310 207.980 641.630 208.040 ;
        RECT 743.890 207.980 744.210 208.040 ;
        RECT 641.310 207.840 744.210 207.980 ;
        RECT 641.310 207.780 641.630 207.840 ;
        RECT 743.890 207.780 744.210 207.840 ;
        RECT 639.010 20.640 639.330 20.700 ;
        RECT 641.310 20.640 641.630 20.700 ;
        RECT 639.010 20.500 641.630 20.640 ;
        RECT 639.010 20.440 639.330 20.500 ;
        RECT 641.310 20.440 641.630 20.500 ;
      LAYER via ;
        RECT 641.340 207.780 641.600 208.040 ;
        RECT 743.920 207.780 744.180 208.040 ;
        RECT 639.040 20.440 639.300 20.700 ;
        RECT 641.340 20.440 641.600 20.700 ;
      LAYER met2 ;
        RECT 743.960 220.000 744.240 224.000 ;
        RECT 743.980 208.070 744.120 220.000 ;
        RECT 641.340 207.750 641.600 208.070 ;
        RECT 743.920 207.750 744.180 208.070 ;
        RECT 641.400 20.730 641.540 207.750 ;
        RECT 639.040 20.410 639.300 20.730 ;
        RECT 641.340 20.410 641.600 20.730 ;
        RECT 639.100 2.400 639.240 20.410 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2213.200 220.730 2213.480 224.000 ;
        RECT 2213.200 220.590 2214.740 220.730 ;
        RECT 2213.200 220.000 2213.480 220.590 ;
        RECT 2214.600 16.845 2214.740 220.590 ;
        RECT 2214.530 16.475 2214.810 16.845 ;
        RECT 2422.910 16.475 2423.190 16.845 ;
        RECT 2422.980 2.400 2423.120 16.475 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
      LAYER via2 ;
        RECT 2214.530 16.520 2214.810 16.800 ;
        RECT 2422.910 16.520 2423.190 16.800 ;
      LAYER met3 ;
        RECT 2214.505 16.810 2214.835 16.825 ;
        RECT 2422.885 16.810 2423.215 16.825 ;
        RECT 2214.505 16.510 2423.215 16.810 ;
        RECT 2214.505 16.495 2214.835 16.510 ;
        RECT 2422.885 16.495 2423.215 16.510 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2227.850 210.360 2228.170 210.420 ;
        RECT 2418.750 210.360 2419.070 210.420 ;
        RECT 2227.850 210.220 2419.070 210.360 ;
        RECT 2227.850 210.160 2228.170 210.220 ;
        RECT 2418.750 210.160 2419.070 210.220 ;
        RECT 2418.750 16.220 2419.070 16.280 ;
        RECT 2440.830 16.220 2441.150 16.280 ;
        RECT 2418.750 16.080 2441.150 16.220 ;
        RECT 2418.750 16.020 2419.070 16.080 ;
        RECT 2440.830 16.020 2441.150 16.080 ;
      LAYER via ;
        RECT 2227.880 210.160 2228.140 210.420 ;
        RECT 2418.780 210.160 2419.040 210.420 ;
        RECT 2418.780 16.020 2419.040 16.280 ;
        RECT 2440.860 16.020 2441.120 16.280 ;
      LAYER met2 ;
        RECT 2227.920 220.000 2228.200 224.000 ;
        RECT 2227.940 210.450 2228.080 220.000 ;
        RECT 2227.880 210.130 2228.140 210.450 ;
        RECT 2418.780 210.130 2419.040 210.450 ;
        RECT 2418.840 16.310 2418.980 210.130 ;
        RECT 2418.780 15.990 2419.040 16.310 ;
        RECT 2440.860 15.990 2441.120 16.310 ;
        RECT 2440.920 2.400 2441.060 15.990 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2242.570 207.300 2242.890 207.360 ;
        RECT 2248.550 207.300 2248.870 207.360 ;
        RECT 2242.570 207.160 2248.870 207.300 ;
        RECT 2242.570 207.100 2242.890 207.160 ;
        RECT 2248.550 207.100 2248.870 207.160 ;
        RECT 2458.770 19.280 2459.090 19.340 ;
        RECT 2262.900 19.140 2459.090 19.280 ;
        RECT 2248.550 18.940 2248.870 19.000 ;
        RECT 2262.900 18.940 2263.040 19.140 ;
        RECT 2458.770 19.080 2459.090 19.140 ;
        RECT 2248.550 18.800 2263.040 18.940 ;
        RECT 2248.550 18.740 2248.870 18.800 ;
      LAYER via ;
        RECT 2242.600 207.100 2242.860 207.360 ;
        RECT 2248.580 207.100 2248.840 207.360 ;
        RECT 2248.580 18.740 2248.840 19.000 ;
        RECT 2458.800 19.080 2459.060 19.340 ;
      LAYER met2 ;
        RECT 2242.640 220.000 2242.920 224.000 ;
        RECT 2242.660 207.390 2242.800 220.000 ;
        RECT 2242.600 207.070 2242.860 207.390 ;
        RECT 2248.580 207.070 2248.840 207.390 ;
        RECT 2248.640 19.030 2248.780 207.070 ;
        RECT 2458.800 19.050 2459.060 19.370 ;
        RECT 2248.580 18.710 2248.840 19.030 ;
        RECT 2458.860 2.400 2459.000 19.050 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2286.805 17.085 2286.975 19.635 ;
      LAYER mcon ;
        RECT 2286.805 19.465 2286.975 19.635 ;
      LAYER met1 ;
        RECT 2257.290 207.300 2257.610 207.360 ;
        RECT 2262.810 207.300 2263.130 207.360 ;
        RECT 2257.290 207.160 2263.130 207.300 ;
        RECT 2257.290 207.100 2257.610 207.160 ;
        RECT 2262.810 207.100 2263.130 207.160 ;
        RECT 2286.745 19.620 2287.035 19.665 ;
        RECT 2476.710 19.620 2477.030 19.680 ;
        RECT 2286.745 19.480 2477.030 19.620 ;
        RECT 2286.745 19.435 2287.035 19.480 ;
        RECT 2476.710 19.420 2477.030 19.480 ;
        RECT 2262.810 17.240 2263.130 17.300 ;
        RECT 2286.745 17.240 2287.035 17.285 ;
        RECT 2262.810 17.100 2287.035 17.240 ;
        RECT 2262.810 17.040 2263.130 17.100 ;
        RECT 2286.745 17.055 2287.035 17.100 ;
      LAYER via ;
        RECT 2257.320 207.100 2257.580 207.360 ;
        RECT 2262.840 207.100 2263.100 207.360 ;
        RECT 2476.740 19.420 2477.000 19.680 ;
        RECT 2262.840 17.040 2263.100 17.300 ;
      LAYER met2 ;
        RECT 2257.360 220.000 2257.640 224.000 ;
        RECT 2257.380 207.390 2257.520 220.000 ;
        RECT 2257.320 207.070 2257.580 207.390 ;
        RECT 2262.840 207.070 2263.100 207.390 ;
        RECT 2262.900 17.330 2263.040 207.070 ;
        RECT 2476.740 19.390 2477.000 19.710 ;
        RECT 2262.840 17.010 2263.100 17.330 ;
        RECT 2476.800 2.400 2476.940 19.390 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2272.010 207.300 2272.330 207.360 ;
        RECT 2276.610 207.300 2276.930 207.360 ;
        RECT 2272.010 207.160 2276.930 207.300 ;
        RECT 2272.010 207.100 2272.330 207.160 ;
        RECT 2276.610 207.100 2276.930 207.160 ;
        RECT 2276.610 18.940 2276.930 19.000 ;
        RECT 2494.650 18.940 2494.970 19.000 ;
        RECT 2276.610 18.800 2494.970 18.940 ;
        RECT 2276.610 18.740 2276.930 18.800 ;
        RECT 2494.650 18.740 2494.970 18.800 ;
      LAYER via ;
        RECT 2272.040 207.100 2272.300 207.360 ;
        RECT 2276.640 207.100 2276.900 207.360 ;
        RECT 2276.640 18.740 2276.900 19.000 ;
        RECT 2494.680 18.740 2494.940 19.000 ;
      LAYER met2 ;
        RECT 2272.080 220.000 2272.360 224.000 ;
        RECT 2272.100 207.390 2272.240 220.000 ;
        RECT 2272.040 207.070 2272.300 207.390 ;
        RECT 2276.640 207.070 2276.900 207.390 ;
        RECT 2276.700 19.030 2276.840 207.070 ;
        RECT 2276.640 18.710 2276.900 19.030 ;
        RECT 2494.680 18.710 2494.940 19.030 ;
        RECT 2494.740 2.400 2494.880 18.710 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2511.670 18.260 2511.990 18.320 ;
        RECT 2298.320 18.120 2511.990 18.260 ;
        RECT 2290.410 17.920 2290.730 17.980 ;
        RECT 2298.320 17.920 2298.460 18.120 ;
        RECT 2511.670 18.060 2511.990 18.120 ;
        RECT 2290.410 17.780 2298.460 17.920 ;
        RECT 2290.410 17.720 2290.730 17.780 ;
      LAYER via ;
        RECT 2290.440 17.720 2290.700 17.980 ;
        RECT 2511.700 18.060 2511.960 18.320 ;
      LAYER met2 ;
        RECT 2286.800 220.730 2287.080 224.000 ;
        RECT 2286.800 220.590 2290.640 220.730 ;
        RECT 2286.800 220.000 2287.080 220.590 ;
        RECT 2290.500 18.010 2290.640 220.590 ;
        RECT 2511.700 18.030 2511.960 18.350 ;
        RECT 2290.440 17.690 2290.700 18.010 ;
        RECT 2511.760 17.410 2511.900 18.030 ;
        RECT 2511.760 17.270 2512.360 17.410 ;
        RECT 2512.220 2.400 2512.360 17.270 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2530.070 18.260 2530.390 18.320 ;
        RECT 2512.220 18.120 2530.390 18.260 ;
        RECT 2304.210 17.920 2304.530 17.980 ;
        RECT 2512.220 17.920 2512.360 18.120 ;
        RECT 2530.070 18.060 2530.390 18.120 ;
        RECT 2304.210 17.780 2512.360 17.920 ;
        RECT 2304.210 17.720 2304.530 17.780 ;
      LAYER via ;
        RECT 2304.240 17.720 2304.500 17.980 ;
        RECT 2530.100 18.060 2530.360 18.320 ;
      LAYER met2 ;
        RECT 2301.060 220.730 2301.340 224.000 ;
        RECT 2301.060 220.590 2304.440 220.730 ;
        RECT 2301.060 220.000 2301.340 220.590 ;
        RECT 2304.300 18.010 2304.440 220.590 ;
        RECT 2530.100 18.030 2530.360 18.350 ;
        RECT 2304.240 17.690 2304.500 18.010 ;
        RECT 2530.160 2.400 2530.300 18.030 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2315.710 209.000 2316.030 209.060 ;
        RECT 2507.990 209.000 2508.310 209.060 ;
        RECT 2315.710 208.860 2508.310 209.000 ;
        RECT 2315.710 208.800 2316.030 208.860 ;
        RECT 2507.990 208.800 2508.310 208.860 ;
        RECT 2507.990 19.280 2508.310 19.340 ;
        RECT 2507.990 19.140 2531.220 19.280 ;
        RECT 2507.990 19.080 2508.310 19.140 ;
        RECT 2531.080 18.600 2531.220 19.140 ;
        RECT 2548.010 18.600 2548.330 18.660 ;
        RECT 2531.080 18.460 2548.330 18.600 ;
        RECT 2548.010 18.400 2548.330 18.460 ;
      LAYER via ;
        RECT 2315.740 208.800 2316.000 209.060 ;
        RECT 2508.020 208.800 2508.280 209.060 ;
        RECT 2508.020 19.080 2508.280 19.340 ;
        RECT 2548.040 18.400 2548.300 18.660 ;
      LAYER met2 ;
        RECT 2315.780 220.000 2316.060 224.000 ;
        RECT 2315.800 209.090 2315.940 220.000 ;
        RECT 2315.740 208.770 2316.000 209.090 ;
        RECT 2508.020 208.770 2508.280 209.090 ;
        RECT 2508.080 19.370 2508.220 208.770 ;
        RECT 2508.020 19.050 2508.280 19.370 ;
        RECT 2548.040 18.370 2548.300 18.690 ;
        RECT 2548.100 2.400 2548.240 18.370 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2331.810 17.580 2332.130 17.640 ;
        RECT 2331.810 17.440 2556.060 17.580 ;
        RECT 2331.810 17.380 2332.130 17.440 ;
        RECT 2555.920 17.240 2556.060 17.440 ;
        RECT 2565.950 17.240 2566.270 17.300 ;
        RECT 2555.920 17.100 2566.270 17.240 ;
        RECT 2565.950 17.040 2566.270 17.100 ;
      LAYER via ;
        RECT 2331.840 17.380 2332.100 17.640 ;
        RECT 2565.980 17.040 2566.240 17.300 ;
      LAYER met2 ;
        RECT 2330.500 220.730 2330.780 224.000 ;
        RECT 2330.500 220.590 2332.040 220.730 ;
        RECT 2330.500 220.000 2330.780 220.590 ;
        RECT 2331.900 17.670 2332.040 220.590 ;
        RECT 2331.840 17.350 2332.100 17.670 ;
        RECT 2565.980 17.010 2566.240 17.330 ;
        RECT 2566.040 2.400 2566.180 17.010 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2345.150 211.380 2345.470 211.440 ;
        RECT 2390.690 211.380 2391.010 211.440 ;
        RECT 2345.150 211.240 2391.010 211.380 ;
        RECT 2345.150 211.180 2345.470 211.240 ;
        RECT 2390.690 211.180 2391.010 211.240 ;
        RECT 2390.690 15.200 2391.010 15.260 ;
        RECT 2583.890 15.200 2584.210 15.260 ;
        RECT 2390.690 15.060 2584.210 15.200 ;
        RECT 2390.690 15.000 2391.010 15.060 ;
        RECT 2583.890 15.000 2584.210 15.060 ;
      LAYER via ;
        RECT 2345.180 211.180 2345.440 211.440 ;
        RECT 2390.720 211.180 2390.980 211.440 ;
        RECT 2390.720 15.000 2390.980 15.260 ;
        RECT 2583.920 15.000 2584.180 15.260 ;
      LAYER met2 ;
        RECT 2345.220 220.000 2345.500 224.000 ;
        RECT 2345.240 211.470 2345.380 220.000 ;
        RECT 2345.180 211.150 2345.440 211.470 ;
        RECT 2390.720 211.150 2390.980 211.470 ;
        RECT 2390.780 15.290 2390.920 211.150 ;
        RECT 2390.720 14.970 2390.980 15.290 ;
        RECT 2583.920 14.970 2584.180 15.290 ;
        RECT 2583.980 2.400 2584.120 14.970 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 820.710 210.700 821.030 210.760 ;
        RECT 890.630 210.700 890.950 210.760 ;
        RECT 820.710 210.560 890.950 210.700 ;
        RECT 820.710 210.500 821.030 210.560 ;
        RECT 890.630 210.500 890.950 210.560 ;
        RECT 817.490 17.580 817.810 17.640 ;
        RECT 820.710 17.580 821.030 17.640 ;
        RECT 817.490 17.440 821.030 17.580 ;
        RECT 817.490 17.380 817.810 17.440 ;
        RECT 820.710 17.380 821.030 17.440 ;
      LAYER via ;
        RECT 820.740 210.500 821.000 210.760 ;
        RECT 890.660 210.500 890.920 210.760 ;
        RECT 817.520 17.380 817.780 17.640 ;
        RECT 820.740 17.380 821.000 17.640 ;
      LAYER met2 ;
        RECT 890.700 220.000 890.980 224.000 ;
        RECT 890.720 210.790 890.860 220.000 ;
        RECT 820.740 210.470 821.000 210.790 ;
        RECT 890.660 210.470 890.920 210.790 ;
        RECT 820.800 17.670 820.940 210.470 ;
        RECT 817.520 17.350 817.780 17.670 ;
        RECT 820.740 17.350 821.000 17.670 ;
        RECT 817.580 2.400 817.720 17.350 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2359.870 212.740 2360.190 212.800 ;
        RECT 2418.290 212.740 2418.610 212.800 ;
        RECT 2359.870 212.600 2418.610 212.740 ;
        RECT 2359.870 212.540 2360.190 212.600 ;
        RECT 2418.290 212.540 2418.610 212.600 ;
        RECT 2418.290 14.860 2418.610 14.920 ;
        RECT 2601.370 14.860 2601.690 14.920 ;
        RECT 2418.290 14.720 2601.690 14.860 ;
        RECT 2418.290 14.660 2418.610 14.720 ;
        RECT 2601.370 14.660 2601.690 14.720 ;
      LAYER via ;
        RECT 2359.900 212.540 2360.160 212.800 ;
        RECT 2418.320 212.540 2418.580 212.800 ;
        RECT 2418.320 14.660 2418.580 14.920 ;
        RECT 2601.400 14.660 2601.660 14.920 ;
      LAYER met2 ;
        RECT 2359.940 220.000 2360.220 224.000 ;
        RECT 2359.960 212.830 2360.100 220.000 ;
        RECT 2359.900 212.510 2360.160 212.830 ;
        RECT 2418.320 212.510 2418.580 212.830 ;
        RECT 2418.380 14.950 2418.520 212.510 ;
        RECT 2418.320 14.630 2418.580 14.950 ;
        RECT 2601.400 14.630 2601.660 14.950 ;
        RECT 2601.460 2.400 2601.600 14.630 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2374.590 207.300 2374.910 207.360 ;
        RECT 2380.110 207.300 2380.430 207.360 ;
        RECT 2374.590 207.160 2380.430 207.300 ;
        RECT 2374.590 207.100 2374.910 207.160 ;
        RECT 2380.110 207.100 2380.430 207.160 ;
        RECT 2380.110 16.560 2380.430 16.620 ;
        RECT 2619.310 16.560 2619.630 16.620 ;
        RECT 2380.110 16.420 2619.630 16.560 ;
        RECT 2380.110 16.360 2380.430 16.420 ;
        RECT 2619.310 16.360 2619.630 16.420 ;
      LAYER via ;
        RECT 2374.620 207.100 2374.880 207.360 ;
        RECT 2380.140 207.100 2380.400 207.360 ;
        RECT 2380.140 16.360 2380.400 16.620 ;
        RECT 2619.340 16.360 2619.600 16.620 ;
      LAYER met2 ;
        RECT 2374.660 220.000 2374.940 224.000 ;
        RECT 2374.680 207.390 2374.820 220.000 ;
        RECT 2374.620 207.070 2374.880 207.390 ;
        RECT 2380.140 207.070 2380.400 207.390 ;
        RECT 2380.200 16.650 2380.340 207.070 ;
        RECT 2380.140 16.330 2380.400 16.650 ;
        RECT 2619.340 16.330 2619.600 16.650 ;
        RECT 2619.400 2.400 2619.540 16.330 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2389.310 211.040 2389.630 211.100 ;
        RECT 2635.870 211.040 2636.190 211.100 ;
        RECT 2389.310 210.900 2636.190 211.040 ;
        RECT 2389.310 210.840 2389.630 210.900 ;
        RECT 2635.870 210.840 2636.190 210.900 ;
      LAYER via ;
        RECT 2389.340 210.840 2389.600 211.100 ;
        RECT 2635.900 210.840 2636.160 211.100 ;
      LAYER met2 ;
        RECT 2389.380 220.000 2389.660 224.000 ;
        RECT 2389.400 211.130 2389.540 220.000 ;
        RECT 2389.340 210.810 2389.600 211.130 ;
        RECT 2635.900 210.810 2636.160 211.130 ;
        RECT 2635.960 17.410 2636.100 210.810 ;
        RECT 2635.960 17.270 2637.480 17.410 ;
        RECT 2637.340 2.400 2637.480 17.270 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2404.030 207.300 2404.350 207.360 ;
        RECT 2407.710 207.300 2408.030 207.360 ;
        RECT 2404.030 207.160 2408.030 207.300 ;
        RECT 2404.030 207.100 2404.350 207.160 ;
        RECT 2407.710 207.100 2408.030 207.160 ;
        RECT 2407.710 15.540 2408.030 15.600 ;
        RECT 2655.190 15.540 2655.510 15.600 ;
        RECT 2407.710 15.400 2655.510 15.540 ;
        RECT 2407.710 15.340 2408.030 15.400 ;
        RECT 2655.190 15.340 2655.510 15.400 ;
      LAYER via ;
        RECT 2404.060 207.100 2404.320 207.360 ;
        RECT 2407.740 207.100 2408.000 207.360 ;
        RECT 2407.740 15.340 2408.000 15.600 ;
        RECT 2655.220 15.340 2655.480 15.600 ;
      LAYER met2 ;
        RECT 2404.100 220.000 2404.380 224.000 ;
        RECT 2404.120 207.390 2404.260 220.000 ;
        RECT 2404.060 207.070 2404.320 207.390 ;
        RECT 2407.740 207.070 2408.000 207.390 ;
        RECT 2407.800 15.630 2407.940 207.070 ;
        RECT 2407.740 15.310 2408.000 15.630 ;
        RECT 2655.220 15.310 2655.480 15.630 ;
        RECT 2655.280 2.400 2655.420 15.310 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2418.750 212.060 2419.070 212.120 ;
        RECT 2652.890 212.060 2653.210 212.120 ;
        RECT 2418.750 211.920 2653.210 212.060 ;
        RECT 2418.750 211.860 2419.070 211.920 ;
        RECT 2652.890 211.860 2653.210 211.920 ;
        RECT 2652.890 16.560 2653.210 16.620 ;
        RECT 2672.670 16.560 2672.990 16.620 ;
        RECT 2652.890 16.420 2672.990 16.560 ;
        RECT 2652.890 16.360 2653.210 16.420 ;
        RECT 2672.670 16.360 2672.990 16.420 ;
      LAYER via ;
        RECT 2418.780 211.860 2419.040 212.120 ;
        RECT 2652.920 211.860 2653.180 212.120 ;
        RECT 2652.920 16.360 2653.180 16.620 ;
        RECT 2672.700 16.360 2672.960 16.620 ;
      LAYER met2 ;
        RECT 2418.820 220.000 2419.100 224.000 ;
        RECT 2418.840 212.150 2418.980 220.000 ;
        RECT 2418.780 211.830 2419.040 212.150 ;
        RECT 2652.920 211.830 2653.180 212.150 ;
        RECT 2652.980 16.650 2653.120 211.830 ;
        RECT 2652.920 16.330 2653.180 16.650 ;
        RECT 2672.700 16.330 2672.960 16.650 ;
        RECT 2672.760 2.400 2672.900 16.330 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2433.470 212.740 2433.790 212.800 ;
        RECT 2659.790 212.740 2660.110 212.800 ;
        RECT 2433.470 212.600 2660.110 212.740 ;
        RECT 2433.470 212.540 2433.790 212.600 ;
        RECT 2659.790 212.540 2660.110 212.600 ;
        RECT 2659.790 14.860 2660.110 14.920 ;
        RECT 2690.610 14.860 2690.930 14.920 ;
        RECT 2659.790 14.720 2690.930 14.860 ;
        RECT 2659.790 14.660 2660.110 14.720 ;
        RECT 2690.610 14.660 2690.930 14.720 ;
      LAYER via ;
        RECT 2433.500 212.540 2433.760 212.800 ;
        RECT 2659.820 212.540 2660.080 212.800 ;
        RECT 2659.820 14.660 2660.080 14.920 ;
        RECT 2690.640 14.660 2690.900 14.920 ;
      LAYER met2 ;
        RECT 2433.540 220.000 2433.820 224.000 ;
        RECT 2433.560 212.830 2433.700 220.000 ;
        RECT 2433.500 212.510 2433.760 212.830 ;
        RECT 2659.820 212.510 2660.080 212.830 ;
        RECT 2659.880 14.950 2660.020 212.510 ;
        RECT 2659.820 14.630 2660.080 14.950 ;
        RECT 2690.640 14.630 2690.900 14.950 ;
        RECT 2690.700 2.400 2690.840 14.630 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2697.585 16.065 2697.755 16.915 ;
      LAYER mcon ;
        RECT 2697.585 16.745 2697.755 16.915 ;
      LAYER met1 ;
        RECT 2449.110 16.900 2449.430 16.960 ;
        RECT 2697.525 16.900 2697.815 16.945 ;
        RECT 2449.110 16.760 2697.815 16.900 ;
        RECT 2449.110 16.700 2449.430 16.760 ;
        RECT 2697.525 16.715 2697.815 16.760 ;
        RECT 2697.525 16.220 2697.815 16.265 ;
        RECT 2708.550 16.220 2708.870 16.280 ;
        RECT 2697.525 16.080 2708.870 16.220 ;
        RECT 2697.525 16.035 2697.815 16.080 ;
        RECT 2708.550 16.020 2708.870 16.080 ;
      LAYER via ;
        RECT 2449.140 16.700 2449.400 16.960 ;
        RECT 2708.580 16.020 2708.840 16.280 ;
      LAYER met2 ;
        RECT 2448.260 220.730 2448.540 224.000 ;
        RECT 2448.260 220.590 2449.340 220.730 ;
        RECT 2448.260 220.000 2448.540 220.590 ;
        RECT 2449.200 16.990 2449.340 220.590 ;
        RECT 2449.140 16.670 2449.400 16.990 ;
        RECT 2708.580 15.990 2708.840 16.310 ;
        RECT 2708.640 2.400 2708.780 15.990 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2462.910 20.300 2463.230 20.360 ;
        RECT 2726.490 20.300 2726.810 20.360 ;
        RECT 2462.910 20.160 2726.810 20.300 ;
        RECT 2462.910 20.100 2463.230 20.160 ;
        RECT 2726.490 20.100 2726.810 20.160 ;
      LAYER via ;
        RECT 2462.940 20.100 2463.200 20.360 ;
        RECT 2726.520 20.100 2726.780 20.360 ;
      LAYER met2 ;
        RECT 2462.980 220.000 2463.260 224.000 ;
        RECT 2463.000 20.390 2463.140 220.000 ;
        RECT 2462.940 20.070 2463.200 20.390 ;
        RECT 2726.520 20.070 2726.780 20.390 ;
        RECT 2726.580 2.400 2726.720 20.070 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2477.630 209.340 2477.950 209.400 ;
        RECT 2666.690 209.340 2667.010 209.400 ;
        RECT 2477.630 209.200 2667.010 209.340 ;
        RECT 2477.630 209.140 2477.950 209.200 ;
        RECT 2666.690 209.140 2667.010 209.200 ;
        RECT 2744.430 14.860 2744.750 14.920 ;
        RECT 2715.080 14.720 2744.750 14.860 ;
        RECT 2666.690 14.180 2667.010 14.240 ;
        RECT 2715.080 14.180 2715.220 14.720 ;
        RECT 2744.430 14.660 2744.750 14.720 ;
        RECT 2666.690 14.040 2715.220 14.180 ;
        RECT 2666.690 13.980 2667.010 14.040 ;
      LAYER via ;
        RECT 2477.660 209.140 2477.920 209.400 ;
        RECT 2666.720 209.140 2666.980 209.400 ;
        RECT 2666.720 13.980 2666.980 14.240 ;
        RECT 2744.460 14.660 2744.720 14.920 ;
      LAYER met2 ;
        RECT 2477.700 220.000 2477.980 224.000 ;
        RECT 2477.720 209.430 2477.860 220.000 ;
        RECT 2477.660 209.110 2477.920 209.430 ;
        RECT 2666.720 209.110 2666.980 209.430 ;
        RECT 2666.780 14.270 2666.920 209.110 ;
        RECT 2744.460 14.630 2744.720 14.950 ;
        RECT 2666.720 13.950 2666.980 14.270 ;
        RECT 2744.520 2.400 2744.660 14.630 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2492.350 207.300 2492.670 207.360 ;
        RECT 2497.410 207.300 2497.730 207.360 ;
        RECT 2492.350 207.160 2497.730 207.300 ;
        RECT 2492.350 207.100 2492.670 207.160 ;
        RECT 2497.410 207.100 2497.730 207.160 ;
        RECT 2497.410 20.640 2497.730 20.700 ;
        RECT 2761.910 20.640 2762.230 20.700 ;
        RECT 2497.410 20.500 2762.230 20.640 ;
        RECT 2497.410 20.440 2497.730 20.500 ;
        RECT 2761.910 20.440 2762.230 20.500 ;
      LAYER via ;
        RECT 2492.380 207.100 2492.640 207.360 ;
        RECT 2497.440 207.100 2497.700 207.360 ;
        RECT 2497.440 20.440 2497.700 20.700 ;
        RECT 2761.940 20.440 2762.200 20.700 ;
      LAYER met2 ;
        RECT 2492.420 220.000 2492.700 224.000 ;
        RECT 2492.440 207.390 2492.580 220.000 ;
        RECT 2492.380 207.070 2492.640 207.390 ;
        RECT 2497.440 207.070 2497.700 207.390 ;
        RECT 2497.500 20.730 2497.640 207.070 ;
        RECT 2497.440 20.410 2497.700 20.730 ;
        RECT 2761.940 20.410 2762.200 20.730 ;
        RECT 2762.000 2.400 2762.140 20.410 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 841.410 212.740 841.730 212.800 ;
        RECT 905.350 212.740 905.670 212.800 ;
        RECT 841.410 212.600 905.670 212.740 ;
        RECT 841.410 212.540 841.730 212.600 ;
        RECT 905.350 212.540 905.670 212.600 ;
        RECT 835.430 15.540 835.750 15.600 ;
        RECT 841.410 15.540 841.730 15.600 ;
        RECT 835.430 15.400 841.730 15.540 ;
        RECT 835.430 15.340 835.750 15.400 ;
        RECT 841.410 15.340 841.730 15.400 ;
      LAYER via ;
        RECT 841.440 212.540 841.700 212.800 ;
        RECT 905.380 212.540 905.640 212.800 ;
        RECT 835.460 15.340 835.720 15.600 ;
        RECT 841.440 15.340 841.700 15.600 ;
      LAYER met2 ;
        RECT 905.420 220.000 905.700 224.000 ;
        RECT 905.440 212.830 905.580 220.000 ;
        RECT 841.440 212.510 841.700 212.830 ;
        RECT 905.380 212.510 905.640 212.830 ;
        RECT 841.500 15.630 841.640 212.510 ;
        RECT 835.460 15.310 835.720 15.630 ;
        RECT 841.440 15.310 841.700 15.630 ;
        RECT 835.520 2.400 835.660 15.310 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2714.605 15.045 2715.695 15.215 ;
        RECT 2714.605 14.365 2714.775 15.045 ;
      LAYER mcon ;
        RECT 2715.525 15.045 2715.695 15.215 ;
      LAYER met1 ;
        RECT 2507.070 208.660 2507.390 208.720 ;
        RECT 2673.590 208.660 2673.910 208.720 ;
        RECT 2507.070 208.520 2673.910 208.660 ;
        RECT 2507.070 208.460 2507.390 208.520 ;
        RECT 2673.590 208.460 2673.910 208.520 ;
        RECT 2715.465 15.200 2715.755 15.245 ;
        RECT 2779.850 15.200 2780.170 15.260 ;
        RECT 2715.465 15.060 2780.170 15.200 ;
        RECT 2715.465 15.015 2715.755 15.060 ;
        RECT 2779.850 15.000 2780.170 15.060 ;
        RECT 2673.590 14.520 2673.910 14.580 ;
        RECT 2714.545 14.520 2714.835 14.565 ;
        RECT 2673.590 14.380 2714.835 14.520 ;
        RECT 2673.590 14.320 2673.910 14.380 ;
        RECT 2714.545 14.335 2714.835 14.380 ;
      LAYER via ;
        RECT 2507.100 208.460 2507.360 208.720 ;
        RECT 2673.620 208.460 2673.880 208.720 ;
        RECT 2779.880 15.000 2780.140 15.260 ;
        RECT 2673.620 14.320 2673.880 14.580 ;
      LAYER met2 ;
        RECT 2507.140 220.000 2507.420 224.000 ;
        RECT 2507.160 208.750 2507.300 220.000 ;
        RECT 2507.100 208.430 2507.360 208.750 ;
        RECT 2673.620 208.430 2673.880 208.750 ;
        RECT 2673.680 14.610 2673.820 208.430 ;
        RECT 2779.880 14.970 2780.140 15.290 ;
        RECT 2673.620 14.290 2673.880 14.610 ;
        RECT 2779.940 2.400 2780.080 14.970 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2570.165 18.105 2570.335 19.635 ;
      LAYER mcon ;
        RECT 2570.165 19.465 2570.335 19.635 ;
      LAYER met1 ;
        RECT 2570.105 19.620 2570.395 19.665 ;
        RECT 2797.790 19.620 2798.110 19.680 ;
        RECT 2570.105 19.480 2798.110 19.620 ;
        RECT 2570.105 19.435 2570.395 19.480 ;
        RECT 2797.790 19.420 2798.110 19.480 ;
        RECT 2525.010 18.600 2525.330 18.660 ;
        RECT 2525.010 18.460 2530.760 18.600 ;
        RECT 2525.010 18.400 2525.330 18.460 ;
        RECT 2530.620 18.260 2530.760 18.460 ;
        RECT 2570.105 18.260 2570.395 18.305 ;
        RECT 2530.620 18.120 2570.395 18.260 ;
        RECT 2570.105 18.075 2570.395 18.120 ;
      LAYER via ;
        RECT 2797.820 19.420 2798.080 19.680 ;
        RECT 2525.040 18.400 2525.300 18.660 ;
      LAYER met2 ;
        RECT 2521.860 220.730 2522.140 224.000 ;
        RECT 2521.860 220.590 2525.240 220.730 ;
        RECT 2521.860 220.000 2522.140 220.590 ;
        RECT 2525.100 18.690 2525.240 220.590 ;
        RECT 2797.820 19.390 2798.080 19.710 ;
        RECT 2525.040 18.370 2525.300 18.690 ;
        RECT 2797.880 2.400 2798.020 19.390 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2536.510 209.680 2536.830 209.740 ;
        RECT 2687.390 209.680 2687.710 209.740 ;
        RECT 2536.510 209.540 2687.710 209.680 ;
        RECT 2536.510 209.480 2536.830 209.540 ;
        RECT 2687.390 209.480 2687.710 209.540 ;
        RECT 2815.730 15.540 2816.050 15.600 ;
        RECT 2715.080 15.400 2816.050 15.540 ;
        RECT 2687.390 15.200 2687.710 15.260 ;
        RECT 2715.080 15.200 2715.220 15.400 ;
        RECT 2815.730 15.340 2816.050 15.400 ;
        RECT 2687.390 15.060 2715.220 15.200 ;
        RECT 2687.390 15.000 2687.710 15.060 ;
      LAYER via ;
        RECT 2536.540 209.480 2536.800 209.740 ;
        RECT 2687.420 209.480 2687.680 209.740 ;
        RECT 2687.420 15.000 2687.680 15.260 ;
        RECT 2815.760 15.340 2816.020 15.600 ;
      LAYER met2 ;
        RECT 2536.580 220.000 2536.860 224.000 ;
        RECT 2536.600 209.770 2536.740 220.000 ;
        RECT 2536.540 209.450 2536.800 209.770 ;
        RECT 2687.420 209.450 2687.680 209.770 ;
        RECT 2687.480 15.290 2687.620 209.450 ;
        RECT 2815.760 15.310 2816.020 15.630 ;
        RECT 2687.420 14.970 2687.680 15.290 ;
        RECT 2815.820 2.400 2815.960 15.310 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2590.865 14.025 2591.035 18.615 ;
      LAYER mcon ;
        RECT 2590.865 18.445 2591.035 18.615 ;
      LAYER met1 ;
        RECT 2590.805 18.600 2591.095 18.645 ;
        RECT 2833.670 18.600 2833.990 18.660 ;
        RECT 2590.805 18.460 2833.990 18.600 ;
        RECT 2590.805 18.415 2591.095 18.460 ;
        RECT 2833.670 18.400 2833.990 18.460 ;
        RECT 2552.610 14.180 2552.930 14.240 ;
        RECT 2590.805 14.180 2591.095 14.225 ;
        RECT 2552.610 14.040 2591.095 14.180 ;
        RECT 2552.610 13.980 2552.930 14.040 ;
        RECT 2590.805 13.995 2591.095 14.040 ;
      LAYER via ;
        RECT 2833.700 18.400 2833.960 18.660 ;
        RECT 2552.640 13.980 2552.900 14.240 ;
      LAYER met2 ;
        RECT 2550.840 220.730 2551.120 224.000 ;
        RECT 2550.840 220.590 2552.840 220.730 ;
        RECT 2550.840 220.000 2551.120 220.590 ;
        RECT 2552.700 14.270 2552.840 220.590 ;
        RECT 2833.700 18.370 2833.960 18.690 ;
        RECT 2552.640 13.950 2552.900 14.270 ;
        RECT 2833.760 2.400 2833.900 18.370 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2707.705 15.725 2709.715 15.895 ;
        RECT 2693.905 14.705 2694.075 15.555 ;
        RECT 2707.705 14.705 2707.875 15.725 ;
      LAYER mcon ;
        RECT 2709.545 15.725 2709.715 15.895 ;
        RECT 2693.905 15.385 2694.075 15.555 ;
      LAYER met1 ;
        RECT 2565.490 209.000 2565.810 209.060 ;
        RECT 2687.850 209.000 2688.170 209.060 ;
        RECT 2565.490 208.860 2688.170 209.000 ;
        RECT 2565.490 208.800 2565.810 208.860 ;
        RECT 2687.850 208.800 2688.170 208.860 ;
        RECT 2709.485 15.880 2709.775 15.925 ;
        RECT 2851.150 15.880 2851.470 15.940 ;
        RECT 2709.485 15.740 2851.470 15.880 ;
        RECT 2709.485 15.695 2709.775 15.740 ;
        RECT 2851.150 15.680 2851.470 15.740 ;
        RECT 2687.850 15.540 2688.170 15.600 ;
        RECT 2693.845 15.540 2694.135 15.585 ;
        RECT 2687.850 15.400 2694.135 15.540 ;
        RECT 2687.850 15.340 2688.170 15.400 ;
        RECT 2693.845 15.355 2694.135 15.400 ;
        RECT 2693.845 14.860 2694.135 14.905 ;
        RECT 2707.645 14.860 2707.935 14.905 ;
        RECT 2693.845 14.720 2707.935 14.860 ;
        RECT 2693.845 14.675 2694.135 14.720 ;
        RECT 2707.645 14.675 2707.935 14.720 ;
      LAYER via ;
        RECT 2565.520 208.800 2565.780 209.060 ;
        RECT 2687.880 208.800 2688.140 209.060 ;
        RECT 2851.180 15.680 2851.440 15.940 ;
        RECT 2687.880 15.340 2688.140 15.600 ;
      LAYER met2 ;
        RECT 2565.560 220.000 2565.840 224.000 ;
        RECT 2565.580 209.090 2565.720 220.000 ;
        RECT 2565.520 208.770 2565.780 209.090 ;
        RECT 2687.880 208.770 2688.140 209.090 ;
        RECT 2687.940 15.630 2688.080 208.770 ;
        RECT 2851.180 15.650 2851.440 15.970 ;
        RECT 2687.880 15.310 2688.140 15.630 ;
        RECT 2851.240 2.400 2851.380 15.650 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2580.210 18.260 2580.530 18.320 ;
        RECT 2580.210 18.120 2590.100 18.260 ;
        RECT 2580.210 18.060 2580.530 18.120 ;
        RECT 2589.960 17.920 2590.100 18.120 ;
        RECT 2869.090 17.920 2869.410 17.980 ;
        RECT 2589.960 17.780 2869.410 17.920 ;
        RECT 2869.090 17.720 2869.410 17.780 ;
      LAYER via ;
        RECT 2580.240 18.060 2580.500 18.320 ;
        RECT 2869.120 17.720 2869.380 17.980 ;
      LAYER met2 ;
        RECT 2580.280 220.000 2580.560 224.000 ;
        RECT 2580.300 18.350 2580.440 220.000 ;
        RECT 2580.240 18.030 2580.500 18.350 ;
        RECT 2869.120 17.690 2869.380 18.010 ;
        RECT 2869.180 2.400 2869.320 17.690 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2594.930 208.320 2595.250 208.380 ;
        RECT 2694.290 208.320 2694.610 208.380 ;
        RECT 2594.930 208.180 2694.610 208.320 ;
        RECT 2594.930 208.120 2595.250 208.180 ;
        RECT 2694.290 208.120 2694.610 208.180 ;
        RECT 2887.030 16.220 2887.350 16.280 ;
        RECT 2709.100 16.080 2887.350 16.220 ;
        RECT 2694.290 15.540 2694.610 15.600 ;
        RECT 2709.100 15.540 2709.240 16.080 ;
        RECT 2887.030 16.020 2887.350 16.080 ;
        RECT 2694.290 15.400 2709.240 15.540 ;
        RECT 2694.290 15.340 2694.610 15.400 ;
      LAYER via ;
        RECT 2594.960 208.120 2595.220 208.380 ;
        RECT 2694.320 208.120 2694.580 208.380 ;
        RECT 2694.320 15.340 2694.580 15.600 ;
        RECT 2887.060 16.020 2887.320 16.280 ;
      LAYER met2 ;
        RECT 2595.000 220.000 2595.280 224.000 ;
        RECT 2595.020 208.410 2595.160 220.000 ;
        RECT 2594.960 208.090 2595.220 208.410 ;
        RECT 2694.320 208.090 2694.580 208.410 ;
        RECT 2694.380 15.630 2694.520 208.090 ;
        RECT 2887.060 15.990 2887.320 16.310 ;
        RECT 2694.320 15.310 2694.580 15.630 ;
        RECT 2887.120 2.400 2887.260 15.990 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2609.650 207.300 2609.970 207.360 ;
        RECT 2614.710 207.300 2615.030 207.360 ;
        RECT 2609.650 207.160 2615.030 207.300 ;
        RECT 2609.650 207.100 2609.970 207.160 ;
        RECT 2614.710 207.100 2615.030 207.160 ;
        RECT 2614.710 17.240 2615.030 17.300 ;
        RECT 2904.970 17.240 2905.290 17.300 ;
        RECT 2614.710 17.100 2905.290 17.240 ;
        RECT 2614.710 17.040 2615.030 17.100 ;
        RECT 2904.970 17.040 2905.290 17.100 ;
      LAYER via ;
        RECT 2609.680 207.100 2609.940 207.360 ;
        RECT 2614.740 207.100 2615.000 207.360 ;
        RECT 2614.740 17.040 2615.000 17.300 ;
        RECT 2905.000 17.040 2905.260 17.300 ;
      LAYER met2 ;
        RECT 2609.720 220.000 2610.000 224.000 ;
        RECT 2609.740 207.390 2609.880 220.000 ;
        RECT 2609.680 207.070 2609.940 207.390 ;
        RECT 2614.740 207.070 2615.000 207.390 ;
        RECT 2614.800 17.330 2614.940 207.070 ;
        RECT 2614.740 17.010 2615.000 17.330 ;
        RECT 2905.000 17.010 2905.260 17.330 ;
        RECT 2905.060 2.400 2905.200 17.010 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 855.210 211.720 855.530 211.780 ;
        RECT 920.070 211.720 920.390 211.780 ;
        RECT 855.210 211.580 920.390 211.720 ;
        RECT 855.210 211.520 855.530 211.580 ;
        RECT 920.070 211.520 920.390 211.580 ;
        RECT 852.910 20.640 853.230 20.700 ;
        RECT 855.210 20.640 855.530 20.700 ;
        RECT 852.910 20.500 855.530 20.640 ;
        RECT 852.910 20.440 853.230 20.500 ;
        RECT 855.210 20.440 855.530 20.500 ;
      LAYER via ;
        RECT 855.240 211.520 855.500 211.780 ;
        RECT 920.100 211.520 920.360 211.780 ;
        RECT 852.940 20.440 853.200 20.700 ;
        RECT 855.240 20.440 855.500 20.700 ;
      LAYER met2 ;
        RECT 920.140 220.000 920.420 224.000 ;
        RECT 920.160 211.810 920.300 220.000 ;
        RECT 855.240 211.490 855.500 211.810 ;
        RECT 920.100 211.490 920.360 211.810 ;
        RECT 855.300 20.730 855.440 211.490 ;
        RECT 852.940 20.410 853.200 20.730 ;
        RECT 855.240 20.410 855.500 20.730 ;
        RECT 853.000 2.400 853.140 20.410 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 875.065 144.925 875.235 179.435 ;
      LAYER mcon ;
        RECT 875.065 179.265 875.235 179.435 ;
      LAYER met1 ;
        RECT 875.910 212.400 876.230 212.460 ;
        RECT 934.790 212.400 935.110 212.460 ;
        RECT 875.910 212.260 935.110 212.400 ;
        RECT 875.910 212.200 876.230 212.260 ;
        RECT 934.790 212.200 935.110 212.260 ;
        RECT 875.005 179.420 875.295 179.465 ;
        RECT 875.910 179.420 876.230 179.480 ;
        RECT 875.005 179.280 876.230 179.420 ;
        RECT 875.005 179.235 875.295 179.280 ;
        RECT 875.910 179.220 876.230 179.280 ;
        RECT 874.990 145.080 875.310 145.140 ;
        RECT 874.795 144.940 875.310 145.080 ;
        RECT 874.990 144.880 875.310 144.940 ;
        RECT 874.990 110.740 875.310 110.800 ;
        RECT 874.160 110.600 875.310 110.740 ;
        RECT 874.160 110.460 874.300 110.600 ;
        RECT 874.990 110.540 875.310 110.600 ;
        RECT 874.070 110.200 874.390 110.460 ;
        RECT 870.850 15.200 871.170 15.260 ;
        RECT 874.070 15.200 874.390 15.260 ;
        RECT 870.850 15.060 874.390 15.200 ;
        RECT 870.850 15.000 871.170 15.060 ;
        RECT 874.070 15.000 874.390 15.060 ;
      LAYER via ;
        RECT 875.940 212.200 876.200 212.460 ;
        RECT 934.820 212.200 935.080 212.460 ;
        RECT 875.940 179.220 876.200 179.480 ;
        RECT 875.020 144.880 875.280 145.140 ;
        RECT 875.020 110.540 875.280 110.800 ;
        RECT 874.100 110.200 874.360 110.460 ;
        RECT 870.880 15.000 871.140 15.260 ;
        RECT 874.100 15.000 874.360 15.260 ;
      LAYER met2 ;
        RECT 934.860 220.000 935.140 224.000 ;
        RECT 934.880 212.490 935.020 220.000 ;
        RECT 875.940 212.170 876.200 212.490 ;
        RECT 934.820 212.170 935.080 212.490 ;
        RECT 876.000 179.510 876.140 212.170 ;
        RECT 875.940 179.190 876.200 179.510 ;
        RECT 875.020 144.850 875.280 145.170 ;
        RECT 875.080 110.830 875.220 144.850 ;
        RECT 875.020 110.510 875.280 110.830 ;
        RECT 874.100 110.170 874.360 110.490 ;
        RECT 874.160 15.290 874.300 110.170 ;
        RECT 870.880 14.970 871.140 15.290 ;
        RECT 874.100 14.970 874.360 15.290 ;
        RECT 870.940 2.400 871.080 14.970 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 889.710 210.360 890.030 210.420 ;
        RECT 949.510 210.360 949.830 210.420 ;
        RECT 889.710 210.220 949.830 210.360 ;
        RECT 889.710 210.160 890.030 210.220 ;
        RECT 949.510 210.160 949.830 210.220 ;
      LAYER via ;
        RECT 889.740 210.160 890.000 210.420 ;
        RECT 949.540 210.160 949.800 210.420 ;
      LAYER met2 ;
        RECT 949.580 220.000 949.860 224.000 ;
        RECT 949.600 210.450 949.740 220.000 ;
        RECT 889.740 210.130 890.000 210.450 ;
        RECT 949.540 210.130 949.800 210.450 ;
        RECT 889.800 17.410 889.940 210.130 ;
        RECT 888.880 17.270 889.940 17.410 ;
        RECT 888.880 2.400 889.020 17.270 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 910.870 212.740 911.190 212.800 ;
        RECT 964.230 212.740 964.550 212.800 ;
        RECT 910.870 212.600 964.550 212.740 ;
        RECT 910.870 212.540 911.190 212.600 ;
        RECT 964.230 212.540 964.550 212.600 ;
        RECT 906.730 15.540 907.050 15.600 ;
        RECT 910.410 15.540 910.730 15.600 ;
        RECT 906.730 15.400 910.730 15.540 ;
        RECT 906.730 15.340 907.050 15.400 ;
        RECT 910.410 15.340 910.730 15.400 ;
      LAYER via ;
        RECT 910.900 212.540 911.160 212.800 ;
        RECT 964.260 212.540 964.520 212.800 ;
        RECT 906.760 15.340 907.020 15.600 ;
        RECT 910.440 15.340 910.700 15.600 ;
      LAYER met2 ;
        RECT 964.300 220.000 964.580 224.000 ;
        RECT 964.320 212.830 964.460 220.000 ;
        RECT 910.900 212.510 911.160 212.830 ;
        RECT 964.260 212.510 964.520 212.830 ;
        RECT 910.960 210.530 911.100 212.510 ;
        RECT 910.500 210.390 911.100 210.530 ;
        RECT 910.500 15.630 910.640 210.390 ;
        RECT 906.760 15.310 907.020 15.630 ;
        RECT 910.440 15.310 910.700 15.630 ;
        RECT 906.820 2.400 906.960 15.310 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 923.750 211.040 924.070 211.100 ;
        RECT 978.950 211.040 979.270 211.100 ;
        RECT 923.750 210.900 979.270 211.040 ;
        RECT 923.750 210.840 924.070 210.900 ;
        RECT 978.950 210.840 979.270 210.900 ;
      LAYER via ;
        RECT 923.780 210.840 924.040 211.100 ;
        RECT 978.980 210.840 979.240 211.100 ;
      LAYER met2 ;
        RECT 979.020 220.000 979.300 224.000 ;
        RECT 979.040 211.130 979.180 220.000 ;
        RECT 923.780 210.810 924.040 211.130 ;
        RECT 978.980 210.810 979.240 211.130 ;
        RECT 923.840 17.410 923.980 210.810 ;
        RECT 923.840 17.270 924.440 17.410 ;
        RECT 924.300 2.400 924.440 17.270 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 944.910 211.720 945.230 211.780 ;
        RECT 993.670 211.720 993.990 211.780 ;
        RECT 944.910 211.580 993.990 211.720 ;
        RECT 944.910 211.520 945.230 211.580 ;
        RECT 993.670 211.520 993.990 211.580 ;
        RECT 942.150 17.580 942.470 17.640 ;
        RECT 944.910 17.580 945.230 17.640 ;
        RECT 942.150 17.440 945.230 17.580 ;
        RECT 942.150 17.380 942.470 17.440 ;
        RECT 944.910 17.380 945.230 17.440 ;
      LAYER via ;
        RECT 944.940 211.520 945.200 211.780 ;
        RECT 993.700 211.520 993.960 211.780 ;
        RECT 942.180 17.380 942.440 17.640 ;
        RECT 944.940 17.380 945.200 17.640 ;
      LAYER met2 ;
        RECT 993.740 220.000 994.020 224.000 ;
        RECT 993.760 211.810 993.900 220.000 ;
        RECT 944.940 211.490 945.200 211.810 ;
        RECT 993.700 211.490 993.960 211.810 ;
        RECT 945.000 17.670 945.140 211.490 ;
        RECT 942.180 17.350 942.440 17.670 ;
        RECT 944.940 17.350 945.200 17.670 ;
        RECT 942.240 2.400 942.380 17.350 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 965.610 210.700 965.930 210.760 ;
        RECT 1008.390 210.700 1008.710 210.760 ;
        RECT 965.610 210.560 1008.710 210.700 ;
        RECT 965.610 210.500 965.930 210.560 ;
        RECT 1008.390 210.500 1008.710 210.560 ;
        RECT 960.090 17.580 960.410 17.640 ;
        RECT 965.610 17.580 965.930 17.640 ;
        RECT 960.090 17.440 965.930 17.580 ;
        RECT 960.090 17.380 960.410 17.440 ;
        RECT 965.610 17.380 965.930 17.440 ;
      LAYER via ;
        RECT 965.640 210.500 965.900 210.760 ;
        RECT 1008.420 210.500 1008.680 210.760 ;
        RECT 960.120 17.380 960.380 17.640 ;
        RECT 965.640 17.380 965.900 17.640 ;
      LAYER met2 ;
        RECT 1008.460 220.000 1008.740 224.000 ;
        RECT 1008.480 210.790 1008.620 220.000 ;
        RECT 965.640 210.470 965.900 210.790 ;
        RECT 1008.420 210.470 1008.680 210.790 ;
        RECT 965.700 17.670 965.840 210.470 ;
        RECT 960.120 17.350 960.380 17.670 ;
        RECT 965.640 17.350 965.900 17.670 ;
        RECT 960.180 2.400 960.320 17.350 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 979.410 211.040 979.730 211.100 ;
        RECT 1023.110 211.040 1023.430 211.100 ;
        RECT 979.410 210.900 1023.430 211.040 ;
        RECT 979.410 210.840 979.730 210.900 ;
        RECT 1023.110 210.840 1023.430 210.900 ;
      LAYER via ;
        RECT 979.440 210.840 979.700 211.100 ;
        RECT 1023.140 210.840 1023.400 211.100 ;
      LAYER met2 ;
        RECT 1023.180 220.000 1023.460 224.000 ;
        RECT 1023.200 211.130 1023.340 220.000 ;
        RECT 979.440 210.810 979.700 211.130 ;
        RECT 1023.140 210.810 1023.400 211.130 ;
        RECT 979.500 17.410 979.640 210.810 ;
        RECT 978.120 17.270 979.640 17.410 ;
        RECT 978.120 2.400 978.260 17.270 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 208.320 662.330 208.380 ;
        RECT 757.230 208.320 757.550 208.380 ;
        RECT 662.010 208.180 757.550 208.320 ;
        RECT 662.010 208.120 662.330 208.180 ;
        RECT 757.230 208.120 757.550 208.180 ;
        RECT 656.950 17.580 657.270 17.640 ;
        RECT 662.010 17.580 662.330 17.640 ;
        RECT 656.950 17.440 662.330 17.580 ;
        RECT 656.950 17.380 657.270 17.440 ;
        RECT 662.010 17.380 662.330 17.440 ;
      LAYER via ;
        RECT 662.040 208.120 662.300 208.380 ;
        RECT 757.260 208.120 757.520 208.380 ;
        RECT 656.980 17.380 657.240 17.640 ;
        RECT 662.040 17.380 662.300 17.640 ;
      LAYER met2 ;
        RECT 758.680 220.730 758.960 224.000 ;
        RECT 757.320 220.590 758.960 220.730 ;
        RECT 757.320 208.410 757.460 220.590 ;
        RECT 758.680 220.000 758.960 220.590 ;
        RECT 662.040 208.090 662.300 208.410 ;
        RECT 757.260 208.090 757.520 208.410 ;
        RECT 662.100 17.670 662.240 208.090 ;
        RECT 656.980 17.350 657.240 17.670 ;
        RECT 662.040 17.350 662.300 17.670 ;
        RECT 657.040 2.400 657.180 17.350 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1000.110 211.720 1000.430 211.780 ;
        RECT 1037.830 211.720 1038.150 211.780 ;
        RECT 1000.110 211.580 1038.150 211.720 ;
        RECT 1000.110 211.520 1000.430 211.580 ;
        RECT 1037.830 211.520 1038.150 211.580 ;
        RECT 995.970 17.580 996.290 17.640 ;
        RECT 1000.110 17.580 1000.430 17.640 ;
        RECT 995.970 17.440 1000.430 17.580 ;
        RECT 995.970 17.380 996.290 17.440 ;
        RECT 1000.110 17.380 1000.430 17.440 ;
      LAYER via ;
        RECT 1000.140 211.520 1000.400 211.780 ;
        RECT 1037.860 211.520 1038.120 211.780 ;
        RECT 996.000 17.380 996.260 17.640 ;
        RECT 1000.140 17.380 1000.400 17.640 ;
      LAYER met2 ;
        RECT 1037.900 220.000 1038.180 224.000 ;
        RECT 1037.920 211.810 1038.060 220.000 ;
        RECT 1000.140 211.490 1000.400 211.810 ;
        RECT 1037.860 211.490 1038.120 211.810 ;
        RECT 1000.200 17.670 1000.340 211.490 ;
        RECT 996.000 17.350 996.260 17.670 ;
        RECT 1000.140 17.350 1000.400 17.670 ;
        RECT 996.060 2.400 996.200 17.350 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 210.700 1014.230 210.760 ;
        RECT 1052.090 210.700 1052.410 210.760 ;
        RECT 1013.910 210.560 1052.410 210.700 ;
        RECT 1013.910 210.500 1014.230 210.560 ;
        RECT 1052.090 210.500 1052.410 210.560 ;
      LAYER via ;
        RECT 1013.940 210.500 1014.200 210.760 ;
        RECT 1052.120 210.500 1052.380 210.760 ;
      LAYER met2 ;
        RECT 1052.160 220.000 1052.440 224.000 ;
        RECT 1052.180 210.790 1052.320 220.000 ;
        RECT 1013.940 210.470 1014.200 210.790 ;
        RECT 1052.120 210.470 1052.380 210.790 ;
        RECT 1014.000 17.410 1014.140 210.470 ;
        RECT 1013.540 17.270 1014.140 17.410 ;
        RECT 1013.540 2.400 1013.680 17.270 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1034.610 211.040 1034.930 211.100 ;
        RECT 1066.810 211.040 1067.130 211.100 ;
        RECT 1034.610 210.900 1067.130 211.040 ;
        RECT 1034.610 210.840 1034.930 210.900 ;
        RECT 1066.810 210.840 1067.130 210.900 ;
        RECT 1031.390 15.200 1031.710 15.260 ;
        RECT 1034.610 15.200 1034.930 15.260 ;
        RECT 1031.390 15.060 1034.930 15.200 ;
        RECT 1031.390 15.000 1031.710 15.060 ;
        RECT 1034.610 15.000 1034.930 15.060 ;
      LAYER via ;
        RECT 1034.640 210.840 1034.900 211.100 ;
        RECT 1066.840 210.840 1067.100 211.100 ;
        RECT 1031.420 15.000 1031.680 15.260 ;
        RECT 1034.640 15.000 1034.900 15.260 ;
      LAYER met2 ;
        RECT 1066.880 220.000 1067.160 224.000 ;
        RECT 1066.900 211.130 1067.040 220.000 ;
        RECT 1034.640 210.810 1034.900 211.130 ;
        RECT 1066.840 210.810 1067.100 211.130 ;
        RECT 1034.700 15.290 1034.840 210.810 ;
        RECT 1031.420 14.970 1031.680 15.290 ;
        RECT 1034.640 14.970 1034.900 15.290 ;
        RECT 1031.480 2.400 1031.620 14.970 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1054.850 207.980 1055.170 208.040 ;
        RECT 1081.530 207.980 1081.850 208.040 ;
        RECT 1054.850 207.840 1081.850 207.980 ;
        RECT 1054.850 207.780 1055.170 207.840 ;
        RECT 1081.530 207.780 1081.850 207.840 ;
        RECT 1049.330 17.580 1049.650 17.640 ;
        RECT 1054.850 17.580 1055.170 17.640 ;
        RECT 1049.330 17.440 1055.170 17.580 ;
        RECT 1049.330 17.380 1049.650 17.440 ;
        RECT 1054.850 17.380 1055.170 17.440 ;
      LAYER via ;
        RECT 1054.880 207.780 1055.140 208.040 ;
        RECT 1081.560 207.780 1081.820 208.040 ;
        RECT 1049.360 17.380 1049.620 17.640 ;
        RECT 1054.880 17.380 1055.140 17.640 ;
      LAYER met2 ;
        RECT 1081.600 220.000 1081.880 224.000 ;
        RECT 1081.620 208.070 1081.760 220.000 ;
        RECT 1054.880 207.750 1055.140 208.070 ;
        RECT 1081.560 207.750 1081.820 208.070 ;
        RECT 1054.940 17.670 1055.080 207.750 ;
        RECT 1049.360 17.350 1049.620 17.670 ;
        RECT 1054.880 17.350 1055.140 17.670 ;
        RECT 1049.420 2.400 1049.560 17.350 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1069.110 211.040 1069.430 211.100 ;
        RECT 1096.250 211.040 1096.570 211.100 ;
        RECT 1069.110 210.900 1096.570 211.040 ;
        RECT 1069.110 210.840 1069.430 210.900 ;
        RECT 1096.250 210.840 1096.570 210.900 ;
      LAYER via ;
        RECT 1069.140 210.840 1069.400 211.100 ;
        RECT 1096.280 210.840 1096.540 211.100 ;
      LAYER met2 ;
        RECT 1096.320 220.000 1096.600 224.000 ;
        RECT 1096.340 211.130 1096.480 220.000 ;
        RECT 1069.140 210.810 1069.400 211.130 ;
        RECT 1096.280 210.810 1096.540 211.130 ;
        RECT 1069.200 17.410 1069.340 210.810 ;
        RECT 1067.360 17.270 1069.340 17.410 ;
        RECT 1067.360 2.400 1067.500 17.270 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1089.810 210.700 1090.130 210.760 ;
        RECT 1110.970 210.700 1111.290 210.760 ;
        RECT 1089.810 210.560 1111.290 210.700 ;
        RECT 1089.810 210.500 1090.130 210.560 ;
        RECT 1110.970 210.500 1111.290 210.560 ;
        RECT 1085.210 17.580 1085.530 17.640 ;
        RECT 1089.810 17.580 1090.130 17.640 ;
        RECT 1085.210 17.440 1090.130 17.580 ;
        RECT 1085.210 17.380 1085.530 17.440 ;
        RECT 1089.810 17.380 1090.130 17.440 ;
      LAYER via ;
        RECT 1089.840 210.500 1090.100 210.760 ;
        RECT 1111.000 210.500 1111.260 210.760 ;
        RECT 1085.240 17.380 1085.500 17.640 ;
        RECT 1089.840 17.380 1090.100 17.640 ;
      LAYER met2 ;
        RECT 1111.040 220.000 1111.320 224.000 ;
        RECT 1111.060 210.790 1111.200 220.000 ;
        RECT 1089.840 210.470 1090.100 210.790 ;
        RECT 1111.000 210.470 1111.260 210.790 ;
        RECT 1089.900 17.670 1090.040 210.470 ;
        RECT 1085.240 17.350 1085.500 17.670 ;
        RECT 1089.840 17.350 1090.100 17.670 ;
        RECT 1085.300 2.400 1085.440 17.350 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1103.610 208.320 1103.930 208.380 ;
        RECT 1125.690 208.320 1126.010 208.380 ;
        RECT 1103.610 208.180 1126.010 208.320 ;
        RECT 1103.610 208.120 1103.930 208.180 ;
        RECT 1125.690 208.120 1126.010 208.180 ;
      LAYER via ;
        RECT 1103.640 208.120 1103.900 208.380 ;
        RECT 1125.720 208.120 1125.980 208.380 ;
      LAYER met2 ;
        RECT 1125.760 220.000 1126.040 224.000 ;
        RECT 1125.780 208.410 1125.920 220.000 ;
        RECT 1103.640 208.090 1103.900 208.410 ;
        RECT 1125.720 208.090 1125.980 208.410 ;
        RECT 1103.700 17.410 1103.840 208.090 ;
        RECT 1102.780 17.270 1103.840 17.410 ;
        RECT 1102.780 2.400 1102.920 17.270 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1124.310 207.980 1124.630 208.040 ;
        RECT 1140.410 207.980 1140.730 208.040 ;
        RECT 1124.310 207.840 1140.730 207.980 ;
        RECT 1124.310 207.780 1124.630 207.840 ;
        RECT 1140.410 207.780 1140.730 207.840 ;
        RECT 1120.630 17.580 1120.950 17.640 ;
        RECT 1124.310 17.580 1124.630 17.640 ;
        RECT 1120.630 17.440 1124.630 17.580 ;
        RECT 1120.630 17.380 1120.950 17.440 ;
        RECT 1124.310 17.380 1124.630 17.440 ;
      LAYER via ;
        RECT 1124.340 207.780 1124.600 208.040 ;
        RECT 1140.440 207.780 1140.700 208.040 ;
        RECT 1120.660 17.380 1120.920 17.640 ;
        RECT 1124.340 17.380 1124.600 17.640 ;
      LAYER met2 ;
        RECT 1140.480 220.000 1140.760 224.000 ;
        RECT 1140.500 208.070 1140.640 220.000 ;
        RECT 1124.340 207.750 1124.600 208.070 ;
        RECT 1140.440 207.750 1140.700 208.070 ;
        RECT 1124.400 17.670 1124.540 207.750 ;
        RECT 1120.660 17.350 1120.920 17.670 ;
        RECT 1124.340 17.350 1124.600 17.670 ;
        RECT 1120.720 2.400 1120.860 17.350 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1138.570 18.600 1138.890 18.660 ;
        RECT 1152.830 18.600 1153.150 18.660 ;
        RECT 1138.570 18.460 1153.150 18.600 ;
        RECT 1138.570 18.400 1138.890 18.460 ;
        RECT 1152.830 18.400 1153.150 18.460 ;
      LAYER via ;
        RECT 1138.600 18.400 1138.860 18.660 ;
        RECT 1152.860 18.400 1153.120 18.660 ;
      LAYER met2 ;
        RECT 1155.200 220.730 1155.480 224.000 ;
        RECT 1152.920 220.590 1155.480 220.730 ;
        RECT 1152.920 18.690 1153.060 220.590 ;
        RECT 1155.200 220.000 1155.480 220.590 ;
        RECT 1138.600 18.370 1138.860 18.690 ;
        RECT 1152.860 18.370 1153.120 18.690 ;
        RECT 1138.660 2.400 1138.800 18.370 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1158.810 207.300 1159.130 207.360 ;
        RECT 1169.850 207.300 1170.170 207.360 ;
        RECT 1158.810 207.160 1170.170 207.300 ;
        RECT 1158.810 207.100 1159.130 207.160 ;
        RECT 1169.850 207.100 1170.170 207.160 ;
        RECT 1156.510 17.580 1156.830 17.640 ;
        RECT 1158.810 17.580 1159.130 17.640 ;
        RECT 1156.510 17.440 1159.130 17.580 ;
        RECT 1156.510 17.380 1156.830 17.440 ;
        RECT 1158.810 17.380 1159.130 17.440 ;
      LAYER via ;
        RECT 1158.840 207.100 1159.100 207.360 ;
        RECT 1169.880 207.100 1170.140 207.360 ;
        RECT 1156.540 17.380 1156.800 17.640 ;
        RECT 1158.840 17.380 1159.100 17.640 ;
      LAYER met2 ;
        RECT 1169.920 220.000 1170.200 224.000 ;
        RECT 1169.940 207.390 1170.080 220.000 ;
        RECT 1158.840 207.070 1159.100 207.390 ;
        RECT 1169.880 207.070 1170.140 207.390 ;
        RECT 1158.900 17.670 1159.040 207.070 ;
        RECT 1156.540 17.350 1156.800 17.670 ;
        RECT 1158.840 17.350 1159.100 17.670 ;
        RECT 1156.600 2.400 1156.740 17.350 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 680.945 209.185 681.115 213.095 ;
      LAYER mcon ;
        RECT 680.945 212.925 681.115 213.095 ;
      LAYER met1 ;
        RECT 680.885 213.080 681.175 213.125 ;
        RECT 773.330 213.080 773.650 213.140 ;
        RECT 680.885 212.940 773.650 213.080 ;
        RECT 680.885 212.895 681.175 212.940 ;
        RECT 773.330 212.880 773.650 212.940 ;
        RECT 675.810 209.340 676.130 209.400 ;
        RECT 680.885 209.340 681.175 209.385 ;
        RECT 675.810 209.200 681.175 209.340 ;
        RECT 675.810 209.140 676.130 209.200 ;
        RECT 680.885 209.155 681.175 209.200 ;
      LAYER via ;
        RECT 773.360 212.880 773.620 213.140 ;
        RECT 675.840 209.140 676.100 209.400 ;
      LAYER met2 ;
        RECT 773.400 220.000 773.680 224.000 ;
        RECT 773.420 213.170 773.560 220.000 ;
        RECT 773.360 212.850 773.620 213.170 ;
        RECT 675.840 209.110 676.100 209.430 ;
        RECT 675.900 17.410 676.040 209.110 ;
        RECT 674.520 17.270 676.040 17.410 ;
        RECT 674.520 2.400 674.660 17.270 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1173.990 17.580 1174.310 17.640 ;
        RECT 1180.890 17.580 1181.210 17.640 ;
        RECT 1173.990 17.440 1181.210 17.580 ;
        RECT 1173.990 17.380 1174.310 17.440 ;
        RECT 1180.890 17.380 1181.210 17.440 ;
      LAYER via ;
        RECT 1174.020 17.380 1174.280 17.640 ;
        RECT 1180.920 17.380 1181.180 17.640 ;
      LAYER met2 ;
        RECT 1184.640 220.730 1184.920 224.000 ;
        RECT 1180.980 220.590 1184.920 220.730 ;
        RECT 1180.980 17.670 1181.120 220.590 ;
        RECT 1184.640 220.000 1184.920 220.590 ;
        RECT 1174.020 17.350 1174.280 17.670 ;
        RECT 1180.920 17.350 1181.180 17.670 ;
        RECT 1174.080 2.400 1174.220 17.350 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1194.230 200.160 1194.550 200.220 ;
        RECT 1197.910 200.160 1198.230 200.220 ;
        RECT 1194.230 200.020 1198.230 200.160 ;
        RECT 1194.230 199.960 1194.550 200.020 ;
        RECT 1197.910 199.960 1198.230 200.020 ;
        RECT 1191.930 20.640 1192.250 20.700 ;
        RECT 1194.230 20.640 1194.550 20.700 ;
        RECT 1191.930 20.500 1194.550 20.640 ;
        RECT 1191.930 20.440 1192.250 20.500 ;
        RECT 1194.230 20.440 1194.550 20.500 ;
      LAYER via ;
        RECT 1194.260 199.960 1194.520 200.220 ;
        RECT 1197.940 199.960 1198.200 200.220 ;
        RECT 1191.960 20.440 1192.220 20.700 ;
        RECT 1194.260 20.440 1194.520 20.700 ;
      LAYER met2 ;
        RECT 1199.360 220.730 1199.640 224.000 ;
        RECT 1198.000 220.590 1199.640 220.730 ;
        RECT 1198.000 200.250 1198.140 220.590 ;
        RECT 1199.360 220.000 1199.640 220.590 ;
        RECT 1194.260 199.930 1194.520 200.250 ;
        RECT 1197.940 199.930 1198.200 200.250 ;
        RECT 1194.320 20.730 1194.460 199.930 ;
        RECT 1191.960 20.410 1192.220 20.730 ;
        RECT 1194.260 20.410 1194.520 20.730 ;
        RECT 1192.020 2.400 1192.160 20.410 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1208.030 179.760 1208.350 179.820 ;
        RECT 1212.630 179.760 1212.950 179.820 ;
        RECT 1208.030 179.620 1212.950 179.760 ;
        RECT 1208.030 179.560 1208.350 179.620 ;
        RECT 1212.630 179.560 1212.950 179.620 ;
      LAYER via ;
        RECT 1208.060 179.560 1208.320 179.820 ;
        RECT 1212.660 179.560 1212.920 179.820 ;
      LAYER met2 ;
        RECT 1214.080 220.730 1214.360 224.000 ;
        RECT 1212.720 220.590 1214.360 220.730 ;
        RECT 1212.720 179.850 1212.860 220.590 ;
        RECT 1214.080 220.000 1214.360 220.590 ;
        RECT 1208.060 179.530 1208.320 179.850 ;
        RECT 1212.660 179.530 1212.920 179.850 ;
        RECT 1208.120 24.210 1208.260 179.530 ;
        RECT 1208.120 24.070 1210.100 24.210 ;
        RECT 1209.960 2.400 1210.100 24.070 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1228.800 220.000 1229.080 224.000 ;
        RECT 1228.820 213.930 1228.960 220.000 ;
        RECT 1227.900 213.790 1228.960 213.930 ;
        RECT 1227.900 2.400 1228.040 213.790 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1242.530 20.640 1242.850 20.700 ;
        RECT 1245.750 20.640 1246.070 20.700 ;
        RECT 1242.530 20.500 1246.070 20.640 ;
        RECT 1242.530 20.440 1242.850 20.500 ;
        RECT 1245.750 20.440 1246.070 20.500 ;
      LAYER via ;
        RECT 1242.560 20.440 1242.820 20.700 ;
        RECT 1245.780 20.440 1246.040 20.700 ;
      LAYER met2 ;
        RECT 1243.520 220.730 1243.800 224.000 ;
        RECT 1242.620 220.590 1243.800 220.730 ;
        RECT 1242.620 20.730 1242.760 220.590 ;
        RECT 1243.520 220.000 1243.800 220.590 ;
        RECT 1242.560 20.410 1242.820 20.730 ;
        RECT 1245.780 20.410 1246.040 20.730 ;
        RECT 1245.840 2.400 1245.980 20.410 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1258.170 213.760 1258.490 213.820 ;
        RECT 1262.310 213.760 1262.630 213.820 ;
        RECT 1258.170 213.620 1262.630 213.760 ;
        RECT 1258.170 213.560 1258.490 213.620 ;
        RECT 1262.310 213.560 1262.630 213.620 ;
        RECT 1261.390 62.120 1261.710 62.180 ;
        RECT 1262.310 62.120 1262.630 62.180 ;
        RECT 1261.390 61.980 1262.630 62.120 ;
        RECT 1261.390 61.920 1261.710 61.980 ;
        RECT 1262.310 61.920 1262.630 61.980 ;
        RECT 1261.390 20.300 1261.710 20.360 ;
        RECT 1263.230 20.300 1263.550 20.360 ;
        RECT 1261.390 20.160 1263.550 20.300 ;
        RECT 1261.390 20.100 1261.710 20.160 ;
        RECT 1263.230 20.100 1263.550 20.160 ;
      LAYER via ;
        RECT 1258.200 213.560 1258.460 213.820 ;
        RECT 1262.340 213.560 1262.600 213.820 ;
        RECT 1261.420 61.920 1261.680 62.180 ;
        RECT 1262.340 61.920 1262.600 62.180 ;
        RECT 1261.420 20.100 1261.680 20.360 ;
        RECT 1263.260 20.100 1263.520 20.360 ;
      LAYER met2 ;
        RECT 1258.240 220.000 1258.520 224.000 ;
        RECT 1258.260 213.850 1258.400 220.000 ;
        RECT 1258.200 213.530 1258.460 213.850 ;
        RECT 1262.340 213.530 1262.600 213.850 ;
        RECT 1262.400 62.210 1262.540 213.530 ;
        RECT 1261.420 61.890 1261.680 62.210 ;
        RECT 1262.340 61.890 1262.600 62.210 ;
        RECT 1261.480 20.390 1261.620 61.890 ;
        RECT 1261.420 20.070 1261.680 20.390 ;
        RECT 1263.260 20.070 1263.520 20.390 ;
        RECT 1263.320 2.400 1263.460 20.070 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1276.110 17.580 1276.430 17.640 ;
        RECT 1281.170 17.580 1281.490 17.640 ;
        RECT 1276.110 17.440 1281.490 17.580 ;
        RECT 1276.110 17.380 1276.430 17.440 ;
        RECT 1281.170 17.380 1281.490 17.440 ;
      LAYER via ;
        RECT 1276.140 17.380 1276.400 17.640 ;
        RECT 1281.200 17.380 1281.460 17.640 ;
      LAYER met2 ;
        RECT 1272.960 220.730 1273.240 224.000 ;
        RECT 1272.960 220.590 1276.340 220.730 ;
        RECT 1272.960 220.000 1273.240 220.590 ;
        RECT 1276.200 17.670 1276.340 220.590 ;
        RECT 1276.140 17.350 1276.400 17.670 ;
        RECT 1281.200 17.350 1281.460 17.670 ;
        RECT 1281.260 2.400 1281.400 17.350 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1287.610 207.640 1287.930 207.700 ;
        RECT 1293.590 207.640 1293.910 207.700 ;
        RECT 1287.610 207.500 1293.910 207.640 ;
        RECT 1287.610 207.440 1287.930 207.500 ;
        RECT 1293.590 207.440 1293.910 207.500 ;
        RECT 1293.590 17.580 1293.910 17.640 ;
        RECT 1299.110 17.580 1299.430 17.640 ;
        RECT 1293.590 17.440 1299.430 17.580 ;
        RECT 1293.590 17.380 1293.910 17.440 ;
        RECT 1299.110 17.380 1299.430 17.440 ;
      LAYER via ;
        RECT 1287.640 207.440 1287.900 207.700 ;
        RECT 1293.620 207.440 1293.880 207.700 ;
        RECT 1293.620 17.380 1293.880 17.640 ;
        RECT 1299.140 17.380 1299.400 17.640 ;
      LAYER met2 ;
        RECT 1287.680 220.000 1287.960 224.000 ;
        RECT 1287.700 207.730 1287.840 220.000 ;
        RECT 1287.640 207.410 1287.900 207.730 ;
        RECT 1293.620 207.410 1293.880 207.730 ;
        RECT 1293.680 17.670 1293.820 207.410 ;
        RECT 1293.620 17.350 1293.880 17.670 ;
        RECT 1299.140 17.350 1299.400 17.670 ;
        RECT 1299.200 2.400 1299.340 17.350 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1303.710 16.900 1304.030 16.960 ;
        RECT 1317.050 16.900 1317.370 16.960 ;
        RECT 1303.710 16.760 1317.370 16.900 ;
        RECT 1303.710 16.700 1304.030 16.760 ;
        RECT 1317.050 16.700 1317.370 16.760 ;
      LAYER via ;
        RECT 1303.740 16.700 1304.000 16.960 ;
        RECT 1317.080 16.700 1317.340 16.960 ;
      LAYER met2 ;
        RECT 1301.940 220.730 1302.220 224.000 ;
        RECT 1301.940 220.590 1303.940 220.730 ;
        RECT 1301.940 220.000 1302.220 220.590 ;
        RECT 1303.800 16.990 1303.940 220.590 ;
        RECT 1303.740 16.670 1304.000 16.990 ;
        RECT 1317.080 16.670 1317.340 16.990 ;
        RECT 1317.140 2.400 1317.280 16.670 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.510 17.920 1317.830 17.980 ;
        RECT 1334.990 17.920 1335.310 17.980 ;
        RECT 1317.510 17.780 1335.310 17.920 ;
        RECT 1317.510 17.720 1317.830 17.780 ;
        RECT 1334.990 17.720 1335.310 17.780 ;
      LAYER via ;
        RECT 1317.540 17.720 1317.800 17.980 ;
        RECT 1335.020 17.720 1335.280 17.980 ;
      LAYER met2 ;
        RECT 1316.660 220.730 1316.940 224.000 ;
        RECT 1316.660 220.590 1317.740 220.730 ;
        RECT 1316.660 220.000 1316.940 220.590 ;
        RECT 1317.600 18.010 1317.740 220.590 ;
        RECT 1317.540 17.690 1317.800 18.010 ;
        RECT 1335.020 17.690 1335.280 18.010 ;
        RECT 1335.080 2.400 1335.220 17.690 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 696.510 212.400 696.830 212.460 ;
        RECT 788.050 212.400 788.370 212.460 ;
        RECT 696.510 212.260 788.370 212.400 ;
        RECT 696.510 212.200 696.830 212.260 ;
        RECT 788.050 212.200 788.370 212.260 ;
        RECT 692.370 17.580 692.690 17.640 ;
        RECT 696.510 17.580 696.830 17.640 ;
        RECT 692.370 17.440 696.830 17.580 ;
        RECT 692.370 17.380 692.690 17.440 ;
        RECT 696.510 17.380 696.830 17.440 ;
      LAYER via ;
        RECT 696.540 212.200 696.800 212.460 ;
        RECT 788.080 212.200 788.340 212.460 ;
        RECT 692.400 17.380 692.660 17.640 ;
        RECT 696.540 17.380 696.800 17.640 ;
      LAYER met2 ;
        RECT 788.120 220.000 788.400 224.000 ;
        RECT 788.140 212.490 788.280 220.000 ;
        RECT 696.540 212.170 696.800 212.490 ;
        RECT 788.080 212.170 788.340 212.490 ;
        RECT 696.600 17.670 696.740 212.170 ;
        RECT 692.400 17.350 692.660 17.670 ;
        RECT 696.540 17.350 696.800 17.670 ;
        RECT 692.460 2.400 692.600 17.350 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1331.310 17.580 1331.630 17.640 ;
        RECT 1352.470 17.580 1352.790 17.640 ;
        RECT 1331.310 17.440 1352.790 17.580 ;
        RECT 1331.310 17.380 1331.630 17.440 ;
        RECT 1352.470 17.380 1352.790 17.440 ;
      LAYER via ;
        RECT 1331.340 17.380 1331.600 17.640 ;
        RECT 1352.500 17.380 1352.760 17.640 ;
      LAYER met2 ;
        RECT 1331.380 220.000 1331.660 224.000 ;
        RECT 1331.400 17.670 1331.540 220.000 ;
        RECT 1331.340 17.350 1331.600 17.670 ;
        RECT 1352.500 17.350 1352.760 17.670 ;
        RECT 1352.560 2.400 1352.700 17.350 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1346.030 207.300 1346.350 207.360 ;
        RECT 1352.010 207.300 1352.330 207.360 ;
        RECT 1346.030 207.160 1352.330 207.300 ;
        RECT 1346.030 207.100 1346.350 207.160 ;
        RECT 1352.010 207.100 1352.330 207.160 ;
        RECT 1352.010 17.920 1352.330 17.980 ;
        RECT 1370.410 17.920 1370.730 17.980 ;
        RECT 1352.010 17.780 1370.730 17.920 ;
        RECT 1352.010 17.720 1352.330 17.780 ;
        RECT 1370.410 17.720 1370.730 17.780 ;
      LAYER via ;
        RECT 1346.060 207.100 1346.320 207.360 ;
        RECT 1352.040 207.100 1352.300 207.360 ;
        RECT 1352.040 17.720 1352.300 17.980 ;
        RECT 1370.440 17.720 1370.700 17.980 ;
      LAYER met2 ;
        RECT 1346.100 220.000 1346.380 224.000 ;
        RECT 1346.120 207.390 1346.260 220.000 ;
        RECT 1346.060 207.070 1346.320 207.390 ;
        RECT 1352.040 207.070 1352.300 207.390 ;
        RECT 1352.100 18.010 1352.240 207.070 ;
        RECT 1352.040 17.690 1352.300 18.010 ;
        RECT 1370.440 17.690 1370.700 18.010 ;
        RECT 1370.500 2.400 1370.640 17.690 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1360.750 207.300 1361.070 207.360 ;
        RECT 1365.350 207.300 1365.670 207.360 ;
        RECT 1360.750 207.160 1365.670 207.300 ;
        RECT 1360.750 207.100 1361.070 207.160 ;
        RECT 1365.350 207.100 1365.670 207.160 ;
        RECT 1365.350 15.540 1365.670 15.600 ;
        RECT 1388.350 15.540 1388.670 15.600 ;
        RECT 1365.350 15.400 1388.670 15.540 ;
        RECT 1365.350 15.340 1365.670 15.400 ;
        RECT 1388.350 15.340 1388.670 15.400 ;
      LAYER via ;
        RECT 1360.780 207.100 1361.040 207.360 ;
        RECT 1365.380 207.100 1365.640 207.360 ;
        RECT 1365.380 15.340 1365.640 15.600 ;
        RECT 1388.380 15.340 1388.640 15.600 ;
      LAYER met2 ;
        RECT 1360.820 220.000 1361.100 224.000 ;
        RECT 1360.840 207.390 1360.980 220.000 ;
        RECT 1360.780 207.070 1361.040 207.390 ;
        RECT 1365.380 207.070 1365.640 207.390 ;
        RECT 1365.440 15.630 1365.580 207.070 ;
        RECT 1365.380 15.310 1365.640 15.630 ;
        RECT 1388.380 15.310 1388.640 15.630 ;
        RECT 1388.440 2.400 1388.580 15.310 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1375.470 207.300 1375.790 207.360 ;
        RECT 1379.610 207.300 1379.930 207.360 ;
        RECT 1375.470 207.160 1379.930 207.300 ;
        RECT 1375.470 207.100 1375.790 207.160 ;
        RECT 1379.610 207.100 1379.930 207.160 ;
        RECT 1379.610 18.260 1379.930 18.320 ;
        RECT 1406.290 18.260 1406.610 18.320 ;
        RECT 1379.610 18.120 1406.610 18.260 ;
        RECT 1379.610 18.060 1379.930 18.120 ;
        RECT 1406.290 18.060 1406.610 18.120 ;
      LAYER via ;
        RECT 1375.500 207.100 1375.760 207.360 ;
        RECT 1379.640 207.100 1379.900 207.360 ;
        RECT 1379.640 18.060 1379.900 18.320 ;
        RECT 1406.320 18.060 1406.580 18.320 ;
      LAYER met2 ;
        RECT 1375.540 220.000 1375.820 224.000 ;
        RECT 1375.560 207.390 1375.700 220.000 ;
        RECT 1375.500 207.070 1375.760 207.390 ;
        RECT 1379.640 207.070 1379.900 207.390 ;
        RECT 1379.700 18.350 1379.840 207.070 ;
        RECT 1379.640 18.030 1379.900 18.350 ;
        RECT 1406.320 18.030 1406.580 18.350 ;
        RECT 1406.380 2.400 1406.520 18.030 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1393.410 16.560 1393.730 16.620 ;
        RECT 1423.770 16.560 1424.090 16.620 ;
        RECT 1393.410 16.420 1424.090 16.560 ;
        RECT 1393.410 16.360 1393.730 16.420 ;
        RECT 1423.770 16.360 1424.090 16.420 ;
      LAYER via ;
        RECT 1393.440 16.360 1393.700 16.620 ;
        RECT 1423.800 16.360 1424.060 16.620 ;
      LAYER met2 ;
        RECT 1390.260 220.730 1390.540 224.000 ;
        RECT 1390.260 220.590 1393.640 220.730 ;
        RECT 1390.260 220.000 1390.540 220.590 ;
        RECT 1393.500 16.650 1393.640 220.590 ;
        RECT 1393.440 16.330 1393.700 16.650 ;
        RECT 1423.800 16.330 1424.060 16.650 ;
        RECT 1423.860 2.400 1424.000 16.330 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1407.210 16.900 1407.530 16.960 ;
        RECT 1441.710 16.900 1442.030 16.960 ;
        RECT 1407.210 16.760 1442.030 16.900 ;
        RECT 1407.210 16.700 1407.530 16.760 ;
        RECT 1441.710 16.700 1442.030 16.760 ;
      LAYER via ;
        RECT 1407.240 16.700 1407.500 16.960 ;
        RECT 1441.740 16.700 1442.000 16.960 ;
      LAYER met2 ;
        RECT 1404.980 220.730 1405.260 224.000 ;
        RECT 1404.980 220.590 1407.440 220.730 ;
        RECT 1404.980 220.000 1405.260 220.590 ;
        RECT 1407.300 16.990 1407.440 220.590 ;
        RECT 1407.240 16.670 1407.500 16.990 ;
        RECT 1441.740 16.670 1442.000 16.990 ;
        RECT 1441.800 2.400 1441.940 16.670 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1421.010 18.940 1421.330 19.000 ;
        RECT 1459.650 18.940 1459.970 19.000 ;
        RECT 1421.010 18.800 1459.970 18.940 ;
        RECT 1421.010 18.740 1421.330 18.800 ;
        RECT 1459.650 18.740 1459.970 18.800 ;
      LAYER via ;
        RECT 1421.040 18.740 1421.300 19.000 ;
        RECT 1459.680 18.740 1459.940 19.000 ;
      LAYER met2 ;
        RECT 1419.700 220.730 1419.980 224.000 ;
        RECT 1419.700 220.590 1421.240 220.730 ;
        RECT 1419.700 220.000 1419.980 220.590 ;
        RECT 1421.100 19.030 1421.240 220.590 ;
        RECT 1421.040 18.710 1421.300 19.030 ;
        RECT 1459.680 18.710 1459.940 19.030 ;
        RECT 1459.740 2.400 1459.880 18.710 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1434.810 17.240 1435.130 17.300 ;
        RECT 1477.590 17.240 1477.910 17.300 ;
        RECT 1434.810 17.100 1477.910 17.240 ;
        RECT 1434.810 17.040 1435.130 17.100 ;
        RECT 1477.590 17.040 1477.910 17.100 ;
      LAYER via ;
        RECT 1434.840 17.040 1435.100 17.300 ;
        RECT 1477.620 17.040 1477.880 17.300 ;
      LAYER met2 ;
        RECT 1434.420 220.730 1434.700 224.000 ;
        RECT 1434.420 220.590 1435.040 220.730 ;
        RECT 1434.420 220.000 1434.700 220.590 ;
        RECT 1434.900 17.330 1435.040 220.590 ;
        RECT 1434.840 17.010 1435.100 17.330 ;
        RECT 1477.620 17.010 1477.880 17.330 ;
        RECT 1477.680 2.400 1477.820 17.010 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1449.070 207.300 1449.390 207.360 ;
        RECT 1455.510 207.300 1455.830 207.360 ;
        RECT 1449.070 207.160 1455.830 207.300 ;
        RECT 1449.070 207.100 1449.390 207.160 ;
        RECT 1455.510 207.100 1455.830 207.160 ;
        RECT 1455.510 14.860 1455.830 14.920 ;
        RECT 1495.530 14.860 1495.850 14.920 ;
        RECT 1455.510 14.720 1495.850 14.860 ;
        RECT 1455.510 14.660 1455.830 14.720 ;
        RECT 1495.530 14.660 1495.850 14.720 ;
      LAYER via ;
        RECT 1449.100 207.100 1449.360 207.360 ;
        RECT 1455.540 207.100 1455.800 207.360 ;
        RECT 1455.540 14.660 1455.800 14.920 ;
        RECT 1495.560 14.660 1495.820 14.920 ;
      LAYER met2 ;
        RECT 1449.140 220.000 1449.420 224.000 ;
        RECT 1449.160 207.390 1449.300 220.000 ;
        RECT 1449.100 207.070 1449.360 207.390 ;
        RECT 1455.540 207.070 1455.800 207.390 ;
        RECT 1455.600 14.950 1455.740 207.070 ;
        RECT 1455.540 14.630 1455.800 14.950 ;
        RECT 1495.560 14.630 1495.820 14.950 ;
        RECT 1495.620 2.400 1495.760 14.630 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1463.790 207.300 1464.110 207.360 ;
        RECT 1468.850 207.300 1469.170 207.360 ;
        RECT 1463.790 207.160 1469.170 207.300 ;
        RECT 1463.790 207.100 1464.110 207.160 ;
        RECT 1468.850 207.100 1469.170 207.160 ;
        RECT 1468.850 19.280 1469.170 19.340 ;
        RECT 1513.010 19.280 1513.330 19.340 ;
        RECT 1468.850 19.140 1513.330 19.280 ;
        RECT 1468.850 19.080 1469.170 19.140 ;
        RECT 1513.010 19.080 1513.330 19.140 ;
      LAYER via ;
        RECT 1463.820 207.100 1464.080 207.360 ;
        RECT 1468.880 207.100 1469.140 207.360 ;
        RECT 1468.880 19.080 1469.140 19.340 ;
        RECT 1513.040 19.080 1513.300 19.340 ;
      LAYER met2 ;
        RECT 1463.860 220.000 1464.140 224.000 ;
        RECT 1463.880 207.390 1464.020 220.000 ;
        RECT 1463.820 207.070 1464.080 207.390 ;
        RECT 1468.880 207.070 1469.140 207.390 ;
        RECT 1468.940 19.370 1469.080 207.070 ;
        RECT 1468.880 19.050 1469.140 19.370 ;
        RECT 1513.040 19.050 1513.300 19.370 ;
        RECT 1513.100 2.400 1513.240 19.050 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 710.310 210.360 710.630 210.420 ;
        RECT 802.310 210.360 802.630 210.420 ;
        RECT 710.310 210.220 802.630 210.360 ;
        RECT 710.310 210.160 710.630 210.220 ;
        RECT 802.310 210.160 802.630 210.220 ;
      LAYER via ;
        RECT 710.340 210.160 710.600 210.420 ;
        RECT 802.340 210.160 802.600 210.420 ;
      LAYER met2 ;
        RECT 802.380 220.000 802.660 224.000 ;
        RECT 802.400 210.450 802.540 220.000 ;
        RECT 710.340 210.130 710.600 210.450 ;
        RECT 802.340 210.130 802.600 210.450 ;
        RECT 710.400 2.400 710.540 210.130 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1478.510 207.300 1478.830 207.360 ;
        RECT 1482.650 207.300 1482.970 207.360 ;
        RECT 1478.510 207.160 1482.970 207.300 ;
        RECT 1478.510 207.100 1478.830 207.160 ;
        RECT 1482.650 207.100 1482.970 207.160 ;
        RECT 1482.650 16.900 1482.970 16.960 ;
        RECT 1530.950 16.900 1531.270 16.960 ;
        RECT 1482.650 16.760 1531.270 16.900 ;
        RECT 1482.650 16.700 1482.970 16.760 ;
        RECT 1530.950 16.700 1531.270 16.760 ;
      LAYER via ;
        RECT 1478.540 207.100 1478.800 207.360 ;
        RECT 1482.680 207.100 1482.940 207.360 ;
        RECT 1482.680 16.700 1482.940 16.960 ;
        RECT 1530.980 16.700 1531.240 16.960 ;
      LAYER met2 ;
        RECT 1478.580 220.000 1478.860 224.000 ;
        RECT 1478.600 207.390 1478.740 220.000 ;
        RECT 1478.540 207.070 1478.800 207.390 ;
        RECT 1482.680 207.070 1482.940 207.390 ;
        RECT 1482.740 16.990 1482.880 207.070 ;
        RECT 1482.680 16.670 1482.940 16.990 ;
        RECT 1530.980 16.670 1531.240 16.990 ;
        RECT 1531.040 2.400 1531.180 16.670 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1493.230 207.300 1493.550 207.360 ;
        RECT 1496.910 207.300 1497.230 207.360 ;
        RECT 1493.230 207.160 1497.230 207.300 ;
        RECT 1493.230 207.100 1493.550 207.160 ;
        RECT 1496.910 207.100 1497.230 207.160 ;
        RECT 1496.910 17.580 1497.230 17.640 ;
        RECT 1548.890 17.580 1549.210 17.640 ;
        RECT 1496.910 17.440 1549.210 17.580 ;
        RECT 1496.910 17.380 1497.230 17.440 ;
        RECT 1548.890 17.380 1549.210 17.440 ;
      LAYER via ;
        RECT 1493.260 207.100 1493.520 207.360 ;
        RECT 1496.940 207.100 1497.200 207.360 ;
        RECT 1496.940 17.380 1497.200 17.640 ;
        RECT 1548.920 17.380 1549.180 17.640 ;
      LAYER met2 ;
        RECT 1493.300 220.000 1493.580 224.000 ;
        RECT 1493.320 207.390 1493.460 220.000 ;
        RECT 1493.260 207.070 1493.520 207.390 ;
        RECT 1496.940 207.070 1497.200 207.390 ;
        RECT 1497.000 17.670 1497.140 207.070 ;
        RECT 1496.940 17.350 1497.200 17.670 ;
        RECT 1548.920 17.350 1549.180 17.670 ;
        RECT 1548.980 2.400 1549.120 17.350 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1510.710 18.940 1511.030 19.000 ;
        RECT 1566.830 18.940 1567.150 19.000 ;
        RECT 1510.710 18.800 1567.150 18.940 ;
        RECT 1510.710 18.740 1511.030 18.800 ;
        RECT 1566.830 18.740 1567.150 18.800 ;
      LAYER via ;
        RECT 1510.740 18.740 1511.000 19.000 ;
        RECT 1566.860 18.740 1567.120 19.000 ;
      LAYER met2 ;
        RECT 1508.020 220.730 1508.300 224.000 ;
        RECT 1508.020 220.590 1510.940 220.730 ;
        RECT 1508.020 220.000 1508.300 220.590 ;
        RECT 1510.800 19.030 1510.940 220.590 ;
        RECT 1510.740 18.710 1511.000 19.030 ;
        RECT 1566.860 18.710 1567.120 19.030 ;
        RECT 1566.920 2.400 1567.060 18.710 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1524.510 16.560 1524.830 16.620 ;
        RECT 1584.770 16.560 1585.090 16.620 ;
        RECT 1524.510 16.420 1585.090 16.560 ;
        RECT 1524.510 16.360 1524.830 16.420 ;
        RECT 1584.770 16.360 1585.090 16.420 ;
      LAYER via ;
        RECT 1524.540 16.360 1524.800 16.620 ;
        RECT 1584.800 16.360 1585.060 16.620 ;
      LAYER met2 ;
        RECT 1522.740 220.730 1523.020 224.000 ;
        RECT 1522.740 220.590 1524.740 220.730 ;
        RECT 1522.740 220.000 1523.020 220.590 ;
        RECT 1524.600 16.650 1524.740 220.590 ;
        RECT 1524.540 16.330 1524.800 16.650 ;
        RECT 1584.800 16.330 1585.060 16.650 ;
        RECT 1584.860 2.400 1585.000 16.330 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1538.310 17.240 1538.630 17.300 ;
        RECT 1602.250 17.240 1602.570 17.300 ;
        RECT 1538.310 17.100 1602.570 17.240 ;
        RECT 1538.310 17.040 1538.630 17.100 ;
        RECT 1602.250 17.040 1602.570 17.100 ;
      LAYER via ;
        RECT 1538.340 17.040 1538.600 17.300 ;
        RECT 1602.280 17.040 1602.540 17.300 ;
      LAYER met2 ;
        RECT 1537.460 220.730 1537.740 224.000 ;
        RECT 1537.460 220.590 1538.540 220.730 ;
        RECT 1537.460 220.000 1537.740 220.590 ;
        RECT 1538.400 17.330 1538.540 220.590 ;
        RECT 1538.340 17.010 1538.600 17.330 ;
        RECT 1602.280 17.010 1602.540 17.330 ;
        RECT 1602.340 2.400 1602.480 17.010 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1552.110 17.580 1552.430 17.640 ;
        RECT 1620.190 17.580 1620.510 17.640 ;
        RECT 1552.110 17.440 1620.510 17.580 ;
        RECT 1552.110 17.380 1552.430 17.440 ;
        RECT 1620.190 17.380 1620.510 17.440 ;
      LAYER via ;
        RECT 1552.140 17.380 1552.400 17.640 ;
        RECT 1620.220 17.380 1620.480 17.640 ;
      LAYER met2 ;
        RECT 1551.720 220.730 1552.000 224.000 ;
        RECT 1551.720 220.590 1552.340 220.730 ;
        RECT 1551.720 220.000 1552.000 220.590 ;
        RECT 1552.200 17.670 1552.340 220.590 ;
        RECT 1552.140 17.350 1552.400 17.670 ;
        RECT 1620.220 17.350 1620.480 17.670 ;
        RECT 1620.280 2.400 1620.420 17.350 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1566.370 207.300 1566.690 207.360 ;
        RECT 1572.810 207.300 1573.130 207.360 ;
        RECT 1566.370 207.160 1573.130 207.300 ;
        RECT 1566.370 207.100 1566.690 207.160 ;
        RECT 1572.810 207.100 1573.130 207.160 ;
        RECT 1572.810 20.640 1573.130 20.700 ;
        RECT 1638.130 20.640 1638.450 20.700 ;
        RECT 1572.810 20.500 1638.450 20.640 ;
        RECT 1572.810 20.440 1573.130 20.500 ;
        RECT 1638.130 20.440 1638.450 20.500 ;
      LAYER via ;
        RECT 1566.400 207.100 1566.660 207.360 ;
        RECT 1572.840 207.100 1573.100 207.360 ;
        RECT 1572.840 20.440 1573.100 20.700 ;
        RECT 1638.160 20.440 1638.420 20.700 ;
      LAYER met2 ;
        RECT 1566.440 220.000 1566.720 224.000 ;
        RECT 1566.460 207.390 1566.600 220.000 ;
        RECT 1566.400 207.070 1566.660 207.390 ;
        RECT 1572.840 207.070 1573.100 207.390 ;
        RECT 1572.900 20.730 1573.040 207.070 ;
        RECT 1572.840 20.410 1573.100 20.730 ;
        RECT 1638.160 20.410 1638.420 20.730 ;
        RECT 1638.220 2.400 1638.360 20.410 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1581.090 207.300 1581.410 207.360 ;
        RECT 1586.150 207.300 1586.470 207.360 ;
        RECT 1581.090 207.160 1586.470 207.300 ;
        RECT 1581.090 207.100 1581.410 207.160 ;
        RECT 1586.150 207.100 1586.470 207.160 ;
        RECT 1586.150 18.600 1586.470 18.660 ;
        RECT 1656.070 18.600 1656.390 18.660 ;
        RECT 1586.150 18.460 1656.390 18.600 ;
        RECT 1586.150 18.400 1586.470 18.460 ;
        RECT 1656.070 18.400 1656.390 18.460 ;
      LAYER via ;
        RECT 1581.120 207.100 1581.380 207.360 ;
        RECT 1586.180 207.100 1586.440 207.360 ;
        RECT 1586.180 18.400 1586.440 18.660 ;
        RECT 1656.100 18.400 1656.360 18.660 ;
      LAYER met2 ;
        RECT 1581.160 220.000 1581.440 224.000 ;
        RECT 1581.180 207.390 1581.320 220.000 ;
        RECT 1581.120 207.070 1581.380 207.390 ;
        RECT 1586.180 207.070 1586.440 207.390 ;
        RECT 1586.240 18.690 1586.380 207.070 ;
        RECT 1586.180 18.370 1586.440 18.690 ;
        RECT 1656.100 18.370 1656.360 18.690 ;
        RECT 1656.160 2.400 1656.300 18.370 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1595.810 207.300 1596.130 207.360 ;
        RECT 1600.410 207.300 1600.730 207.360 ;
        RECT 1595.810 207.160 1600.730 207.300 ;
        RECT 1595.810 207.100 1596.130 207.160 ;
        RECT 1600.410 207.100 1600.730 207.160 ;
        RECT 1600.410 15.540 1600.730 15.600 ;
        RECT 1673.550 15.540 1673.870 15.600 ;
        RECT 1600.410 15.400 1673.870 15.540 ;
        RECT 1600.410 15.340 1600.730 15.400 ;
        RECT 1673.550 15.340 1673.870 15.400 ;
      LAYER via ;
        RECT 1595.840 207.100 1596.100 207.360 ;
        RECT 1600.440 207.100 1600.700 207.360 ;
        RECT 1600.440 15.340 1600.700 15.600 ;
        RECT 1673.580 15.340 1673.840 15.600 ;
      LAYER met2 ;
        RECT 1595.880 220.000 1596.160 224.000 ;
        RECT 1595.900 207.390 1596.040 220.000 ;
        RECT 1595.840 207.070 1596.100 207.390 ;
        RECT 1600.440 207.070 1600.700 207.390 ;
        RECT 1600.500 15.630 1600.640 207.070 ;
        RECT 1600.440 15.310 1600.700 15.630 ;
        RECT 1673.580 15.310 1673.840 15.630 ;
        RECT 1673.640 2.400 1673.780 15.310 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1614.210 17.920 1614.530 17.980 ;
        RECT 1691.490 17.920 1691.810 17.980 ;
        RECT 1614.210 17.780 1691.810 17.920 ;
        RECT 1614.210 17.720 1614.530 17.780 ;
        RECT 1691.490 17.720 1691.810 17.780 ;
      LAYER via ;
        RECT 1614.240 17.720 1614.500 17.980 ;
        RECT 1691.520 17.720 1691.780 17.980 ;
      LAYER met2 ;
        RECT 1610.600 220.730 1610.880 224.000 ;
        RECT 1610.600 220.590 1614.440 220.730 ;
        RECT 1610.600 220.000 1610.880 220.590 ;
        RECT 1614.300 18.010 1614.440 220.590 ;
        RECT 1614.240 17.690 1614.500 18.010 ;
        RECT 1691.520 17.690 1691.780 18.010 ;
        RECT 1691.580 2.400 1691.720 17.690 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 731.010 211.380 731.330 211.440 ;
        RECT 817.030 211.380 817.350 211.440 ;
        RECT 731.010 211.240 817.350 211.380 ;
        RECT 731.010 211.180 731.330 211.240 ;
        RECT 817.030 211.180 817.350 211.240 ;
        RECT 728.250 17.580 728.570 17.640 ;
        RECT 731.010 17.580 731.330 17.640 ;
        RECT 728.250 17.440 731.330 17.580 ;
        RECT 728.250 17.380 728.570 17.440 ;
        RECT 731.010 17.380 731.330 17.440 ;
      LAYER via ;
        RECT 731.040 211.180 731.300 211.440 ;
        RECT 817.060 211.180 817.320 211.440 ;
        RECT 728.280 17.380 728.540 17.640 ;
        RECT 731.040 17.380 731.300 17.640 ;
      LAYER met2 ;
        RECT 817.100 220.000 817.380 224.000 ;
        RECT 817.120 211.470 817.260 220.000 ;
        RECT 731.040 211.150 731.300 211.470 ;
        RECT 817.060 211.150 817.320 211.470 ;
        RECT 731.100 17.670 731.240 211.150 ;
        RECT 728.280 17.350 728.540 17.670 ;
        RECT 731.040 17.350 731.300 17.670 ;
        RECT 728.340 2.400 728.480 17.350 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1628.010 20.300 1628.330 20.360 ;
        RECT 1709.430 20.300 1709.750 20.360 ;
        RECT 1628.010 20.160 1709.750 20.300 ;
        RECT 1628.010 20.100 1628.330 20.160 ;
        RECT 1709.430 20.100 1709.750 20.160 ;
      LAYER via ;
        RECT 1628.040 20.100 1628.300 20.360 ;
        RECT 1709.460 20.100 1709.720 20.360 ;
      LAYER met2 ;
        RECT 1625.320 220.730 1625.600 224.000 ;
        RECT 1625.320 220.590 1628.240 220.730 ;
        RECT 1625.320 220.000 1625.600 220.590 ;
        RECT 1628.100 20.390 1628.240 220.590 ;
        RECT 1628.040 20.070 1628.300 20.390 ;
        RECT 1709.460 20.070 1709.720 20.390 ;
        RECT 1709.520 2.400 1709.660 20.070 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1641.810 20.640 1642.130 20.700 ;
        RECT 1727.370 20.640 1727.690 20.700 ;
        RECT 1641.810 20.500 1727.690 20.640 ;
        RECT 1641.810 20.440 1642.130 20.500 ;
        RECT 1727.370 20.440 1727.690 20.500 ;
      LAYER via ;
        RECT 1641.840 20.440 1642.100 20.700 ;
        RECT 1727.400 20.440 1727.660 20.700 ;
      LAYER met2 ;
        RECT 1640.040 220.730 1640.320 224.000 ;
        RECT 1640.040 220.590 1642.040 220.730 ;
        RECT 1640.040 220.000 1640.320 220.590 ;
        RECT 1641.900 20.730 1642.040 220.590 ;
        RECT 1641.840 20.410 1642.100 20.730 ;
        RECT 1727.400 20.410 1727.660 20.730 ;
        RECT 1727.460 2.400 1727.600 20.410 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1655.610 14.860 1655.930 14.920 ;
        RECT 1745.310 14.860 1745.630 14.920 ;
        RECT 1655.610 14.720 1745.630 14.860 ;
        RECT 1655.610 14.660 1655.930 14.720 ;
        RECT 1745.310 14.660 1745.630 14.720 ;
      LAYER via ;
        RECT 1655.640 14.660 1655.900 14.920 ;
        RECT 1745.340 14.660 1745.600 14.920 ;
      LAYER met2 ;
        RECT 1654.760 220.730 1655.040 224.000 ;
        RECT 1654.760 220.590 1655.840 220.730 ;
        RECT 1654.760 220.000 1655.040 220.590 ;
        RECT 1655.700 14.950 1655.840 220.590 ;
        RECT 1655.640 14.630 1655.900 14.950 ;
        RECT 1745.340 14.630 1745.600 14.950 ;
        RECT 1745.400 2.400 1745.540 14.630 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1669.410 18.600 1669.730 18.660 ;
        RECT 1762.790 18.600 1763.110 18.660 ;
        RECT 1669.410 18.460 1763.110 18.600 ;
        RECT 1669.410 18.400 1669.730 18.460 ;
        RECT 1762.790 18.400 1763.110 18.460 ;
      LAYER via ;
        RECT 1669.440 18.400 1669.700 18.660 ;
        RECT 1762.820 18.400 1763.080 18.660 ;
      LAYER met2 ;
        RECT 1669.480 220.000 1669.760 224.000 ;
        RECT 1669.500 18.690 1669.640 220.000 ;
        RECT 1669.440 18.370 1669.700 18.690 ;
        RECT 1762.820 18.370 1763.080 18.690 ;
        RECT 1762.880 2.400 1763.020 18.370 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1684.130 207.300 1684.450 207.360 ;
        RECT 1690.110 207.300 1690.430 207.360 ;
        RECT 1684.130 207.160 1690.430 207.300 ;
        RECT 1684.130 207.100 1684.450 207.160 ;
        RECT 1690.110 207.100 1690.430 207.160 ;
        RECT 1690.110 15.880 1690.430 15.940 ;
        RECT 1780.730 15.880 1781.050 15.940 ;
        RECT 1690.110 15.740 1781.050 15.880 ;
        RECT 1690.110 15.680 1690.430 15.740 ;
        RECT 1780.730 15.680 1781.050 15.740 ;
      LAYER via ;
        RECT 1684.160 207.100 1684.420 207.360 ;
        RECT 1690.140 207.100 1690.400 207.360 ;
        RECT 1690.140 15.680 1690.400 15.940 ;
        RECT 1780.760 15.680 1781.020 15.940 ;
      LAYER met2 ;
        RECT 1684.200 220.000 1684.480 224.000 ;
        RECT 1684.220 207.390 1684.360 220.000 ;
        RECT 1684.160 207.070 1684.420 207.390 ;
        RECT 1690.140 207.070 1690.400 207.390 ;
        RECT 1690.200 15.970 1690.340 207.070 ;
        RECT 1690.140 15.650 1690.400 15.970 ;
        RECT 1780.760 15.650 1781.020 15.970 ;
        RECT 1780.820 2.400 1780.960 15.650 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1698.850 207.300 1699.170 207.360 ;
        RECT 1703.910 207.300 1704.230 207.360 ;
        RECT 1698.850 207.160 1704.230 207.300 ;
        RECT 1698.850 207.100 1699.170 207.160 ;
        RECT 1703.910 207.100 1704.230 207.160 ;
        RECT 1702.530 26.760 1702.850 26.820 ;
        RECT 1703.910 26.760 1704.230 26.820 ;
        RECT 1702.530 26.620 1704.230 26.760 ;
        RECT 1702.530 26.560 1702.850 26.620 ;
        RECT 1703.910 26.560 1704.230 26.620 ;
        RECT 1702.530 15.540 1702.850 15.600 ;
        RECT 1798.670 15.540 1798.990 15.600 ;
        RECT 1702.530 15.400 1798.990 15.540 ;
        RECT 1702.530 15.340 1702.850 15.400 ;
        RECT 1798.670 15.340 1798.990 15.400 ;
      LAYER via ;
        RECT 1698.880 207.100 1699.140 207.360 ;
        RECT 1703.940 207.100 1704.200 207.360 ;
        RECT 1702.560 26.560 1702.820 26.820 ;
        RECT 1703.940 26.560 1704.200 26.820 ;
        RECT 1702.560 15.340 1702.820 15.600 ;
        RECT 1798.700 15.340 1798.960 15.600 ;
      LAYER met2 ;
        RECT 1698.920 220.000 1699.200 224.000 ;
        RECT 1698.940 207.390 1699.080 220.000 ;
        RECT 1698.880 207.070 1699.140 207.390 ;
        RECT 1703.940 207.070 1704.200 207.390 ;
        RECT 1704.000 26.850 1704.140 207.070 ;
        RECT 1702.560 26.530 1702.820 26.850 ;
        RECT 1703.940 26.530 1704.200 26.850 ;
        RECT 1702.620 15.630 1702.760 26.530 ;
        RECT 1702.560 15.310 1702.820 15.630 ;
        RECT 1798.700 15.310 1798.960 15.630 ;
        RECT 1798.760 2.400 1798.900 15.310 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1713.570 207.300 1713.890 207.360 ;
        RECT 1717.710 207.300 1718.030 207.360 ;
        RECT 1713.570 207.160 1718.030 207.300 ;
        RECT 1713.570 207.100 1713.890 207.160 ;
        RECT 1717.710 207.100 1718.030 207.160 ;
        RECT 1717.710 18.260 1718.030 18.320 ;
        RECT 1816.610 18.260 1816.930 18.320 ;
        RECT 1717.710 18.120 1816.930 18.260 ;
        RECT 1717.710 18.060 1718.030 18.120 ;
        RECT 1816.610 18.060 1816.930 18.120 ;
      LAYER via ;
        RECT 1713.600 207.100 1713.860 207.360 ;
        RECT 1717.740 207.100 1718.000 207.360 ;
        RECT 1717.740 18.060 1718.000 18.320 ;
        RECT 1816.640 18.060 1816.900 18.320 ;
      LAYER met2 ;
        RECT 1713.640 220.000 1713.920 224.000 ;
        RECT 1713.660 207.390 1713.800 220.000 ;
        RECT 1713.600 207.070 1713.860 207.390 ;
        RECT 1717.740 207.070 1718.000 207.390 ;
        RECT 1717.800 18.350 1717.940 207.070 ;
        RECT 1717.740 18.030 1718.000 18.350 ;
        RECT 1816.640 18.030 1816.900 18.350 ;
        RECT 1816.700 2.400 1816.840 18.030 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1731.510 20.640 1731.830 20.700 ;
        RECT 1834.550 20.640 1834.870 20.700 ;
        RECT 1731.510 20.500 1834.870 20.640 ;
        RECT 1731.510 20.440 1731.830 20.500 ;
        RECT 1834.550 20.440 1834.870 20.500 ;
      LAYER via ;
        RECT 1731.540 20.440 1731.800 20.700 ;
        RECT 1834.580 20.440 1834.840 20.700 ;
      LAYER met2 ;
        RECT 1728.360 220.730 1728.640 224.000 ;
        RECT 1728.360 220.590 1731.740 220.730 ;
        RECT 1728.360 220.000 1728.640 220.590 ;
        RECT 1731.600 20.730 1731.740 220.590 ;
        RECT 1731.540 20.410 1731.800 20.730 ;
        RECT 1834.580 20.410 1834.840 20.730 ;
        RECT 1834.640 2.400 1834.780 20.410 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1745.310 19.620 1745.630 19.680 ;
        RECT 1852.030 19.620 1852.350 19.680 ;
        RECT 1745.310 19.480 1852.350 19.620 ;
        RECT 1745.310 19.420 1745.630 19.480 ;
        RECT 1852.030 19.420 1852.350 19.480 ;
      LAYER via ;
        RECT 1745.340 19.420 1745.600 19.680 ;
        RECT 1852.060 19.420 1852.320 19.680 ;
      LAYER met2 ;
        RECT 1743.080 220.730 1743.360 224.000 ;
        RECT 1743.080 220.590 1745.540 220.730 ;
        RECT 1743.080 220.000 1743.360 220.590 ;
        RECT 1745.400 19.710 1745.540 220.590 ;
        RECT 1745.340 19.390 1745.600 19.710 ;
        RECT 1852.060 19.390 1852.320 19.710 ;
        RECT 1852.120 2.400 1852.260 19.390 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1759.110 16.560 1759.430 16.620 ;
        RECT 1869.970 16.560 1870.290 16.620 ;
        RECT 1759.110 16.420 1870.290 16.560 ;
        RECT 1759.110 16.360 1759.430 16.420 ;
        RECT 1869.970 16.360 1870.290 16.420 ;
      LAYER via ;
        RECT 1759.140 16.360 1759.400 16.620 ;
        RECT 1870.000 16.360 1870.260 16.620 ;
      LAYER met2 ;
        RECT 1757.800 220.730 1758.080 224.000 ;
        RECT 1757.800 220.590 1759.340 220.730 ;
        RECT 1757.800 220.000 1758.080 220.590 ;
        RECT 1759.200 16.650 1759.340 220.590 ;
        RECT 1759.140 16.330 1759.400 16.650 ;
        RECT 1870.000 16.330 1870.260 16.650 ;
        RECT 1870.060 2.400 1870.200 16.330 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 751.710 207.980 752.030 208.040 ;
        RECT 831.750 207.980 832.070 208.040 ;
        RECT 751.710 207.840 832.070 207.980 ;
        RECT 751.710 207.780 752.030 207.840 ;
        RECT 831.750 207.780 832.070 207.840 ;
        RECT 746.190 17.580 746.510 17.640 ;
        RECT 751.710 17.580 752.030 17.640 ;
        RECT 746.190 17.440 752.030 17.580 ;
        RECT 746.190 17.380 746.510 17.440 ;
        RECT 751.710 17.380 752.030 17.440 ;
      LAYER via ;
        RECT 751.740 207.780 752.000 208.040 ;
        RECT 831.780 207.780 832.040 208.040 ;
        RECT 746.220 17.380 746.480 17.640 ;
        RECT 751.740 17.380 752.000 17.640 ;
      LAYER met2 ;
        RECT 831.820 220.000 832.100 224.000 ;
        RECT 831.840 208.070 831.980 220.000 ;
        RECT 751.740 207.750 752.000 208.070 ;
        RECT 831.780 207.750 832.040 208.070 ;
        RECT 751.800 17.670 751.940 207.750 ;
        RECT 746.220 17.350 746.480 17.670 ;
        RECT 751.740 17.350 752.000 17.670 ;
        RECT 746.280 2.400 746.420 17.350 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.910 18.940 1773.230 19.000 ;
        RECT 1887.910 18.940 1888.230 19.000 ;
        RECT 1772.910 18.800 1888.230 18.940 ;
        RECT 1772.910 18.740 1773.230 18.800 ;
        RECT 1887.910 18.740 1888.230 18.800 ;
      LAYER via ;
        RECT 1772.940 18.740 1773.200 19.000 ;
        RECT 1887.940 18.740 1888.200 19.000 ;
      LAYER met2 ;
        RECT 1772.520 220.730 1772.800 224.000 ;
        RECT 1772.520 220.590 1773.140 220.730 ;
        RECT 1772.520 220.000 1772.800 220.590 ;
        RECT 1773.000 19.030 1773.140 220.590 ;
        RECT 1772.940 18.710 1773.200 19.030 ;
        RECT 1887.940 18.710 1888.200 19.030 ;
        RECT 1888.000 2.400 1888.140 18.710 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1787.170 207.300 1787.490 207.360 ;
        RECT 1793.610 207.300 1793.930 207.360 ;
        RECT 1787.170 207.160 1793.930 207.300 ;
        RECT 1787.170 207.100 1787.490 207.160 ;
        RECT 1793.610 207.100 1793.930 207.160 ;
        RECT 1793.610 18.600 1793.930 18.660 ;
        RECT 1905.850 18.600 1906.170 18.660 ;
        RECT 1793.610 18.460 1906.170 18.600 ;
        RECT 1793.610 18.400 1793.930 18.460 ;
        RECT 1905.850 18.400 1906.170 18.460 ;
      LAYER via ;
        RECT 1787.200 207.100 1787.460 207.360 ;
        RECT 1793.640 207.100 1793.900 207.360 ;
        RECT 1793.640 18.400 1793.900 18.660 ;
        RECT 1905.880 18.400 1906.140 18.660 ;
      LAYER met2 ;
        RECT 1787.240 220.000 1787.520 224.000 ;
        RECT 1787.260 207.390 1787.400 220.000 ;
        RECT 1787.200 207.070 1787.460 207.390 ;
        RECT 1793.640 207.070 1793.900 207.390 ;
        RECT 1793.700 18.690 1793.840 207.070 ;
        RECT 1793.640 18.370 1793.900 18.690 ;
        RECT 1905.880 18.370 1906.140 18.690 ;
        RECT 1905.940 2.400 1906.080 18.370 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1801.430 207.300 1801.750 207.360 ;
        RECT 1807.410 207.300 1807.730 207.360 ;
        RECT 1801.430 207.160 1807.730 207.300 ;
        RECT 1801.430 207.100 1801.750 207.160 ;
        RECT 1807.410 207.100 1807.730 207.160 ;
        RECT 1807.410 15.540 1807.730 15.600 ;
        RECT 1923.330 15.540 1923.650 15.600 ;
        RECT 1807.410 15.400 1923.650 15.540 ;
        RECT 1807.410 15.340 1807.730 15.400 ;
        RECT 1923.330 15.340 1923.650 15.400 ;
      LAYER via ;
        RECT 1801.460 207.100 1801.720 207.360 ;
        RECT 1807.440 207.100 1807.700 207.360 ;
        RECT 1807.440 15.340 1807.700 15.600 ;
        RECT 1923.360 15.340 1923.620 15.600 ;
      LAYER met2 ;
        RECT 1801.500 220.000 1801.780 224.000 ;
        RECT 1801.520 207.390 1801.660 220.000 ;
        RECT 1801.460 207.070 1801.720 207.390 ;
        RECT 1807.440 207.070 1807.700 207.390 ;
        RECT 1807.500 15.630 1807.640 207.070 ;
        RECT 1807.440 15.310 1807.700 15.630 ;
        RECT 1923.360 15.310 1923.620 15.630 ;
        RECT 1923.420 2.400 1923.560 15.310 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1816.150 207.300 1816.470 207.360 ;
        RECT 1821.210 207.300 1821.530 207.360 ;
        RECT 1816.150 207.160 1821.530 207.300 ;
        RECT 1816.150 207.100 1816.470 207.160 ;
        RECT 1821.210 207.100 1821.530 207.160 ;
        RECT 1821.210 18.260 1821.530 18.320 ;
        RECT 1941.270 18.260 1941.590 18.320 ;
        RECT 1821.210 18.120 1941.590 18.260 ;
        RECT 1821.210 18.060 1821.530 18.120 ;
        RECT 1941.270 18.060 1941.590 18.120 ;
      LAYER via ;
        RECT 1816.180 207.100 1816.440 207.360 ;
        RECT 1821.240 207.100 1821.500 207.360 ;
        RECT 1821.240 18.060 1821.500 18.320 ;
        RECT 1941.300 18.060 1941.560 18.320 ;
      LAYER met2 ;
        RECT 1816.220 220.000 1816.500 224.000 ;
        RECT 1816.240 207.390 1816.380 220.000 ;
        RECT 1816.180 207.070 1816.440 207.390 ;
        RECT 1821.240 207.070 1821.500 207.390 ;
        RECT 1821.300 18.350 1821.440 207.070 ;
        RECT 1821.240 18.030 1821.500 18.350 ;
        RECT 1941.300 18.030 1941.560 18.350 ;
        RECT 1941.360 2.400 1941.500 18.030 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1830.870 207.300 1831.190 207.360 ;
        RECT 1835.010 207.300 1835.330 207.360 ;
        RECT 1830.870 207.160 1835.330 207.300 ;
        RECT 1830.870 207.100 1831.190 207.160 ;
        RECT 1835.010 207.100 1835.330 207.160 ;
        RECT 1835.010 15.880 1835.330 15.940 ;
        RECT 1959.210 15.880 1959.530 15.940 ;
        RECT 1835.010 15.740 1959.530 15.880 ;
        RECT 1835.010 15.680 1835.330 15.740 ;
        RECT 1959.210 15.680 1959.530 15.740 ;
      LAYER via ;
        RECT 1830.900 207.100 1831.160 207.360 ;
        RECT 1835.040 207.100 1835.300 207.360 ;
        RECT 1835.040 15.680 1835.300 15.940 ;
        RECT 1959.240 15.680 1959.500 15.940 ;
      LAYER met2 ;
        RECT 1830.940 220.000 1831.220 224.000 ;
        RECT 1830.960 207.390 1831.100 220.000 ;
        RECT 1830.900 207.070 1831.160 207.390 ;
        RECT 1835.040 207.070 1835.300 207.390 ;
        RECT 1835.100 15.970 1835.240 207.070 ;
        RECT 1835.040 15.650 1835.300 15.970 ;
        RECT 1959.240 15.650 1959.500 15.970 ;
        RECT 1959.300 2.400 1959.440 15.650 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1848.810 16.900 1849.130 16.960 ;
        RECT 1977.150 16.900 1977.470 16.960 ;
        RECT 1848.810 16.760 1977.470 16.900 ;
        RECT 1848.810 16.700 1849.130 16.760 ;
        RECT 1977.150 16.700 1977.470 16.760 ;
      LAYER via ;
        RECT 1848.840 16.700 1849.100 16.960 ;
        RECT 1977.180 16.700 1977.440 16.960 ;
      LAYER met2 ;
        RECT 1845.660 220.730 1845.940 224.000 ;
        RECT 1845.660 220.590 1849.040 220.730 ;
        RECT 1845.660 220.000 1845.940 220.590 ;
        RECT 1848.900 16.990 1849.040 220.590 ;
        RECT 1848.840 16.670 1849.100 16.990 ;
        RECT 1977.180 16.670 1977.440 16.990 ;
        RECT 1977.240 2.400 1977.380 16.670 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1862.610 19.620 1862.930 19.680 ;
        RECT 1995.090 19.620 1995.410 19.680 ;
        RECT 1862.610 19.480 1995.410 19.620 ;
        RECT 1862.610 19.420 1862.930 19.480 ;
        RECT 1995.090 19.420 1995.410 19.480 ;
      LAYER via ;
        RECT 1862.640 19.420 1862.900 19.680 ;
        RECT 1995.120 19.420 1995.380 19.680 ;
      LAYER met2 ;
        RECT 1860.380 220.730 1860.660 224.000 ;
        RECT 1860.380 220.590 1862.840 220.730 ;
        RECT 1860.380 220.000 1860.660 220.590 ;
        RECT 1862.700 19.710 1862.840 220.590 ;
        RECT 1862.640 19.390 1862.900 19.710 ;
        RECT 1995.120 19.390 1995.380 19.710 ;
        RECT 1995.180 2.400 1995.320 19.390 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1876.410 16.560 1876.730 16.620 ;
        RECT 2012.570 16.560 2012.890 16.620 ;
        RECT 1876.410 16.420 2012.890 16.560 ;
        RECT 1876.410 16.360 1876.730 16.420 ;
        RECT 2012.570 16.360 2012.890 16.420 ;
      LAYER via ;
        RECT 1876.440 16.360 1876.700 16.620 ;
        RECT 2012.600 16.360 2012.860 16.620 ;
      LAYER met2 ;
        RECT 1875.100 220.730 1875.380 224.000 ;
        RECT 1875.100 220.590 1876.640 220.730 ;
        RECT 1875.100 220.000 1875.380 220.590 ;
        RECT 1876.500 16.650 1876.640 220.590 ;
        RECT 1876.440 16.330 1876.700 16.650 ;
        RECT 2012.600 16.330 2012.860 16.650 ;
        RECT 2012.660 2.400 2012.800 16.330 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1890.210 18.940 1890.530 19.000 ;
        RECT 2030.510 18.940 2030.830 19.000 ;
        RECT 1890.210 18.800 2030.830 18.940 ;
        RECT 1890.210 18.740 1890.530 18.800 ;
        RECT 2030.510 18.740 2030.830 18.800 ;
      LAYER via ;
        RECT 1890.240 18.740 1890.500 19.000 ;
        RECT 2030.540 18.740 2030.800 19.000 ;
      LAYER met2 ;
        RECT 1889.820 220.730 1890.100 224.000 ;
        RECT 1889.820 220.590 1890.440 220.730 ;
        RECT 1889.820 220.000 1890.100 220.590 ;
        RECT 1890.300 19.030 1890.440 220.590 ;
        RECT 1890.240 18.710 1890.500 19.030 ;
        RECT 2030.540 18.710 2030.800 19.030 ;
        RECT 2030.600 2.400 2030.740 18.710 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1904.470 207.300 1904.790 207.360 ;
        RECT 1910.910 207.300 1911.230 207.360 ;
        RECT 1904.470 207.160 1911.230 207.300 ;
        RECT 1904.470 207.100 1904.790 207.160 ;
        RECT 1910.910 207.100 1911.230 207.160 ;
        RECT 1910.910 14.520 1911.230 14.580 ;
        RECT 2048.450 14.520 2048.770 14.580 ;
        RECT 1910.910 14.380 2048.770 14.520 ;
        RECT 1910.910 14.320 1911.230 14.380 ;
        RECT 2048.450 14.320 2048.770 14.380 ;
      LAYER via ;
        RECT 1904.500 207.100 1904.760 207.360 ;
        RECT 1910.940 207.100 1911.200 207.360 ;
        RECT 1910.940 14.320 1911.200 14.580 ;
        RECT 2048.480 14.320 2048.740 14.580 ;
      LAYER met2 ;
        RECT 1904.540 220.000 1904.820 224.000 ;
        RECT 1904.560 207.390 1904.700 220.000 ;
        RECT 1904.500 207.070 1904.760 207.390 ;
        RECT 1910.940 207.070 1911.200 207.390 ;
        RECT 1911.000 14.610 1911.140 207.070 ;
        RECT 1910.940 14.290 1911.200 14.610 ;
        RECT 2048.480 14.290 2048.740 14.610 ;
        RECT 2048.540 2.400 2048.680 14.290 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 765.510 210.020 765.830 210.080 ;
        RECT 846.470 210.020 846.790 210.080 ;
        RECT 765.510 209.880 846.790 210.020 ;
        RECT 765.510 209.820 765.830 209.880 ;
        RECT 846.470 209.820 846.790 209.880 ;
      LAYER via ;
        RECT 765.540 209.820 765.800 210.080 ;
        RECT 846.500 209.820 846.760 210.080 ;
      LAYER met2 ;
        RECT 846.540 220.000 846.820 224.000 ;
        RECT 846.560 210.110 846.700 220.000 ;
        RECT 765.540 209.790 765.800 210.110 ;
        RECT 846.500 209.790 846.760 210.110 ;
        RECT 765.600 17.410 765.740 209.790 ;
        RECT 763.760 17.270 765.740 17.410 ;
        RECT 763.760 2.400 763.900 17.270 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1919.190 207.300 1919.510 207.360 ;
        RECT 1924.710 207.300 1925.030 207.360 ;
        RECT 1919.190 207.160 1925.030 207.300 ;
        RECT 1919.190 207.100 1919.510 207.160 ;
        RECT 1924.710 207.100 1925.030 207.160 ;
        RECT 1924.710 14.860 1925.030 14.920 ;
        RECT 2066.390 14.860 2066.710 14.920 ;
        RECT 1924.710 14.720 2066.710 14.860 ;
        RECT 1924.710 14.660 1925.030 14.720 ;
        RECT 2066.390 14.660 2066.710 14.720 ;
      LAYER via ;
        RECT 1919.220 207.100 1919.480 207.360 ;
        RECT 1924.740 207.100 1925.000 207.360 ;
        RECT 1924.740 14.660 1925.000 14.920 ;
        RECT 2066.420 14.660 2066.680 14.920 ;
      LAYER met2 ;
        RECT 1919.260 220.000 1919.540 224.000 ;
        RECT 1919.280 207.390 1919.420 220.000 ;
        RECT 1919.220 207.070 1919.480 207.390 ;
        RECT 1924.740 207.070 1925.000 207.390 ;
        RECT 1924.800 14.950 1924.940 207.070 ;
        RECT 1924.740 14.630 1925.000 14.950 ;
        RECT 2066.420 14.630 2066.680 14.950 ;
        RECT 2066.480 2.400 2066.620 14.630 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1933.910 207.300 1934.230 207.360 ;
        RECT 1938.510 207.300 1938.830 207.360 ;
        RECT 1933.910 207.160 1938.830 207.300 ;
        RECT 1933.910 207.100 1934.230 207.160 ;
        RECT 1938.510 207.100 1938.830 207.160 ;
        RECT 1938.510 17.920 1938.830 17.980 ;
        RECT 2084.330 17.920 2084.650 17.980 ;
        RECT 1938.510 17.780 2084.650 17.920 ;
        RECT 1938.510 17.720 1938.830 17.780 ;
        RECT 2084.330 17.720 2084.650 17.780 ;
      LAYER via ;
        RECT 1933.940 207.100 1934.200 207.360 ;
        RECT 1938.540 207.100 1938.800 207.360 ;
        RECT 1938.540 17.720 1938.800 17.980 ;
        RECT 2084.360 17.720 2084.620 17.980 ;
      LAYER met2 ;
        RECT 1933.980 220.000 1934.260 224.000 ;
        RECT 1934.000 207.390 1934.140 220.000 ;
        RECT 1933.940 207.070 1934.200 207.390 ;
        RECT 1938.540 207.070 1938.800 207.390 ;
        RECT 1938.600 18.010 1938.740 207.070 ;
        RECT 1938.540 17.690 1938.800 18.010 ;
        RECT 2084.360 17.690 2084.620 18.010 ;
        RECT 2084.420 2.400 2084.560 17.690 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1948.630 207.300 1948.950 207.360 ;
        RECT 1952.310 207.300 1952.630 207.360 ;
        RECT 1948.630 207.160 1952.630 207.300 ;
        RECT 1948.630 207.100 1948.950 207.160 ;
        RECT 1952.310 207.100 1952.630 207.160 ;
        RECT 1952.310 18.260 1952.630 18.320 ;
        RECT 2101.810 18.260 2102.130 18.320 ;
        RECT 1952.310 18.120 2102.130 18.260 ;
        RECT 1952.310 18.060 1952.630 18.120 ;
        RECT 2101.810 18.060 2102.130 18.120 ;
      LAYER via ;
        RECT 1948.660 207.100 1948.920 207.360 ;
        RECT 1952.340 207.100 1952.600 207.360 ;
        RECT 1952.340 18.060 1952.600 18.320 ;
        RECT 2101.840 18.060 2102.100 18.320 ;
      LAYER met2 ;
        RECT 1948.700 220.000 1948.980 224.000 ;
        RECT 1948.720 207.390 1948.860 220.000 ;
        RECT 1948.660 207.070 1948.920 207.390 ;
        RECT 1952.340 207.070 1952.600 207.390 ;
        RECT 1952.400 18.350 1952.540 207.070 ;
        RECT 1952.340 18.030 1952.600 18.350 ;
        RECT 2101.840 18.030 2102.100 18.350 ;
        RECT 2101.900 2.400 2102.040 18.030 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1966.110 17.580 1966.430 17.640 ;
        RECT 2119.750 17.580 2120.070 17.640 ;
        RECT 1966.110 17.440 2120.070 17.580 ;
        RECT 1966.110 17.380 1966.430 17.440 ;
        RECT 2119.750 17.380 2120.070 17.440 ;
      LAYER via ;
        RECT 1966.140 17.380 1966.400 17.640 ;
        RECT 2119.780 17.380 2120.040 17.640 ;
      LAYER met2 ;
        RECT 1963.420 220.730 1963.700 224.000 ;
        RECT 1963.420 220.590 1966.340 220.730 ;
        RECT 1963.420 220.000 1963.700 220.590 ;
        RECT 1966.200 17.670 1966.340 220.590 ;
        RECT 1966.140 17.350 1966.400 17.670 ;
        RECT 2119.780 17.350 2120.040 17.670 ;
        RECT 2119.840 2.400 2119.980 17.350 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2007.125 16.745 2007.295 19.975 ;
      LAYER mcon ;
        RECT 2007.125 19.805 2007.295 19.975 ;
      LAYER met1 ;
        RECT 1979.910 19.960 1980.230 20.020 ;
        RECT 2007.065 19.960 2007.355 20.005 ;
        RECT 1979.910 19.820 2007.355 19.960 ;
        RECT 1979.910 19.760 1980.230 19.820 ;
        RECT 2007.065 19.775 2007.355 19.820 ;
        RECT 2007.065 16.900 2007.355 16.945 ;
        RECT 2137.690 16.900 2138.010 16.960 ;
        RECT 2007.065 16.760 2138.010 16.900 ;
        RECT 2007.065 16.715 2007.355 16.760 ;
        RECT 2137.690 16.700 2138.010 16.760 ;
      LAYER via ;
        RECT 1979.940 19.760 1980.200 20.020 ;
        RECT 2137.720 16.700 2137.980 16.960 ;
      LAYER met2 ;
        RECT 1978.140 220.730 1978.420 224.000 ;
        RECT 1978.140 220.590 1980.140 220.730 ;
        RECT 1978.140 220.000 1978.420 220.590 ;
        RECT 1980.000 20.050 1980.140 220.590 ;
        RECT 1979.940 19.730 1980.200 20.050 ;
        RECT 2137.720 16.670 2137.980 16.990 ;
        RECT 2137.780 2.400 2137.920 16.670 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1993.710 20.300 1994.030 20.360 ;
        RECT 2155.630 20.300 2155.950 20.360 ;
        RECT 1993.710 20.160 2155.950 20.300 ;
        RECT 1993.710 20.100 1994.030 20.160 ;
        RECT 2155.630 20.100 2155.950 20.160 ;
      LAYER via ;
        RECT 1993.740 20.100 1994.000 20.360 ;
        RECT 2155.660 20.100 2155.920 20.360 ;
      LAYER met2 ;
        RECT 1992.860 220.730 1993.140 224.000 ;
        RECT 1992.860 220.590 1993.940 220.730 ;
        RECT 1992.860 220.000 1993.140 220.590 ;
        RECT 1993.800 20.390 1993.940 220.590 ;
        RECT 1993.740 20.070 1994.000 20.390 ;
        RECT 2155.660 20.070 2155.920 20.390 ;
        RECT 2155.720 2.400 2155.860 20.070 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2115.225 18.785 2115.395 19.975 ;
        RECT 2156.165 16.745 2156.335 18.955 ;
      LAYER mcon ;
        RECT 2115.225 19.805 2115.395 19.975 ;
        RECT 2156.165 18.785 2156.335 18.955 ;
      LAYER met1 ;
        RECT 2007.510 19.960 2007.830 20.020 ;
        RECT 2115.165 19.960 2115.455 20.005 ;
        RECT 2007.510 19.820 2115.455 19.960 ;
        RECT 2007.510 19.760 2007.830 19.820 ;
        RECT 2115.165 19.775 2115.455 19.820 ;
        RECT 2115.165 18.940 2115.455 18.985 ;
        RECT 2156.105 18.940 2156.395 18.985 ;
        RECT 2115.165 18.800 2156.395 18.940 ;
        RECT 2115.165 18.755 2115.455 18.800 ;
        RECT 2156.105 18.755 2156.395 18.800 ;
        RECT 2156.105 16.900 2156.395 16.945 ;
        RECT 2173.110 16.900 2173.430 16.960 ;
        RECT 2156.105 16.760 2173.430 16.900 ;
        RECT 2156.105 16.715 2156.395 16.760 ;
        RECT 2173.110 16.700 2173.430 16.760 ;
      LAYER via ;
        RECT 2007.540 19.760 2007.800 20.020 ;
        RECT 2173.140 16.700 2173.400 16.960 ;
      LAYER met2 ;
        RECT 2007.580 220.000 2007.860 224.000 ;
        RECT 2007.600 20.050 2007.740 220.000 ;
        RECT 2007.540 19.730 2007.800 20.050 ;
        RECT 2173.140 16.670 2173.400 16.990 ;
        RECT 2173.200 2.400 2173.340 16.670 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2022.230 213.420 2022.550 213.480 ;
        RECT 2028.210 213.420 2028.530 213.480 ;
        RECT 2022.230 213.280 2028.530 213.420 ;
        RECT 2022.230 213.220 2022.550 213.280 ;
        RECT 2028.210 213.220 2028.530 213.280 ;
        RECT 2028.210 16.220 2028.530 16.280 ;
        RECT 2191.050 16.220 2191.370 16.280 ;
        RECT 2028.210 16.080 2191.370 16.220 ;
        RECT 2028.210 16.020 2028.530 16.080 ;
        RECT 2191.050 16.020 2191.370 16.080 ;
      LAYER via ;
        RECT 2022.260 213.220 2022.520 213.480 ;
        RECT 2028.240 213.220 2028.500 213.480 ;
        RECT 2028.240 16.020 2028.500 16.280 ;
        RECT 2191.080 16.020 2191.340 16.280 ;
      LAYER met2 ;
        RECT 2022.300 220.000 2022.580 224.000 ;
        RECT 2022.320 213.510 2022.460 220.000 ;
        RECT 2022.260 213.190 2022.520 213.510 ;
        RECT 2028.240 213.190 2028.500 213.510 ;
        RECT 2028.300 16.310 2028.440 213.190 ;
        RECT 2028.240 15.990 2028.500 16.310 ;
        RECT 2191.080 15.990 2191.340 16.310 ;
        RECT 2191.140 2.400 2191.280 15.990 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2114.305 15.725 2114.475 19.635 ;
        RECT 2163.065 15.725 2163.235 19.635 ;
      LAYER mcon ;
        RECT 2114.305 19.465 2114.475 19.635 ;
        RECT 2163.065 19.465 2163.235 19.635 ;
      LAYER met1 ;
        RECT 2036.950 211.040 2037.270 211.100 ;
        RECT 2042.010 211.040 2042.330 211.100 ;
        RECT 2036.950 210.900 2042.330 211.040 ;
        RECT 2036.950 210.840 2037.270 210.900 ;
        RECT 2042.010 210.840 2042.330 210.900 ;
        RECT 2114.245 19.620 2114.535 19.665 ;
        RECT 2055.440 19.480 2114.535 19.620 ;
        RECT 2042.010 18.940 2042.330 19.000 ;
        RECT 2055.440 18.940 2055.580 19.480 ;
        RECT 2114.245 19.435 2114.535 19.480 ;
        RECT 2163.005 19.620 2163.295 19.665 ;
        RECT 2208.990 19.620 2209.310 19.680 ;
        RECT 2163.005 19.480 2209.310 19.620 ;
        RECT 2163.005 19.435 2163.295 19.480 ;
        RECT 2208.990 19.420 2209.310 19.480 ;
        RECT 2042.010 18.800 2055.580 18.940 ;
        RECT 2042.010 18.740 2042.330 18.800 ;
        RECT 2114.245 15.880 2114.535 15.925 ;
        RECT 2163.005 15.880 2163.295 15.925 ;
        RECT 2114.245 15.740 2163.295 15.880 ;
        RECT 2114.245 15.695 2114.535 15.740 ;
        RECT 2163.005 15.695 2163.295 15.740 ;
      LAYER via ;
        RECT 2036.980 210.840 2037.240 211.100 ;
        RECT 2042.040 210.840 2042.300 211.100 ;
        RECT 2042.040 18.740 2042.300 19.000 ;
        RECT 2209.020 19.420 2209.280 19.680 ;
      LAYER met2 ;
        RECT 2037.020 220.000 2037.300 224.000 ;
        RECT 2037.040 211.130 2037.180 220.000 ;
        RECT 2036.980 210.810 2037.240 211.130 ;
        RECT 2042.040 210.810 2042.300 211.130 ;
        RECT 2042.100 19.030 2042.240 210.810 ;
        RECT 2209.020 19.390 2209.280 19.710 ;
        RECT 2042.040 18.710 2042.300 19.030 ;
        RECT 2209.080 2.400 2209.220 19.390 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2051.210 207.300 2051.530 207.360 ;
        RECT 2055.810 207.300 2056.130 207.360 ;
        RECT 2051.210 207.160 2056.130 207.300 ;
        RECT 2051.210 207.100 2051.530 207.160 ;
        RECT 2055.810 207.100 2056.130 207.160 ;
        RECT 2055.810 19.280 2056.130 19.340 ;
        RECT 2226.930 19.280 2227.250 19.340 ;
        RECT 2055.810 19.140 2227.250 19.280 ;
        RECT 2055.810 19.080 2056.130 19.140 ;
        RECT 2226.930 19.080 2227.250 19.140 ;
      LAYER via ;
        RECT 2051.240 207.100 2051.500 207.360 ;
        RECT 2055.840 207.100 2056.100 207.360 ;
        RECT 2055.840 19.080 2056.100 19.340 ;
        RECT 2226.960 19.080 2227.220 19.340 ;
      LAYER met2 ;
        RECT 2051.280 220.000 2051.560 224.000 ;
        RECT 2051.300 207.390 2051.440 220.000 ;
        RECT 2051.240 207.070 2051.500 207.390 ;
        RECT 2055.840 207.070 2056.100 207.390 ;
        RECT 2055.900 19.370 2056.040 207.070 ;
        RECT 2055.840 19.050 2056.100 19.370 ;
        RECT 2226.960 19.050 2227.220 19.370 ;
        RECT 2227.020 2.400 2227.160 19.050 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 786.210 209.340 786.530 209.400 ;
        RECT 861.190 209.340 861.510 209.400 ;
        RECT 786.210 209.200 861.510 209.340 ;
        RECT 786.210 209.140 786.530 209.200 ;
        RECT 861.190 209.140 861.510 209.200 ;
        RECT 781.610 17.580 781.930 17.640 ;
        RECT 786.210 17.580 786.530 17.640 ;
        RECT 781.610 17.440 786.530 17.580 ;
        RECT 781.610 17.380 781.930 17.440 ;
        RECT 786.210 17.380 786.530 17.440 ;
      LAYER via ;
        RECT 786.240 209.140 786.500 209.400 ;
        RECT 861.220 209.140 861.480 209.400 ;
        RECT 781.640 17.380 781.900 17.640 ;
        RECT 786.240 17.380 786.500 17.640 ;
      LAYER met2 ;
        RECT 861.260 220.000 861.540 224.000 ;
        RECT 861.280 209.430 861.420 220.000 ;
        RECT 786.240 209.110 786.500 209.430 ;
        RECT 861.220 209.110 861.480 209.430 ;
        RECT 786.300 17.670 786.440 209.110 ;
        RECT 781.640 17.350 781.900 17.670 ;
        RECT 786.240 17.350 786.500 17.670 ;
        RECT 781.700 2.400 781.840 17.350 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2069.610 18.600 2069.930 18.660 ;
        RECT 2244.870 18.600 2245.190 18.660 ;
        RECT 2069.610 18.460 2245.190 18.600 ;
        RECT 2069.610 18.400 2069.930 18.460 ;
        RECT 2244.870 18.400 2245.190 18.460 ;
      LAYER via ;
        RECT 2069.640 18.400 2069.900 18.660 ;
        RECT 2244.900 18.400 2245.160 18.660 ;
      LAYER met2 ;
        RECT 2066.000 220.730 2066.280 224.000 ;
        RECT 2066.000 220.590 2069.840 220.730 ;
        RECT 2066.000 220.000 2066.280 220.590 ;
        RECT 2069.700 18.690 2069.840 220.590 ;
        RECT 2069.640 18.370 2069.900 18.690 ;
        RECT 2244.900 18.370 2245.160 18.690 ;
        RECT 2244.960 2.400 2245.100 18.370 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2114.765 18.785 2114.935 19.635 ;
        RECT 2158.465 18.785 2158.635 19.635 ;
        RECT 2187.445 18.785 2187.615 20.995 ;
        RECT 2227.465 19.125 2227.635 20.995 ;
      LAYER mcon ;
        RECT 2187.445 20.825 2187.615 20.995 ;
        RECT 2114.765 19.465 2114.935 19.635 ;
        RECT 2158.465 19.465 2158.635 19.635 ;
        RECT 2227.465 20.825 2227.635 20.995 ;
      LAYER met1 ;
        RECT 2187.385 20.980 2187.675 21.025 ;
        RECT 2227.405 20.980 2227.695 21.025 ;
        RECT 2187.385 20.840 2227.695 20.980 ;
        RECT 2187.385 20.795 2187.675 20.840 ;
        RECT 2227.405 20.795 2227.695 20.840 ;
        RECT 2114.705 19.620 2114.995 19.665 ;
        RECT 2158.405 19.620 2158.695 19.665 ;
        RECT 2114.705 19.480 2158.695 19.620 ;
        RECT 2114.705 19.435 2114.995 19.480 ;
        RECT 2158.405 19.435 2158.695 19.480 ;
        RECT 2227.405 19.280 2227.695 19.325 ;
        RECT 2262.350 19.280 2262.670 19.340 ;
        RECT 2227.405 19.140 2262.670 19.280 ;
        RECT 2227.405 19.095 2227.695 19.140 ;
        RECT 2262.350 19.080 2262.670 19.140 ;
        RECT 2083.410 18.940 2083.730 19.000 ;
        RECT 2114.705 18.940 2114.995 18.985 ;
        RECT 2083.410 18.800 2114.995 18.940 ;
        RECT 2083.410 18.740 2083.730 18.800 ;
        RECT 2114.705 18.755 2114.995 18.800 ;
        RECT 2158.405 18.940 2158.695 18.985 ;
        RECT 2187.385 18.940 2187.675 18.985 ;
        RECT 2158.405 18.800 2187.675 18.940 ;
        RECT 2158.405 18.755 2158.695 18.800 ;
        RECT 2187.385 18.755 2187.675 18.800 ;
      LAYER via ;
        RECT 2262.380 19.080 2262.640 19.340 ;
        RECT 2083.440 18.740 2083.700 19.000 ;
      LAYER met2 ;
        RECT 2080.720 220.730 2081.000 224.000 ;
        RECT 2080.720 220.590 2083.640 220.730 ;
        RECT 2080.720 220.000 2081.000 220.590 ;
        RECT 2083.500 19.030 2083.640 220.590 ;
        RECT 2262.380 19.050 2262.640 19.370 ;
        RECT 2083.440 18.710 2083.700 19.030 ;
        RECT 2262.440 2.400 2262.580 19.050 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2097.210 17.920 2097.530 17.980 ;
        RECT 2280.290 17.920 2280.610 17.980 ;
        RECT 2097.210 17.780 2280.610 17.920 ;
        RECT 2097.210 17.720 2097.530 17.780 ;
        RECT 2280.290 17.720 2280.610 17.780 ;
      LAYER via ;
        RECT 2097.240 17.720 2097.500 17.980 ;
        RECT 2280.320 17.720 2280.580 17.980 ;
      LAYER met2 ;
        RECT 2095.440 220.730 2095.720 224.000 ;
        RECT 2095.440 220.590 2097.440 220.730 ;
        RECT 2095.440 220.000 2095.720 220.590 ;
        RECT 2097.300 18.010 2097.440 220.590 ;
        RECT 2097.240 17.690 2097.500 18.010 ;
        RECT 2280.320 17.690 2280.580 18.010 ;
        RECT 2280.380 2.400 2280.520 17.690 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2259.665 17.085 2259.835 18.275 ;
      LAYER mcon ;
        RECT 2259.665 18.105 2259.835 18.275 ;
      LAYER met1 ;
        RECT 2259.605 18.260 2259.895 18.305 ;
        RECT 2297.770 18.260 2298.090 18.320 ;
        RECT 2259.605 18.120 2298.090 18.260 ;
        RECT 2259.605 18.075 2259.895 18.120 ;
        RECT 2297.770 18.060 2298.090 18.120 ;
        RECT 2111.010 17.240 2111.330 17.300 ;
        RECT 2259.605 17.240 2259.895 17.285 ;
        RECT 2111.010 17.100 2259.895 17.240 ;
        RECT 2111.010 17.040 2111.330 17.100 ;
        RECT 2259.605 17.055 2259.895 17.100 ;
      LAYER via ;
        RECT 2297.800 18.060 2298.060 18.320 ;
        RECT 2111.040 17.040 2111.300 17.300 ;
      LAYER met2 ;
        RECT 2110.160 220.730 2110.440 224.000 ;
        RECT 2110.160 220.590 2111.240 220.730 ;
        RECT 2110.160 220.000 2110.440 220.590 ;
        RECT 2111.100 17.330 2111.240 220.590 ;
        RECT 2297.800 18.030 2298.060 18.350 ;
        RECT 2111.040 17.010 2111.300 17.330 ;
        RECT 2297.860 16.730 2298.000 18.030 ;
        RECT 2297.860 16.590 2298.460 16.730 ;
        RECT 2298.320 2.400 2298.460 16.590 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2124.810 17.580 2125.130 17.640 ;
        RECT 2124.810 17.440 2309.500 17.580 ;
        RECT 2124.810 17.380 2125.130 17.440 ;
        RECT 2309.360 17.240 2309.500 17.440 ;
        RECT 2316.170 17.240 2316.490 17.300 ;
        RECT 2309.360 17.100 2316.490 17.240 ;
        RECT 2316.170 17.040 2316.490 17.100 ;
      LAYER via ;
        RECT 2124.840 17.380 2125.100 17.640 ;
        RECT 2316.200 17.040 2316.460 17.300 ;
      LAYER met2 ;
        RECT 2124.880 220.000 2125.160 224.000 ;
        RECT 2124.900 17.670 2125.040 220.000 ;
        RECT 2124.840 17.350 2125.100 17.670 ;
        RECT 2316.200 17.010 2316.460 17.330 ;
        RECT 2316.260 2.400 2316.400 17.010 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2162.145 16.405 2162.315 19.975 ;
        RECT 2174.105 15.385 2174.275 16.575 ;
      LAYER mcon ;
        RECT 2162.145 19.805 2162.315 19.975 ;
        RECT 2174.105 16.405 2174.275 16.575 ;
      LAYER met1 ;
        RECT 2139.530 207.300 2139.850 207.360 ;
        RECT 2145.510 207.300 2145.830 207.360 ;
        RECT 2139.530 207.160 2145.830 207.300 ;
        RECT 2139.530 207.100 2139.850 207.160 ;
        RECT 2145.510 207.100 2145.830 207.160 ;
        RECT 2145.510 19.960 2145.830 20.020 ;
        RECT 2162.085 19.960 2162.375 20.005 ;
        RECT 2145.510 19.820 2162.375 19.960 ;
        RECT 2145.510 19.760 2145.830 19.820 ;
        RECT 2162.085 19.775 2162.375 19.820 ;
        RECT 2162.085 16.560 2162.375 16.605 ;
        RECT 2174.045 16.560 2174.335 16.605 ;
        RECT 2162.085 16.420 2174.335 16.560 ;
        RECT 2162.085 16.375 2162.375 16.420 ;
        RECT 2174.045 16.375 2174.335 16.420 ;
        RECT 2174.045 15.540 2174.335 15.585 ;
        RECT 2334.110 15.540 2334.430 15.600 ;
        RECT 2174.045 15.400 2334.430 15.540 ;
        RECT 2174.045 15.355 2174.335 15.400 ;
        RECT 2334.110 15.340 2334.430 15.400 ;
      LAYER via ;
        RECT 2139.560 207.100 2139.820 207.360 ;
        RECT 2145.540 207.100 2145.800 207.360 ;
        RECT 2145.540 19.760 2145.800 20.020 ;
        RECT 2334.140 15.340 2334.400 15.600 ;
      LAYER met2 ;
        RECT 2139.600 220.000 2139.880 224.000 ;
        RECT 2139.620 207.390 2139.760 220.000 ;
        RECT 2139.560 207.070 2139.820 207.390 ;
        RECT 2145.540 207.070 2145.800 207.390 ;
        RECT 2145.600 20.050 2145.740 207.070 ;
        RECT 2145.540 19.730 2145.800 20.050 ;
        RECT 2334.140 15.310 2334.400 15.630 ;
        RECT 2334.200 2.400 2334.340 15.310 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2172.265 13.685 2172.435 14.875 ;
        RECT 2207.685 13.685 2207.855 15.215 ;
      LAYER mcon ;
        RECT 2207.685 15.045 2207.855 15.215 ;
        RECT 2172.265 14.705 2172.435 14.875 ;
      LAYER met1 ;
        RECT 2154.250 207.300 2154.570 207.360 ;
        RECT 2159.310 207.300 2159.630 207.360 ;
        RECT 2154.250 207.160 2159.630 207.300 ;
        RECT 2154.250 207.100 2154.570 207.160 ;
        RECT 2159.310 207.100 2159.630 207.160 ;
        RECT 2207.625 15.200 2207.915 15.245 ;
        RECT 2351.590 15.200 2351.910 15.260 ;
        RECT 2207.625 15.060 2351.910 15.200 ;
        RECT 2207.625 15.015 2207.915 15.060 ;
        RECT 2351.590 15.000 2351.910 15.060 ;
        RECT 2159.310 14.860 2159.630 14.920 ;
        RECT 2172.205 14.860 2172.495 14.905 ;
        RECT 2159.310 14.720 2172.495 14.860 ;
        RECT 2159.310 14.660 2159.630 14.720 ;
        RECT 2172.205 14.675 2172.495 14.720 ;
        RECT 2172.205 13.840 2172.495 13.885 ;
        RECT 2207.625 13.840 2207.915 13.885 ;
        RECT 2172.205 13.700 2207.915 13.840 ;
        RECT 2172.205 13.655 2172.495 13.700 ;
        RECT 2207.625 13.655 2207.915 13.700 ;
      LAYER via ;
        RECT 2154.280 207.100 2154.540 207.360 ;
        RECT 2159.340 207.100 2159.600 207.360 ;
        RECT 2351.620 15.000 2351.880 15.260 ;
        RECT 2159.340 14.660 2159.600 14.920 ;
      LAYER met2 ;
        RECT 2154.320 220.000 2154.600 224.000 ;
        RECT 2154.340 207.390 2154.480 220.000 ;
        RECT 2154.280 207.070 2154.540 207.390 ;
        RECT 2159.340 207.070 2159.600 207.390 ;
        RECT 2159.400 14.950 2159.540 207.070 ;
        RECT 2351.620 14.970 2351.880 15.290 ;
        RECT 2159.340 14.630 2159.600 14.950 ;
        RECT 2351.680 2.400 2351.820 14.970 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2168.970 207.300 2169.290 207.360 ;
        RECT 2173.110 207.300 2173.430 207.360 ;
        RECT 2168.970 207.160 2173.430 207.300 ;
        RECT 2168.970 207.100 2169.290 207.160 ;
        RECT 2173.110 207.100 2173.430 207.160 ;
        RECT 2211.290 16.560 2211.610 16.620 ;
        RECT 2369.530 16.560 2369.850 16.620 ;
        RECT 2211.290 16.420 2369.850 16.560 ;
        RECT 2211.290 16.360 2211.610 16.420 ;
        RECT 2369.530 16.360 2369.850 16.420 ;
        RECT 2172.650 15.880 2172.970 15.940 ;
        RECT 2211.290 15.880 2211.610 15.940 ;
        RECT 2172.650 15.740 2211.610 15.880 ;
        RECT 2172.650 15.680 2172.970 15.740 ;
        RECT 2211.290 15.680 2211.610 15.740 ;
      LAYER via ;
        RECT 2169.000 207.100 2169.260 207.360 ;
        RECT 2173.140 207.100 2173.400 207.360 ;
        RECT 2211.320 16.360 2211.580 16.620 ;
        RECT 2369.560 16.360 2369.820 16.620 ;
        RECT 2172.680 15.680 2172.940 15.940 ;
        RECT 2211.320 15.680 2211.580 15.940 ;
      LAYER met2 ;
        RECT 2169.040 220.000 2169.320 224.000 ;
        RECT 2169.060 207.390 2169.200 220.000 ;
        RECT 2169.000 207.070 2169.260 207.390 ;
        RECT 2173.140 207.070 2173.400 207.390 ;
        RECT 2173.200 39.170 2173.340 207.070 ;
        RECT 2172.740 39.030 2173.340 39.170 ;
        RECT 2172.740 15.970 2172.880 39.030 ;
        RECT 2211.320 16.330 2211.580 16.650 ;
        RECT 2369.560 16.330 2369.820 16.650 ;
        RECT 2211.380 15.970 2211.520 16.330 ;
        RECT 2172.680 15.650 2172.940 15.970 ;
        RECT 2211.320 15.650 2211.580 15.970 ;
        RECT 2369.620 2.400 2369.760 16.330 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2248.165 18.445 2248.335 19.635 ;
        RECT 2258.745 14.025 2258.915 18.615 ;
      LAYER mcon ;
        RECT 2248.165 19.465 2248.335 19.635 ;
        RECT 2258.745 18.445 2258.915 18.615 ;
      LAYER met1 ;
        RECT 2183.690 207.640 2184.010 207.700 ;
        RECT 2218.190 207.640 2218.510 207.700 ;
        RECT 2183.690 207.500 2218.510 207.640 ;
        RECT 2183.690 207.440 2184.010 207.500 ;
        RECT 2218.190 207.440 2218.510 207.500 ;
        RECT 2218.190 19.620 2218.510 19.680 ;
        RECT 2248.105 19.620 2248.395 19.665 ;
        RECT 2218.190 19.480 2248.395 19.620 ;
        RECT 2218.190 19.420 2218.510 19.480 ;
        RECT 2248.105 19.435 2248.395 19.480 ;
        RECT 2248.105 18.600 2248.395 18.645 ;
        RECT 2258.685 18.600 2258.975 18.645 ;
        RECT 2248.105 18.460 2258.975 18.600 ;
        RECT 2248.105 18.415 2248.395 18.460 ;
        RECT 2258.685 18.415 2258.975 18.460 ;
        RECT 2258.685 14.180 2258.975 14.225 ;
        RECT 2387.470 14.180 2387.790 14.240 ;
        RECT 2258.685 14.040 2387.790 14.180 ;
        RECT 2258.685 13.995 2258.975 14.040 ;
        RECT 2387.470 13.980 2387.790 14.040 ;
      LAYER via ;
        RECT 2183.720 207.440 2183.980 207.700 ;
        RECT 2218.220 207.440 2218.480 207.700 ;
        RECT 2218.220 19.420 2218.480 19.680 ;
        RECT 2387.500 13.980 2387.760 14.240 ;
      LAYER met2 ;
        RECT 2183.760 220.000 2184.040 224.000 ;
        RECT 2183.780 207.730 2183.920 220.000 ;
        RECT 2183.720 207.410 2183.980 207.730 ;
        RECT 2218.220 207.410 2218.480 207.730 ;
        RECT 2218.280 19.710 2218.420 207.410 ;
        RECT 2218.220 19.390 2218.480 19.710 ;
        RECT 2387.500 13.950 2387.760 14.270 ;
        RECT 2387.560 2.400 2387.700 13.950 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2200.710 20.300 2201.030 20.360 ;
        RECT 2405.410 20.300 2405.730 20.360 ;
        RECT 2200.710 20.160 2405.730 20.300 ;
        RECT 2200.710 20.100 2201.030 20.160 ;
        RECT 2405.410 20.100 2405.730 20.160 ;
      LAYER via ;
        RECT 2200.740 20.100 2201.000 20.360 ;
        RECT 2405.440 20.100 2405.700 20.360 ;
      LAYER met2 ;
        RECT 2198.480 220.730 2198.760 224.000 ;
        RECT 2198.480 220.590 2200.940 220.730 ;
        RECT 2198.480 220.000 2198.760 220.590 ;
        RECT 2200.800 20.390 2200.940 220.590 ;
        RECT 2200.740 20.070 2201.000 20.390 ;
        RECT 2405.440 20.070 2405.700 20.390 ;
        RECT 2405.500 2.400 2405.640 20.070 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 800.010 209.680 800.330 209.740 ;
        RECT 874.070 209.680 874.390 209.740 ;
        RECT 800.010 209.540 874.390 209.680 ;
        RECT 800.010 209.480 800.330 209.540 ;
        RECT 874.070 209.480 874.390 209.540 ;
      LAYER via ;
        RECT 800.040 209.480 800.300 209.740 ;
        RECT 874.100 209.480 874.360 209.740 ;
      LAYER met2 ;
        RECT 875.980 220.730 876.260 224.000 ;
        RECT 874.160 220.590 876.260 220.730 ;
        RECT 874.160 209.770 874.300 220.590 ;
        RECT 875.980 220.000 876.260 220.590 ;
        RECT 800.040 209.450 800.300 209.770 ;
        RECT 874.100 209.450 874.360 209.770 ;
        RECT 800.100 17.410 800.240 209.450 ;
        RECT 799.640 17.270 800.240 17.410 ;
        RECT 799.640 2.400 799.780 17.270 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.210 213.420 648.530 213.480 ;
        RECT 748.490 213.420 748.810 213.480 ;
        RECT 648.210 213.280 656.260 213.420 ;
        RECT 648.210 213.220 648.530 213.280 ;
        RECT 656.120 213.080 656.260 213.280 ;
        RECT 679.580 213.280 748.810 213.420 ;
        RECT 679.580 213.080 679.720 213.280 ;
        RECT 748.490 213.220 748.810 213.280 ;
        RECT 656.120 212.940 679.720 213.080 ;
        RECT 644.990 15.200 645.310 15.260 ;
        RECT 648.210 15.200 648.530 15.260 ;
        RECT 644.990 15.060 648.530 15.200 ;
        RECT 644.990 15.000 645.310 15.060 ;
        RECT 648.210 15.000 648.530 15.060 ;
      LAYER via ;
        RECT 648.240 213.220 648.500 213.480 ;
        RECT 748.520 213.220 748.780 213.480 ;
        RECT 645.020 15.000 645.280 15.260 ;
        RECT 648.240 15.000 648.500 15.260 ;
      LAYER met2 ;
        RECT 748.560 220.000 748.840 224.000 ;
        RECT 748.580 213.510 748.720 220.000 ;
        RECT 648.240 213.190 648.500 213.510 ;
        RECT 748.520 213.190 748.780 213.510 ;
        RECT 648.300 15.290 648.440 213.190 ;
        RECT 645.020 14.970 645.280 15.290 ;
        RECT 648.240 14.970 648.500 15.290 ;
        RECT 645.080 2.400 645.220 14.970 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2217.730 210.700 2218.050 210.760 ;
        RECT 2428.870 210.700 2429.190 210.760 ;
        RECT 2217.730 210.560 2429.190 210.700 ;
        RECT 2217.730 210.500 2218.050 210.560 ;
        RECT 2428.870 210.500 2429.190 210.560 ;
      LAYER via ;
        RECT 2217.760 210.500 2218.020 210.760 ;
        RECT 2428.900 210.500 2429.160 210.760 ;
      LAYER met2 ;
        RECT 2217.800 220.000 2218.080 224.000 ;
        RECT 2217.820 210.790 2217.960 220.000 ;
        RECT 2217.760 210.470 2218.020 210.790 ;
        RECT 2428.900 210.470 2429.160 210.790 ;
        RECT 2428.960 2.400 2429.100 210.470 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2232.450 209.340 2232.770 209.400 ;
        RECT 2432.090 209.340 2432.410 209.400 ;
        RECT 2232.450 209.200 2432.410 209.340 ;
        RECT 2232.450 209.140 2232.770 209.200 ;
        RECT 2432.090 209.140 2432.410 209.200 ;
        RECT 2432.090 16.900 2432.410 16.960 ;
        RECT 2446.810 16.900 2447.130 16.960 ;
        RECT 2432.090 16.760 2447.130 16.900 ;
        RECT 2432.090 16.700 2432.410 16.760 ;
        RECT 2446.810 16.700 2447.130 16.760 ;
      LAYER via ;
        RECT 2232.480 209.140 2232.740 209.400 ;
        RECT 2432.120 209.140 2432.380 209.400 ;
        RECT 2432.120 16.700 2432.380 16.960 ;
        RECT 2446.840 16.700 2447.100 16.960 ;
      LAYER met2 ;
        RECT 2232.520 220.000 2232.800 224.000 ;
        RECT 2232.540 209.430 2232.680 220.000 ;
        RECT 2232.480 209.110 2232.740 209.430 ;
        RECT 2432.120 209.110 2432.380 209.430 ;
        RECT 2432.180 16.990 2432.320 209.110 ;
        RECT 2432.120 16.670 2432.380 16.990 ;
        RECT 2446.840 16.670 2447.100 16.990 ;
        RECT 2446.900 2.400 2447.040 16.670 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2259.205 18.955 2259.375 19.635 ;
        RECT 2259.205 18.785 2263.515 18.955 ;
      LAYER mcon ;
        RECT 2259.205 19.465 2259.375 19.635 ;
        RECT 2263.345 18.785 2263.515 18.955 ;
      LAYER met1 ;
        RECT 2249.010 19.620 2249.330 19.680 ;
        RECT 2259.145 19.620 2259.435 19.665 ;
        RECT 2249.010 19.480 2259.435 19.620 ;
        RECT 2249.010 19.420 2249.330 19.480 ;
        RECT 2259.145 19.435 2259.435 19.480 ;
        RECT 2263.285 18.940 2263.575 18.985 ;
        RECT 2263.285 18.800 2269.940 18.940 ;
        RECT 2263.285 18.755 2263.575 18.800 ;
        RECT 2269.800 18.600 2269.940 18.800 ;
        RECT 2464.750 18.600 2465.070 18.660 ;
        RECT 2269.800 18.460 2465.070 18.600 ;
        RECT 2464.750 18.400 2465.070 18.460 ;
      LAYER via ;
        RECT 2249.040 19.420 2249.300 19.680 ;
        RECT 2464.780 18.400 2465.040 18.660 ;
      LAYER met2 ;
        RECT 2247.240 220.730 2247.520 224.000 ;
        RECT 2247.240 220.590 2249.240 220.730 ;
        RECT 2247.240 220.000 2247.520 220.590 ;
        RECT 2249.100 19.710 2249.240 220.590 ;
        RECT 2249.040 19.390 2249.300 19.710 ;
        RECT 2464.780 18.370 2465.040 18.690 ;
        RECT 2464.840 2.400 2464.980 18.370 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2261.890 213.080 2262.210 213.140 ;
        RECT 2473.490 213.080 2473.810 213.140 ;
        RECT 2261.890 212.940 2473.810 213.080 ;
        RECT 2261.890 212.880 2262.210 212.940 ;
        RECT 2473.490 212.880 2473.810 212.940 ;
        RECT 2473.490 18.600 2473.810 18.660 ;
        RECT 2482.690 18.600 2483.010 18.660 ;
        RECT 2473.490 18.460 2483.010 18.600 ;
        RECT 2473.490 18.400 2473.810 18.460 ;
        RECT 2482.690 18.400 2483.010 18.460 ;
      LAYER via ;
        RECT 2261.920 212.880 2262.180 213.140 ;
        RECT 2473.520 212.880 2473.780 213.140 ;
        RECT 2473.520 18.400 2473.780 18.660 ;
        RECT 2482.720 18.400 2482.980 18.660 ;
      LAYER met2 ;
        RECT 2261.960 220.000 2262.240 224.000 ;
        RECT 2261.980 213.170 2262.120 220.000 ;
        RECT 2261.920 212.850 2262.180 213.170 ;
        RECT 2473.520 212.850 2473.780 213.170 ;
        RECT 2473.580 18.690 2473.720 212.850 ;
        RECT 2473.520 18.370 2473.780 18.690 ;
        RECT 2482.720 18.370 2482.980 18.690 ;
        RECT 2482.780 2.400 2482.920 18.370 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2276.610 213.760 2276.930 213.820 ;
        RECT 2498.330 213.760 2498.650 213.820 ;
        RECT 2276.610 213.620 2498.650 213.760 ;
        RECT 2276.610 213.560 2276.930 213.620 ;
        RECT 2498.330 213.560 2498.650 213.620 ;
        RECT 2498.330 2.960 2498.650 3.020 ;
        RECT 2500.630 2.960 2500.950 3.020 ;
        RECT 2498.330 2.820 2500.950 2.960 ;
        RECT 2498.330 2.760 2498.650 2.820 ;
        RECT 2500.630 2.760 2500.950 2.820 ;
      LAYER via ;
        RECT 2276.640 213.560 2276.900 213.820 ;
        RECT 2498.360 213.560 2498.620 213.820 ;
        RECT 2498.360 2.760 2498.620 3.020 ;
        RECT 2500.660 2.760 2500.920 3.020 ;
      LAYER met2 ;
        RECT 2276.680 220.000 2276.960 224.000 ;
        RECT 2276.700 213.850 2276.840 220.000 ;
        RECT 2276.640 213.530 2276.900 213.850 ;
        RECT 2498.360 213.530 2498.620 213.850 ;
        RECT 2498.420 3.050 2498.560 213.530 ;
        RECT 2498.360 2.730 2498.620 3.050 ;
        RECT 2500.660 2.730 2500.920 3.050 ;
        RECT 2500.720 2.400 2500.860 2.730 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2291.330 209.680 2291.650 209.740 ;
        RECT 2512.130 209.680 2512.450 209.740 ;
        RECT 2291.330 209.540 2512.450 209.680 ;
        RECT 2291.330 209.480 2291.650 209.540 ;
        RECT 2512.130 209.480 2512.450 209.540 ;
        RECT 2512.130 18.600 2512.450 18.660 ;
        RECT 2518.110 18.600 2518.430 18.660 ;
        RECT 2512.130 18.460 2518.430 18.600 ;
        RECT 2512.130 18.400 2512.450 18.460 ;
        RECT 2518.110 18.400 2518.430 18.460 ;
      LAYER via ;
        RECT 2291.360 209.480 2291.620 209.740 ;
        RECT 2512.160 209.480 2512.420 209.740 ;
        RECT 2512.160 18.400 2512.420 18.660 ;
        RECT 2518.140 18.400 2518.400 18.660 ;
      LAYER met2 ;
        RECT 2291.400 220.000 2291.680 224.000 ;
        RECT 2291.420 209.770 2291.560 220.000 ;
        RECT 2291.360 209.450 2291.620 209.770 ;
        RECT 2512.160 209.450 2512.420 209.770 ;
        RECT 2512.220 18.690 2512.360 209.450 ;
        RECT 2512.160 18.370 2512.420 18.690 ;
        RECT 2518.140 18.370 2518.400 18.690 ;
        RECT 2518.200 2.400 2518.340 18.370 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2306.050 213.420 2306.370 213.480 ;
        RECT 2532.370 213.420 2532.690 213.480 ;
        RECT 2306.050 213.280 2532.690 213.420 ;
        RECT 2306.050 213.220 2306.370 213.280 ;
        RECT 2532.370 213.220 2532.690 213.280 ;
        RECT 2532.370 2.960 2532.690 3.020 ;
        RECT 2536.050 2.960 2536.370 3.020 ;
        RECT 2532.370 2.820 2536.370 2.960 ;
        RECT 2532.370 2.760 2532.690 2.820 ;
        RECT 2536.050 2.760 2536.370 2.820 ;
      LAYER via ;
        RECT 2306.080 213.220 2306.340 213.480 ;
        RECT 2532.400 213.220 2532.660 213.480 ;
        RECT 2532.400 2.760 2532.660 3.020 ;
        RECT 2536.080 2.760 2536.340 3.020 ;
      LAYER met2 ;
        RECT 2306.120 220.000 2306.400 224.000 ;
        RECT 2306.140 213.510 2306.280 220.000 ;
        RECT 2306.080 213.190 2306.340 213.510 ;
        RECT 2532.400 213.190 2532.660 213.510 ;
        RECT 2532.460 3.050 2532.600 213.190 ;
        RECT 2532.400 2.730 2532.660 3.050 ;
        RECT 2536.080 2.730 2536.340 3.050 ;
        RECT 2536.140 2.400 2536.280 2.730 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2320.770 210.020 2321.090 210.080 ;
        RECT 2542.490 210.020 2542.810 210.080 ;
        RECT 2320.770 209.880 2542.810 210.020 ;
        RECT 2320.770 209.820 2321.090 209.880 ;
        RECT 2542.490 209.820 2542.810 209.880 ;
        RECT 2542.490 19.620 2542.810 19.680 ;
        RECT 2553.990 19.620 2554.310 19.680 ;
        RECT 2542.490 19.480 2554.310 19.620 ;
        RECT 2542.490 19.420 2542.810 19.480 ;
        RECT 2553.990 19.420 2554.310 19.480 ;
      LAYER via ;
        RECT 2320.800 209.820 2321.060 210.080 ;
        RECT 2542.520 209.820 2542.780 210.080 ;
        RECT 2542.520 19.420 2542.780 19.680 ;
        RECT 2554.020 19.420 2554.280 19.680 ;
      LAYER met2 ;
        RECT 2320.840 220.000 2321.120 224.000 ;
        RECT 2320.860 210.110 2321.000 220.000 ;
        RECT 2320.800 209.790 2321.060 210.110 ;
        RECT 2542.520 209.790 2542.780 210.110 ;
        RECT 2542.580 19.710 2542.720 209.790 ;
        RECT 2542.520 19.390 2542.780 19.710 ;
        RECT 2554.020 19.390 2554.280 19.710 ;
        RECT 2554.080 2.400 2554.220 19.390 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2335.490 212.400 2335.810 212.460 ;
        RECT 2563.190 212.400 2563.510 212.460 ;
        RECT 2335.490 212.260 2563.510 212.400 ;
        RECT 2335.490 212.200 2335.810 212.260 ;
        RECT 2563.190 212.200 2563.510 212.260 ;
        RECT 2563.190 17.580 2563.510 17.640 ;
        RECT 2571.930 17.580 2572.250 17.640 ;
        RECT 2563.190 17.440 2572.250 17.580 ;
        RECT 2563.190 17.380 2563.510 17.440 ;
        RECT 2571.930 17.380 2572.250 17.440 ;
      LAYER via ;
        RECT 2335.520 212.200 2335.780 212.460 ;
        RECT 2563.220 212.200 2563.480 212.460 ;
        RECT 2563.220 17.380 2563.480 17.640 ;
        RECT 2571.960 17.380 2572.220 17.640 ;
      LAYER met2 ;
        RECT 2335.560 220.000 2335.840 224.000 ;
        RECT 2335.580 212.490 2335.720 220.000 ;
        RECT 2335.520 212.170 2335.780 212.490 ;
        RECT 2563.220 212.170 2563.480 212.490 ;
        RECT 2563.280 17.670 2563.420 212.170 ;
        RECT 2563.220 17.350 2563.480 17.670 ;
        RECT 2571.960 17.350 2572.220 17.670 ;
        RECT 2572.020 2.400 2572.160 17.350 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2555.445 17.085 2555.615 17.935 ;
      LAYER mcon ;
        RECT 2555.445 17.765 2555.615 17.935 ;
      LAYER met1 ;
        RECT 2555.385 17.920 2555.675 17.965 ;
        RECT 2589.410 17.920 2589.730 17.980 ;
        RECT 2555.385 17.780 2589.730 17.920 ;
        RECT 2555.385 17.735 2555.675 17.780 ;
        RECT 2589.410 17.720 2589.730 17.780 ;
        RECT 2352.510 17.240 2352.830 17.300 ;
        RECT 2555.385 17.240 2555.675 17.285 ;
        RECT 2352.510 17.100 2555.675 17.240 ;
        RECT 2352.510 17.040 2352.830 17.100 ;
        RECT 2555.385 17.055 2555.675 17.100 ;
      LAYER via ;
        RECT 2589.440 17.720 2589.700 17.980 ;
        RECT 2352.540 17.040 2352.800 17.300 ;
      LAYER met2 ;
        RECT 2350.280 220.730 2350.560 224.000 ;
        RECT 2350.280 220.590 2352.740 220.730 ;
        RECT 2350.280 220.000 2350.560 220.590 ;
        RECT 2352.600 17.330 2352.740 220.590 ;
        RECT 2589.440 17.690 2589.700 18.010 ;
        RECT 2352.540 17.010 2352.800 17.330 ;
        RECT 2589.500 2.400 2589.640 17.690 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 827.610 211.380 827.930 211.440 ;
        RECT 895.690 211.380 896.010 211.440 ;
        RECT 827.610 211.240 896.010 211.380 ;
        RECT 827.610 211.180 827.930 211.240 ;
        RECT 895.690 211.180 896.010 211.240 ;
        RECT 823.470 17.240 823.790 17.300 ;
        RECT 827.610 17.240 827.930 17.300 ;
        RECT 823.470 17.100 827.930 17.240 ;
        RECT 823.470 17.040 823.790 17.100 ;
        RECT 827.610 17.040 827.930 17.100 ;
      LAYER via ;
        RECT 827.640 211.180 827.900 211.440 ;
        RECT 895.720 211.180 895.980 211.440 ;
        RECT 823.500 17.040 823.760 17.300 ;
        RECT 827.640 17.040 827.900 17.300 ;
      LAYER met2 ;
        RECT 895.760 220.000 896.040 224.000 ;
        RECT 895.780 211.470 895.920 220.000 ;
        RECT 827.640 211.150 827.900 211.470 ;
        RECT 895.720 211.150 895.980 211.470 ;
        RECT 827.700 17.330 827.840 211.150 ;
        RECT 823.500 17.010 823.760 17.330 ;
        RECT 827.640 17.010 827.900 17.330 ;
        RECT 823.560 2.400 823.700 17.010 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2364.930 211.720 2365.250 211.780 ;
        RECT 2602.290 211.720 2602.610 211.780 ;
        RECT 2364.930 211.580 2602.610 211.720 ;
        RECT 2364.930 211.520 2365.250 211.580 ;
        RECT 2602.290 211.520 2602.610 211.580 ;
      LAYER via ;
        RECT 2364.960 211.520 2365.220 211.780 ;
        RECT 2602.320 211.520 2602.580 211.780 ;
      LAYER met2 ;
        RECT 2365.000 220.000 2365.280 224.000 ;
        RECT 2365.020 211.810 2365.160 220.000 ;
        RECT 2364.960 211.490 2365.220 211.810 ;
        RECT 2602.320 211.490 2602.580 211.810 ;
        RECT 2602.380 17.410 2602.520 211.490 ;
        RECT 2602.380 17.270 2607.580 17.410 ;
        RECT 2607.440 2.400 2607.580 17.270 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2379.650 208.660 2379.970 208.720 ;
        RECT 2480.390 208.660 2480.710 208.720 ;
        RECT 2379.650 208.520 2480.710 208.660 ;
        RECT 2379.650 208.460 2379.970 208.520 ;
        RECT 2480.390 208.460 2480.710 208.520 ;
        RECT 2480.390 14.520 2480.710 14.580 ;
        RECT 2625.290 14.520 2625.610 14.580 ;
        RECT 2480.390 14.380 2625.610 14.520 ;
        RECT 2480.390 14.320 2480.710 14.380 ;
        RECT 2625.290 14.320 2625.610 14.380 ;
      LAYER via ;
        RECT 2379.680 208.460 2379.940 208.720 ;
        RECT 2480.420 208.460 2480.680 208.720 ;
        RECT 2480.420 14.320 2480.680 14.580 ;
        RECT 2625.320 14.320 2625.580 14.580 ;
      LAYER met2 ;
        RECT 2379.720 220.000 2380.000 224.000 ;
        RECT 2379.740 208.750 2379.880 220.000 ;
        RECT 2379.680 208.430 2379.940 208.750 ;
        RECT 2480.420 208.430 2480.680 208.750 ;
        RECT 2480.480 14.610 2480.620 208.430 ;
        RECT 2480.420 14.290 2480.680 14.610 ;
        RECT 2625.320 14.290 2625.580 14.610 ;
        RECT 2625.380 2.400 2625.520 14.290 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2394.370 211.380 2394.690 211.440 ;
        RECT 2642.770 211.380 2643.090 211.440 ;
        RECT 2394.370 211.240 2643.090 211.380 ;
        RECT 2394.370 211.180 2394.690 211.240 ;
        RECT 2642.770 211.180 2643.090 211.240 ;
      LAYER via ;
        RECT 2394.400 211.180 2394.660 211.440 ;
        RECT 2642.800 211.180 2643.060 211.440 ;
      LAYER met2 ;
        RECT 2394.440 220.000 2394.720 224.000 ;
        RECT 2394.460 211.470 2394.600 220.000 ;
        RECT 2394.400 211.150 2394.660 211.470 ;
        RECT 2642.800 211.150 2643.060 211.470 ;
        RECT 2642.860 17.410 2643.000 211.150 ;
        RECT 2642.860 17.270 2643.460 17.410 ;
        RECT 2643.320 2.400 2643.460 17.270 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2409.090 207.300 2409.410 207.360 ;
        RECT 2414.610 207.300 2414.930 207.360 ;
        RECT 2409.090 207.160 2414.930 207.300 ;
        RECT 2409.090 207.100 2409.410 207.160 ;
        RECT 2414.610 207.100 2414.930 207.160 ;
        RECT 2414.610 15.880 2414.930 15.940 ;
        RECT 2661.170 15.880 2661.490 15.940 ;
        RECT 2414.610 15.740 2661.490 15.880 ;
        RECT 2414.610 15.680 2414.930 15.740 ;
        RECT 2661.170 15.680 2661.490 15.740 ;
      LAYER via ;
        RECT 2409.120 207.100 2409.380 207.360 ;
        RECT 2414.640 207.100 2414.900 207.360 ;
        RECT 2414.640 15.680 2414.900 15.940 ;
        RECT 2661.200 15.680 2661.460 15.940 ;
      LAYER met2 ;
        RECT 2409.160 220.000 2409.440 224.000 ;
        RECT 2409.180 207.390 2409.320 220.000 ;
        RECT 2409.120 207.070 2409.380 207.390 ;
        RECT 2414.640 207.070 2414.900 207.390 ;
        RECT 2414.700 15.970 2414.840 207.070 ;
        RECT 2414.640 15.650 2414.900 15.970 ;
        RECT 2661.200 15.650 2661.460 15.970 ;
        RECT 2661.260 2.400 2661.400 15.650 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2423.810 210.360 2424.130 210.420 ;
        RECT 2677.270 210.360 2677.590 210.420 ;
        RECT 2423.810 210.220 2677.590 210.360 ;
        RECT 2423.810 210.160 2424.130 210.220 ;
        RECT 2677.270 210.160 2677.590 210.220 ;
      LAYER via ;
        RECT 2423.840 210.160 2424.100 210.420 ;
        RECT 2677.300 210.160 2677.560 210.420 ;
      LAYER met2 ;
        RECT 2423.880 220.000 2424.160 224.000 ;
        RECT 2423.900 210.450 2424.040 220.000 ;
        RECT 2423.840 210.130 2424.100 210.450 ;
        RECT 2677.300 210.130 2677.560 210.450 ;
        RECT 2677.360 3.130 2677.500 210.130 ;
        RECT 2677.360 2.990 2678.880 3.130 ;
        RECT 2678.740 2.400 2678.880 2.990 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2442.210 16.220 2442.530 16.280 ;
        RECT 2696.590 16.220 2696.910 16.280 ;
        RECT 2442.210 16.080 2696.910 16.220 ;
        RECT 2442.210 16.020 2442.530 16.080 ;
        RECT 2696.590 16.020 2696.910 16.080 ;
      LAYER via ;
        RECT 2442.240 16.020 2442.500 16.280 ;
        RECT 2696.620 16.020 2696.880 16.280 ;
      LAYER met2 ;
        RECT 2438.600 220.730 2438.880 224.000 ;
        RECT 2438.600 220.590 2442.440 220.730 ;
        RECT 2438.600 220.000 2438.880 220.590 ;
        RECT 2442.300 16.310 2442.440 220.590 ;
        RECT 2442.240 15.990 2442.500 16.310 ;
        RECT 2696.620 15.990 2696.880 16.310 ;
        RECT 2696.680 2.400 2696.820 15.990 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2453.250 210.700 2453.570 210.760 ;
        RECT 2701.190 210.700 2701.510 210.760 ;
        RECT 2453.250 210.560 2701.510 210.700 ;
        RECT 2453.250 210.500 2453.570 210.560 ;
        RECT 2701.190 210.500 2701.510 210.560 ;
        RECT 2701.190 16.900 2701.510 16.960 ;
        RECT 2714.530 16.900 2714.850 16.960 ;
        RECT 2701.190 16.760 2714.850 16.900 ;
        RECT 2701.190 16.700 2701.510 16.760 ;
        RECT 2714.530 16.700 2714.850 16.760 ;
      LAYER via ;
        RECT 2453.280 210.500 2453.540 210.760 ;
        RECT 2701.220 210.500 2701.480 210.760 ;
        RECT 2701.220 16.700 2701.480 16.960 ;
        RECT 2714.560 16.700 2714.820 16.960 ;
      LAYER met2 ;
        RECT 2453.320 220.000 2453.600 224.000 ;
        RECT 2453.340 210.790 2453.480 220.000 ;
        RECT 2453.280 210.470 2453.540 210.790 ;
        RECT 2701.220 210.470 2701.480 210.790 ;
        RECT 2701.280 16.990 2701.420 210.470 ;
        RECT 2701.220 16.670 2701.480 16.990 ;
        RECT 2714.560 16.670 2714.820 16.990 ;
        RECT 2714.620 2.400 2714.760 16.670 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2469.810 19.960 2470.130 20.020 ;
        RECT 2732.470 19.960 2732.790 20.020 ;
        RECT 2469.810 19.820 2732.790 19.960 ;
        RECT 2469.810 19.760 2470.130 19.820 ;
        RECT 2732.470 19.760 2732.790 19.820 ;
      LAYER via ;
        RECT 2469.840 19.760 2470.100 20.020 ;
        RECT 2732.500 19.760 2732.760 20.020 ;
      LAYER met2 ;
        RECT 2467.580 220.730 2467.860 224.000 ;
        RECT 2467.580 220.590 2470.040 220.730 ;
        RECT 2467.580 220.000 2467.860 220.590 ;
        RECT 2469.900 20.050 2470.040 220.590 ;
        RECT 2469.840 19.730 2470.100 20.050 ;
        RECT 2732.500 19.730 2732.760 20.050 ;
        RECT 2732.560 2.400 2732.700 19.730 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2714.145 13.685 2714.315 14.875 ;
      LAYER mcon ;
        RECT 2714.145 14.705 2714.315 14.875 ;
      LAYER met1 ;
        RECT 2482.230 213.080 2482.550 213.140 ;
        RECT 2708.090 213.080 2708.410 213.140 ;
        RECT 2482.230 212.940 2708.410 213.080 ;
        RECT 2482.230 212.880 2482.550 212.940 ;
        RECT 2708.090 212.880 2708.410 212.940 ;
        RECT 2708.090 14.860 2708.410 14.920 ;
        RECT 2714.085 14.860 2714.375 14.905 ;
        RECT 2708.090 14.720 2714.375 14.860 ;
        RECT 2708.090 14.660 2708.410 14.720 ;
        RECT 2714.085 14.675 2714.375 14.720 ;
        RECT 2750.410 14.180 2750.730 14.240 ;
        RECT 2715.540 14.040 2750.730 14.180 ;
        RECT 2714.085 13.840 2714.375 13.885 ;
        RECT 2715.540 13.840 2715.680 14.040 ;
        RECT 2750.410 13.980 2750.730 14.040 ;
        RECT 2714.085 13.700 2715.680 13.840 ;
        RECT 2714.085 13.655 2714.375 13.700 ;
      LAYER via ;
        RECT 2482.260 212.880 2482.520 213.140 ;
        RECT 2708.120 212.880 2708.380 213.140 ;
        RECT 2708.120 14.660 2708.380 14.920 ;
        RECT 2750.440 13.980 2750.700 14.240 ;
      LAYER met2 ;
        RECT 2482.300 220.000 2482.580 224.000 ;
        RECT 2482.320 213.170 2482.460 220.000 ;
        RECT 2482.260 212.850 2482.520 213.170 ;
        RECT 2708.120 212.850 2708.380 213.170 ;
        RECT 2708.180 14.950 2708.320 212.850 ;
        RECT 2708.120 14.630 2708.380 14.950 ;
        RECT 2750.440 13.950 2750.700 14.270 ;
        RECT 2750.500 2.400 2750.640 13.950 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2530.605 18.785 2531.695 18.955 ;
      LAYER mcon ;
        RECT 2531.525 18.785 2531.695 18.955 ;
      LAYER met1 ;
        RECT 2496.950 18.940 2497.270 19.000 ;
        RECT 2530.545 18.940 2530.835 18.985 ;
        RECT 2496.950 18.800 2530.835 18.940 ;
        RECT 2496.950 18.740 2497.270 18.800 ;
        RECT 2530.545 18.755 2530.835 18.800 ;
        RECT 2531.465 18.940 2531.755 18.985 ;
        RECT 2767.890 18.940 2768.210 19.000 ;
        RECT 2531.465 18.800 2768.210 18.940 ;
        RECT 2531.465 18.755 2531.755 18.800 ;
        RECT 2767.890 18.740 2768.210 18.800 ;
      LAYER via ;
        RECT 2496.980 18.740 2497.240 19.000 ;
        RECT 2767.920 18.740 2768.180 19.000 ;
      LAYER met2 ;
        RECT 2497.020 220.000 2497.300 224.000 ;
        RECT 2497.040 19.030 2497.180 220.000 ;
        RECT 2496.980 18.710 2497.240 19.030 ;
        RECT 2767.920 18.710 2768.180 19.030 ;
        RECT 2767.980 2.400 2768.120 18.710 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 840.950 211.040 841.270 211.100 ;
        RECT 910.410 211.040 910.730 211.100 ;
        RECT 840.950 210.900 910.730 211.040 ;
        RECT 840.950 210.840 841.270 210.900 ;
        RECT 910.410 210.840 910.730 210.900 ;
      LAYER via ;
        RECT 840.980 210.840 841.240 211.100 ;
        RECT 910.440 210.840 910.700 211.100 ;
      LAYER met2 ;
        RECT 910.480 220.000 910.760 224.000 ;
        RECT 910.500 211.130 910.640 220.000 ;
        RECT 840.980 210.810 841.240 211.130 ;
        RECT 910.440 210.810 910.700 211.130 ;
        RECT 841.040 2.400 841.180 210.810 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2511.670 213.760 2511.990 213.820 ;
        RECT 2714.990 213.760 2715.310 213.820 ;
        RECT 2511.670 213.620 2715.310 213.760 ;
        RECT 2511.670 213.560 2511.990 213.620 ;
        RECT 2714.990 213.560 2715.310 213.620 ;
        RECT 2715.910 14.520 2716.230 14.580 ;
        RECT 2785.830 14.520 2786.150 14.580 ;
        RECT 2715.910 14.380 2786.150 14.520 ;
        RECT 2715.910 14.320 2716.230 14.380 ;
        RECT 2785.830 14.320 2786.150 14.380 ;
      LAYER via ;
        RECT 2511.700 213.560 2511.960 213.820 ;
        RECT 2715.020 213.560 2715.280 213.820 ;
        RECT 2715.940 14.320 2716.200 14.580 ;
        RECT 2785.860 14.320 2786.120 14.580 ;
      LAYER met2 ;
        RECT 2511.740 220.000 2512.020 224.000 ;
        RECT 2511.760 213.850 2511.900 220.000 ;
        RECT 2511.700 213.530 2511.960 213.850 ;
        RECT 2715.020 213.530 2715.280 213.850 ;
        RECT 2715.080 14.010 2715.220 213.530 ;
        RECT 2715.940 14.290 2716.200 14.610 ;
        RECT 2785.860 14.290 2786.120 14.610 ;
        RECT 2716.000 14.010 2716.140 14.290 ;
        RECT 2715.080 13.870 2716.140 14.010 ;
        RECT 2785.920 2.400 2786.060 14.290 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2526.390 207.300 2526.710 207.360 ;
        RECT 2531.910 207.300 2532.230 207.360 ;
        RECT 2526.390 207.160 2532.230 207.300 ;
        RECT 2526.390 207.100 2526.710 207.160 ;
        RECT 2531.910 207.100 2532.230 207.160 ;
        RECT 2531.910 19.280 2532.230 19.340 ;
        RECT 2803.770 19.280 2804.090 19.340 ;
        RECT 2531.910 19.140 2804.090 19.280 ;
        RECT 2531.910 19.080 2532.230 19.140 ;
        RECT 2803.770 19.080 2804.090 19.140 ;
      LAYER via ;
        RECT 2526.420 207.100 2526.680 207.360 ;
        RECT 2531.940 207.100 2532.200 207.360 ;
        RECT 2531.940 19.080 2532.200 19.340 ;
        RECT 2803.800 19.080 2804.060 19.340 ;
      LAYER met2 ;
        RECT 2526.460 220.000 2526.740 224.000 ;
        RECT 2526.480 207.390 2526.620 220.000 ;
        RECT 2526.420 207.070 2526.680 207.390 ;
        RECT 2531.940 207.070 2532.200 207.390 ;
        RECT 2532.000 19.370 2532.140 207.070 ;
        RECT 2531.940 19.050 2532.200 19.370 ;
        RECT 2803.800 19.050 2804.060 19.370 ;
        RECT 2803.860 2.400 2804.000 19.050 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2541.110 213.420 2541.430 213.480 ;
        RECT 2721.890 213.420 2722.210 213.480 ;
        RECT 2541.110 213.280 2722.210 213.420 ;
        RECT 2541.110 213.220 2541.430 213.280 ;
        RECT 2721.890 213.220 2722.210 213.280 ;
        RECT 2721.890 16.900 2722.210 16.960 ;
        RECT 2821.710 16.900 2822.030 16.960 ;
        RECT 2721.890 16.760 2822.030 16.900 ;
        RECT 2721.890 16.700 2722.210 16.760 ;
        RECT 2821.710 16.700 2822.030 16.760 ;
      LAYER via ;
        RECT 2541.140 213.220 2541.400 213.480 ;
        RECT 2721.920 213.220 2722.180 213.480 ;
        RECT 2721.920 16.700 2722.180 16.960 ;
        RECT 2821.740 16.700 2822.000 16.960 ;
      LAYER met2 ;
        RECT 2541.180 220.000 2541.460 224.000 ;
        RECT 2541.200 213.510 2541.340 220.000 ;
        RECT 2541.140 213.190 2541.400 213.510 ;
        RECT 2721.920 213.190 2722.180 213.510 ;
        RECT 2721.980 16.990 2722.120 213.190 ;
        RECT 2721.920 16.670 2722.180 16.990 ;
        RECT 2821.740 16.670 2822.000 16.990 ;
        RECT 2821.800 2.400 2821.940 16.670 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2555.830 207.300 2556.150 207.360 ;
        RECT 2559.510 207.300 2559.830 207.360 ;
        RECT 2555.830 207.160 2559.830 207.300 ;
        RECT 2555.830 207.100 2556.150 207.160 ;
        RECT 2559.510 207.100 2559.830 207.160 ;
        RECT 2559.510 18.600 2559.830 18.660 ;
        RECT 2559.510 18.460 2590.560 18.600 ;
        RECT 2559.510 18.400 2559.830 18.460 ;
        RECT 2590.420 18.260 2590.560 18.460 ;
        RECT 2839.190 18.260 2839.510 18.320 ;
        RECT 2590.420 18.120 2839.510 18.260 ;
        RECT 2839.190 18.060 2839.510 18.120 ;
      LAYER via ;
        RECT 2555.860 207.100 2556.120 207.360 ;
        RECT 2559.540 207.100 2559.800 207.360 ;
        RECT 2559.540 18.400 2559.800 18.660 ;
        RECT 2839.220 18.060 2839.480 18.320 ;
      LAYER met2 ;
        RECT 2555.900 220.000 2556.180 224.000 ;
        RECT 2555.920 207.390 2556.060 220.000 ;
        RECT 2555.860 207.070 2556.120 207.390 ;
        RECT 2559.540 207.070 2559.800 207.390 ;
        RECT 2559.600 18.690 2559.740 207.070 ;
        RECT 2559.540 18.370 2559.800 18.690 ;
        RECT 2839.220 18.030 2839.480 18.350 ;
        RECT 2839.280 2.400 2839.420 18.030 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2570.550 212.400 2570.870 212.460 ;
        RECT 2728.790 212.400 2729.110 212.460 ;
        RECT 2570.550 212.260 2729.110 212.400 ;
        RECT 2570.550 212.200 2570.870 212.260 ;
        RECT 2728.790 212.200 2729.110 212.260 ;
        RECT 2728.790 20.300 2729.110 20.360 ;
        RECT 2857.130 20.300 2857.450 20.360 ;
        RECT 2728.790 20.160 2857.450 20.300 ;
        RECT 2728.790 20.100 2729.110 20.160 ;
        RECT 2857.130 20.100 2857.450 20.160 ;
      LAYER via ;
        RECT 2570.580 212.200 2570.840 212.460 ;
        RECT 2728.820 212.200 2729.080 212.460 ;
        RECT 2728.820 20.100 2729.080 20.360 ;
        RECT 2857.160 20.100 2857.420 20.360 ;
      LAYER met2 ;
        RECT 2570.620 220.000 2570.900 224.000 ;
        RECT 2570.640 212.490 2570.780 220.000 ;
        RECT 2570.580 212.170 2570.840 212.490 ;
        RECT 2728.820 212.170 2729.080 212.490 ;
        RECT 2728.880 20.390 2729.020 212.170 ;
        RECT 2728.820 20.070 2729.080 20.390 ;
        RECT 2857.160 20.070 2857.420 20.390 ;
        RECT 2857.220 2.400 2857.360 20.070 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2587.110 17.580 2587.430 17.640 ;
        RECT 2875.070 17.580 2875.390 17.640 ;
        RECT 2587.110 17.440 2875.390 17.580 ;
        RECT 2587.110 17.380 2587.430 17.440 ;
        RECT 2875.070 17.380 2875.390 17.440 ;
      LAYER via ;
        RECT 2587.140 17.380 2587.400 17.640 ;
        RECT 2875.100 17.380 2875.360 17.640 ;
      LAYER met2 ;
        RECT 2585.340 220.730 2585.620 224.000 ;
        RECT 2585.340 220.590 2587.340 220.730 ;
        RECT 2585.340 220.000 2585.620 220.590 ;
        RECT 2587.200 17.670 2587.340 220.590 ;
        RECT 2587.140 17.350 2587.400 17.670 ;
        RECT 2875.100 17.350 2875.360 17.670 ;
        RECT 2875.160 2.400 2875.300 17.350 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2599.990 210.020 2600.310 210.080 ;
        RECT 2735.690 210.020 2736.010 210.080 ;
        RECT 2599.990 209.880 2736.010 210.020 ;
        RECT 2599.990 209.820 2600.310 209.880 ;
        RECT 2735.690 209.820 2736.010 209.880 ;
        RECT 2735.690 19.960 2736.010 20.020 ;
        RECT 2893.010 19.960 2893.330 20.020 ;
        RECT 2735.690 19.820 2893.330 19.960 ;
        RECT 2735.690 19.760 2736.010 19.820 ;
        RECT 2893.010 19.760 2893.330 19.820 ;
      LAYER via ;
        RECT 2600.020 209.820 2600.280 210.080 ;
        RECT 2735.720 209.820 2735.980 210.080 ;
        RECT 2735.720 19.760 2735.980 20.020 ;
        RECT 2893.040 19.760 2893.300 20.020 ;
      LAYER met2 ;
        RECT 2600.060 220.000 2600.340 224.000 ;
        RECT 2600.080 210.110 2600.220 220.000 ;
        RECT 2600.020 209.790 2600.280 210.110 ;
        RECT 2735.720 209.790 2735.980 210.110 ;
        RECT 2735.780 20.050 2735.920 209.790 ;
        RECT 2735.720 19.730 2735.980 20.050 ;
        RECT 2893.040 19.730 2893.300 20.050 ;
        RECT 2893.100 2.400 2893.240 19.730 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2614.710 211.720 2615.030 211.780 ;
        RECT 2736.150 211.720 2736.470 211.780 ;
        RECT 2614.710 211.580 2736.470 211.720 ;
        RECT 2614.710 211.520 2615.030 211.580 ;
        RECT 2736.150 211.520 2736.470 211.580 ;
      LAYER via ;
        RECT 2614.740 211.520 2615.000 211.780 ;
        RECT 2736.180 211.520 2736.440 211.780 ;
      LAYER met2 ;
        RECT 2614.780 220.000 2615.060 224.000 ;
        RECT 2614.800 211.810 2614.940 220.000 ;
        RECT 2614.740 211.490 2615.000 211.810 ;
        RECT 2736.180 211.490 2736.440 211.810 ;
        RECT 2736.240 16.845 2736.380 211.490 ;
        RECT 2736.170 16.475 2736.450 16.845 ;
        RECT 2910.970 16.475 2911.250 16.845 ;
        RECT 2911.040 2.400 2911.180 16.475 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
      LAYER via2 ;
        RECT 2736.170 16.520 2736.450 16.800 ;
        RECT 2910.970 16.520 2911.250 16.800 ;
      LAYER met3 ;
        RECT 2736.145 16.810 2736.475 16.825 ;
        RECT 2910.945 16.810 2911.275 16.825 ;
        RECT 2736.145 16.510 2911.275 16.810 ;
        RECT 2736.145 16.495 2736.475 16.510 ;
        RECT 2910.945 16.495 2911.275 16.510 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 862.110 213.080 862.430 213.140 ;
        RECT 925.130 213.080 925.450 213.140 ;
        RECT 862.110 212.940 925.450 213.080 ;
        RECT 862.110 212.880 862.430 212.940 ;
        RECT 925.130 212.880 925.450 212.940 ;
        RECT 858.890 20.640 859.210 20.700 ;
        RECT 862.110 20.640 862.430 20.700 ;
        RECT 858.890 20.500 862.430 20.640 ;
        RECT 858.890 20.440 859.210 20.500 ;
        RECT 862.110 20.440 862.430 20.500 ;
      LAYER via ;
        RECT 862.140 212.880 862.400 213.140 ;
        RECT 925.160 212.880 925.420 213.140 ;
        RECT 858.920 20.440 859.180 20.700 ;
        RECT 862.140 20.440 862.400 20.700 ;
      LAYER met2 ;
        RECT 925.200 220.000 925.480 224.000 ;
        RECT 925.220 213.170 925.360 220.000 ;
        RECT 862.140 212.850 862.400 213.170 ;
        RECT 925.160 212.850 925.420 213.170 ;
        RECT 862.200 20.730 862.340 212.850 ;
        RECT 858.920 20.410 859.180 20.730 ;
        RECT 862.140 20.410 862.400 20.730 ;
        RECT 858.980 2.400 859.120 20.410 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.350 212.060 882.670 212.120 ;
        RECT 939.850 212.060 940.170 212.120 ;
        RECT 882.350 211.920 940.170 212.060 ;
        RECT 882.350 211.860 882.670 211.920 ;
        RECT 939.850 211.860 940.170 211.920 ;
        RECT 876.830 16.560 877.150 16.620 ;
        RECT 882.350 16.560 882.670 16.620 ;
        RECT 876.830 16.420 882.670 16.560 ;
        RECT 876.830 16.360 877.150 16.420 ;
        RECT 882.350 16.360 882.670 16.420 ;
      LAYER via ;
        RECT 882.380 211.860 882.640 212.120 ;
        RECT 939.880 211.860 940.140 212.120 ;
        RECT 876.860 16.360 877.120 16.620 ;
        RECT 882.380 16.360 882.640 16.620 ;
      LAYER met2 ;
        RECT 939.920 220.000 940.200 224.000 ;
        RECT 939.940 212.150 940.080 220.000 ;
        RECT 882.380 211.830 882.640 212.150 ;
        RECT 939.880 211.830 940.140 212.150 ;
        RECT 882.440 16.650 882.580 211.830 ;
        RECT 876.860 16.330 877.120 16.650 ;
        RECT 882.380 16.330 882.640 16.650 ;
        RECT 876.920 2.400 877.060 16.330 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 896.610 210.700 896.930 210.760 ;
        RECT 954.570 210.700 954.890 210.760 ;
        RECT 896.610 210.560 954.890 210.700 ;
        RECT 896.610 210.500 896.930 210.560 ;
        RECT 954.570 210.500 954.890 210.560 ;
      LAYER via ;
        RECT 896.640 210.500 896.900 210.760 ;
        RECT 954.600 210.500 954.860 210.760 ;
      LAYER met2 ;
        RECT 954.640 220.000 954.920 224.000 ;
        RECT 954.660 210.790 954.800 220.000 ;
        RECT 896.640 210.470 896.900 210.790 ;
        RECT 954.600 210.470 954.860 210.790 ;
        RECT 896.700 17.410 896.840 210.470 ;
        RECT 894.860 17.270 896.840 17.410 ;
        RECT 894.860 2.400 895.000 17.270 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 917.310 213.420 917.630 213.480 ;
        RECT 968.830 213.420 969.150 213.480 ;
        RECT 917.310 213.280 969.150 213.420 ;
        RECT 917.310 213.220 917.630 213.280 ;
        RECT 968.830 213.220 969.150 213.280 ;
        RECT 912.710 17.580 913.030 17.640 ;
        RECT 917.310 17.580 917.630 17.640 ;
        RECT 912.710 17.440 917.630 17.580 ;
        RECT 912.710 17.380 913.030 17.440 ;
        RECT 917.310 17.380 917.630 17.440 ;
      LAYER via ;
        RECT 917.340 213.220 917.600 213.480 ;
        RECT 968.860 213.220 969.120 213.480 ;
        RECT 912.740 17.380 913.000 17.640 ;
        RECT 917.340 17.380 917.600 17.640 ;
      LAYER met2 ;
        RECT 968.900 220.000 969.180 224.000 ;
        RECT 968.920 213.510 969.060 220.000 ;
        RECT 917.340 213.190 917.600 213.510 ;
        RECT 968.860 213.190 969.120 213.510 ;
        RECT 917.400 17.670 917.540 213.190 ;
        RECT 912.740 17.350 913.000 17.670 ;
        RECT 917.340 17.350 917.600 17.670 ;
        RECT 912.800 2.400 912.940 17.350 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 931.110 213.080 931.430 213.140 ;
        RECT 983.550 213.080 983.870 213.140 ;
        RECT 931.110 212.940 983.870 213.080 ;
        RECT 931.110 212.880 931.430 212.940 ;
        RECT 983.550 212.880 983.870 212.940 ;
      LAYER via ;
        RECT 931.140 212.880 931.400 213.140 ;
        RECT 983.580 212.880 983.840 213.140 ;
      LAYER met2 ;
        RECT 983.620 220.000 983.900 224.000 ;
        RECT 983.640 213.170 983.780 220.000 ;
        RECT 931.140 212.850 931.400 213.170 ;
        RECT 983.580 212.850 983.840 213.170 ;
        RECT 931.200 17.410 931.340 212.850 ;
        RECT 930.280 17.270 931.340 17.410 ;
        RECT 930.280 2.400 930.420 17.270 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 951.810 213.760 952.130 213.820 ;
        RECT 998.270 213.760 998.590 213.820 ;
        RECT 951.810 213.620 998.590 213.760 ;
        RECT 951.810 213.560 952.130 213.620 ;
        RECT 998.270 213.560 998.590 213.620 ;
        RECT 948.130 17.580 948.450 17.640 ;
        RECT 951.810 17.580 952.130 17.640 ;
        RECT 948.130 17.440 952.130 17.580 ;
        RECT 948.130 17.380 948.450 17.440 ;
        RECT 951.810 17.380 952.130 17.440 ;
      LAYER via ;
        RECT 951.840 213.560 952.100 213.820 ;
        RECT 998.300 213.560 998.560 213.820 ;
        RECT 948.160 17.380 948.420 17.640 ;
        RECT 951.840 17.380 952.100 17.640 ;
      LAYER met2 ;
        RECT 998.340 220.000 998.620 224.000 ;
        RECT 998.360 213.850 998.500 220.000 ;
        RECT 951.840 213.530 952.100 213.850 ;
        RECT 998.300 213.530 998.560 213.850 ;
        RECT 951.900 17.670 952.040 213.530 ;
        RECT 948.160 17.350 948.420 17.670 ;
        RECT 951.840 17.350 952.100 17.670 ;
        RECT 948.220 2.400 948.360 17.350 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.510 207.300 972.830 207.360 ;
        RECT 1012.990 207.300 1013.310 207.360 ;
        RECT 972.510 207.160 1013.310 207.300 ;
        RECT 972.510 207.100 972.830 207.160 ;
        RECT 1012.990 207.100 1013.310 207.160 ;
        RECT 966.070 17.580 966.390 17.640 ;
        RECT 972.510 17.580 972.830 17.640 ;
        RECT 966.070 17.440 972.830 17.580 ;
        RECT 966.070 17.380 966.390 17.440 ;
        RECT 972.510 17.380 972.830 17.440 ;
      LAYER via ;
        RECT 972.540 207.100 972.800 207.360 ;
        RECT 1013.020 207.100 1013.280 207.360 ;
        RECT 966.100 17.380 966.360 17.640 ;
        RECT 972.540 17.380 972.800 17.640 ;
      LAYER met2 ;
        RECT 1013.060 220.000 1013.340 224.000 ;
        RECT 1013.080 207.390 1013.220 220.000 ;
        RECT 972.540 207.070 972.800 207.390 ;
        RECT 1013.020 207.070 1013.280 207.390 ;
        RECT 972.600 17.670 972.740 207.070 ;
        RECT 966.100 17.350 966.360 17.670 ;
        RECT 972.540 17.350 972.800 17.670 ;
        RECT 966.160 2.400 966.300 17.350 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 986.310 213.080 986.630 213.140 ;
        RECT 1027.710 213.080 1028.030 213.140 ;
        RECT 986.310 212.940 1028.030 213.080 ;
        RECT 986.310 212.880 986.630 212.940 ;
        RECT 1027.710 212.880 1028.030 212.940 ;
        RECT 984.010 17.580 984.330 17.640 ;
        RECT 986.310 17.580 986.630 17.640 ;
        RECT 984.010 17.440 986.630 17.580 ;
        RECT 984.010 17.380 984.330 17.440 ;
        RECT 986.310 17.380 986.630 17.440 ;
      LAYER via ;
        RECT 986.340 212.880 986.600 213.140 ;
        RECT 1027.740 212.880 1028.000 213.140 ;
        RECT 984.040 17.380 984.300 17.640 ;
        RECT 986.340 17.380 986.600 17.640 ;
      LAYER met2 ;
        RECT 1027.780 220.000 1028.060 224.000 ;
        RECT 1027.800 213.170 1027.940 220.000 ;
        RECT 986.340 212.850 986.600 213.170 ;
        RECT 1027.740 212.850 1028.000 213.170 ;
        RECT 986.400 17.670 986.540 212.850 ;
        RECT 984.040 17.350 984.300 17.670 ;
        RECT 986.340 17.350 986.600 17.670 ;
        RECT 984.100 2.400 984.240 17.350 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.450 210.020 668.770 210.080 ;
        RECT 763.210 210.020 763.530 210.080 ;
        RECT 668.450 209.880 763.530 210.020 ;
        RECT 668.450 209.820 668.770 209.880 ;
        RECT 763.210 209.820 763.530 209.880 ;
        RECT 662.930 17.580 663.250 17.640 ;
        RECT 668.450 17.580 668.770 17.640 ;
        RECT 662.930 17.440 668.770 17.580 ;
        RECT 662.930 17.380 663.250 17.440 ;
        RECT 668.450 17.380 668.770 17.440 ;
      LAYER via ;
        RECT 668.480 209.820 668.740 210.080 ;
        RECT 763.240 209.820 763.500 210.080 ;
        RECT 662.960 17.380 663.220 17.640 ;
        RECT 668.480 17.380 668.740 17.640 ;
      LAYER met2 ;
        RECT 763.280 220.000 763.560 224.000 ;
        RECT 763.300 210.110 763.440 220.000 ;
        RECT 668.480 209.790 668.740 210.110 ;
        RECT 763.240 209.790 763.500 210.110 ;
        RECT 668.540 17.670 668.680 209.790 ;
        RECT 662.960 17.350 663.220 17.670 ;
        RECT 668.480 17.350 668.740 17.670 ;
        RECT 663.020 2.400 663.160 17.350 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.010 208.320 1007.330 208.380 ;
        RECT 1042.430 208.320 1042.750 208.380 ;
        RECT 1007.010 208.180 1042.750 208.320 ;
        RECT 1007.010 208.120 1007.330 208.180 ;
        RECT 1042.430 208.120 1042.750 208.180 ;
        RECT 1001.950 17.580 1002.270 17.640 ;
        RECT 1007.010 17.580 1007.330 17.640 ;
        RECT 1001.950 17.440 1007.330 17.580 ;
        RECT 1001.950 17.380 1002.270 17.440 ;
        RECT 1007.010 17.380 1007.330 17.440 ;
      LAYER via ;
        RECT 1007.040 208.120 1007.300 208.380 ;
        RECT 1042.460 208.120 1042.720 208.380 ;
        RECT 1001.980 17.380 1002.240 17.640 ;
        RECT 1007.040 17.380 1007.300 17.640 ;
      LAYER met2 ;
        RECT 1042.500 220.000 1042.780 224.000 ;
        RECT 1042.520 208.410 1042.660 220.000 ;
        RECT 1007.040 208.090 1007.300 208.410 ;
        RECT 1042.460 208.090 1042.720 208.410 ;
        RECT 1007.100 17.670 1007.240 208.090 ;
        RECT 1001.980 17.350 1002.240 17.670 ;
        RECT 1007.040 17.350 1007.300 17.670 ;
        RECT 1002.040 2.400 1002.180 17.350 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1020.810 207.640 1021.130 207.700 ;
        RECT 1057.150 207.640 1057.470 207.700 ;
        RECT 1020.810 207.500 1057.470 207.640 ;
        RECT 1020.810 207.440 1021.130 207.500 ;
        RECT 1057.150 207.440 1057.470 207.500 ;
      LAYER via ;
        RECT 1020.840 207.440 1021.100 207.700 ;
        RECT 1057.180 207.440 1057.440 207.700 ;
      LAYER met2 ;
        RECT 1057.220 220.000 1057.500 224.000 ;
        RECT 1057.240 207.730 1057.380 220.000 ;
        RECT 1020.840 207.410 1021.100 207.730 ;
        RECT 1057.180 207.410 1057.440 207.730 ;
        RECT 1020.900 17.410 1021.040 207.410 ;
        RECT 1019.520 17.270 1021.040 17.410 ;
        RECT 1019.520 2.400 1019.660 17.270 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1041.510 211.720 1041.830 211.780 ;
        RECT 1071.870 211.720 1072.190 211.780 ;
        RECT 1041.510 211.580 1072.190 211.720 ;
        RECT 1041.510 211.520 1041.830 211.580 ;
        RECT 1071.870 211.520 1072.190 211.580 ;
        RECT 1037.370 17.580 1037.690 17.640 ;
        RECT 1041.510 17.580 1041.830 17.640 ;
        RECT 1037.370 17.440 1041.830 17.580 ;
        RECT 1037.370 17.380 1037.690 17.440 ;
        RECT 1041.510 17.380 1041.830 17.440 ;
      LAYER via ;
        RECT 1041.540 211.520 1041.800 211.780 ;
        RECT 1071.900 211.520 1072.160 211.780 ;
        RECT 1037.400 17.380 1037.660 17.640 ;
        RECT 1041.540 17.380 1041.800 17.640 ;
      LAYER met2 ;
        RECT 1071.940 220.000 1072.220 224.000 ;
        RECT 1071.960 211.810 1072.100 220.000 ;
        RECT 1041.540 211.490 1041.800 211.810 ;
        RECT 1071.900 211.490 1072.160 211.810 ;
        RECT 1041.600 17.670 1041.740 211.490 ;
        RECT 1037.400 17.350 1037.660 17.670 ;
        RECT 1041.540 17.350 1041.800 17.670 ;
        RECT 1037.460 2.400 1037.600 17.350 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1055.310 208.660 1055.630 208.720 ;
        RECT 1086.590 208.660 1086.910 208.720 ;
        RECT 1055.310 208.520 1086.910 208.660 ;
        RECT 1055.310 208.460 1055.630 208.520 ;
        RECT 1086.590 208.460 1086.910 208.520 ;
      LAYER via ;
        RECT 1055.340 208.460 1055.600 208.720 ;
        RECT 1086.620 208.460 1086.880 208.720 ;
      LAYER met2 ;
        RECT 1086.660 220.000 1086.940 224.000 ;
        RECT 1086.680 208.750 1086.820 220.000 ;
        RECT 1055.340 208.430 1055.600 208.750 ;
        RECT 1086.620 208.430 1086.880 208.750 ;
        RECT 1055.400 2.400 1055.540 208.430 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1076.010 207.640 1076.330 207.700 ;
        RECT 1101.310 207.640 1101.630 207.700 ;
        RECT 1076.010 207.500 1101.630 207.640 ;
        RECT 1076.010 207.440 1076.330 207.500 ;
        RECT 1101.310 207.440 1101.630 207.500 ;
        RECT 1073.250 17.580 1073.570 17.640 ;
        RECT 1076.010 17.580 1076.330 17.640 ;
        RECT 1073.250 17.440 1076.330 17.580 ;
        RECT 1073.250 17.380 1073.570 17.440 ;
        RECT 1076.010 17.380 1076.330 17.440 ;
      LAYER via ;
        RECT 1076.040 207.440 1076.300 207.700 ;
        RECT 1101.340 207.440 1101.600 207.700 ;
        RECT 1073.280 17.380 1073.540 17.640 ;
        RECT 1076.040 17.380 1076.300 17.640 ;
      LAYER met2 ;
        RECT 1101.380 220.000 1101.660 224.000 ;
        RECT 1101.400 207.730 1101.540 220.000 ;
        RECT 1076.040 207.410 1076.300 207.730 ;
        RECT 1101.340 207.410 1101.600 207.730 ;
        RECT 1076.100 17.670 1076.240 207.410 ;
        RECT 1073.280 17.350 1073.540 17.670 ;
        RECT 1076.040 17.350 1076.300 17.670 ;
        RECT 1073.340 2.400 1073.480 17.350 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.710 212.060 1097.030 212.120 ;
        RECT 1116.030 212.060 1116.350 212.120 ;
        RECT 1096.710 211.920 1116.350 212.060 ;
        RECT 1096.710 211.860 1097.030 211.920 ;
        RECT 1116.030 211.860 1116.350 211.920 ;
        RECT 1090.730 15.200 1091.050 15.260 ;
        RECT 1096.710 15.200 1097.030 15.260 ;
        RECT 1090.730 15.060 1097.030 15.200 ;
        RECT 1090.730 15.000 1091.050 15.060 ;
        RECT 1096.710 15.000 1097.030 15.060 ;
      LAYER via ;
        RECT 1096.740 211.860 1097.000 212.120 ;
        RECT 1116.060 211.860 1116.320 212.120 ;
        RECT 1090.760 15.000 1091.020 15.260 ;
        RECT 1096.740 15.000 1097.000 15.260 ;
      LAYER met2 ;
        RECT 1116.100 220.000 1116.380 224.000 ;
        RECT 1116.120 212.150 1116.260 220.000 ;
        RECT 1096.740 211.830 1097.000 212.150 ;
        RECT 1116.060 211.830 1116.320 212.150 ;
        RECT 1096.800 15.290 1096.940 211.830 ;
        RECT 1090.760 14.970 1091.020 15.290 ;
        RECT 1096.740 14.970 1097.000 15.290 ;
        RECT 1090.820 2.400 1090.960 14.970 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1110.510 207.640 1110.830 207.700 ;
        RECT 1130.750 207.640 1131.070 207.700 ;
        RECT 1110.510 207.500 1131.070 207.640 ;
        RECT 1110.510 207.440 1110.830 207.500 ;
        RECT 1130.750 207.440 1131.070 207.500 ;
      LAYER via ;
        RECT 1110.540 207.440 1110.800 207.700 ;
        RECT 1130.780 207.440 1131.040 207.700 ;
      LAYER met2 ;
        RECT 1130.820 220.000 1131.100 224.000 ;
        RECT 1130.840 207.730 1130.980 220.000 ;
        RECT 1110.540 207.410 1110.800 207.730 ;
        RECT 1130.780 207.410 1131.040 207.730 ;
        RECT 1110.600 17.410 1110.740 207.410 ;
        RECT 1108.760 17.270 1110.740 17.410 ;
        RECT 1108.760 2.400 1108.900 17.270 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1131.210 207.640 1131.530 207.700 ;
        RECT 1145.470 207.640 1145.790 207.700 ;
        RECT 1131.210 207.500 1145.790 207.640 ;
        RECT 1131.210 207.440 1131.530 207.500 ;
        RECT 1145.470 207.440 1145.790 207.500 ;
        RECT 1126.610 17.580 1126.930 17.640 ;
        RECT 1131.210 17.580 1131.530 17.640 ;
        RECT 1126.610 17.440 1131.530 17.580 ;
        RECT 1126.610 17.380 1126.930 17.440 ;
        RECT 1131.210 17.380 1131.530 17.440 ;
      LAYER via ;
        RECT 1131.240 207.440 1131.500 207.700 ;
        RECT 1145.500 207.440 1145.760 207.700 ;
        RECT 1126.640 17.380 1126.900 17.640 ;
        RECT 1131.240 17.380 1131.500 17.640 ;
      LAYER met2 ;
        RECT 1145.540 220.000 1145.820 224.000 ;
        RECT 1145.560 207.730 1145.700 220.000 ;
        RECT 1131.240 207.410 1131.500 207.730 ;
        RECT 1145.500 207.410 1145.760 207.730 ;
        RECT 1131.300 17.670 1131.440 207.410 ;
        RECT 1126.640 17.350 1126.900 17.670 ;
        RECT 1131.240 17.350 1131.500 17.670 ;
        RECT 1126.700 2.400 1126.840 17.350 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1145.010 210.360 1145.330 210.420 ;
        RECT 1160.190 210.360 1160.510 210.420 ;
        RECT 1145.010 210.220 1160.510 210.360 ;
        RECT 1145.010 210.160 1145.330 210.220 ;
        RECT 1160.190 210.160 1160.510 210.220 ;
      LAYER via ;
        RECT 1145.040 210.160 1145.300 210.420 ;
        RECT 1160.220 210.160 1160.480 210.420 ;
      LAYER met2 ;
        RECT 1160.260 220.000 1160.540 224.000 ;
        RECT 1160.280 210.450 1160.420 220.000 ;
        RECT 1145.040 210.130 1145.300 210.450 ;
        RECT 1160.220 210.130 1160.480 210.450 ;
        RECT 1145.100 17.410 1145.240 210.130 ;
        RECT 1144.640 17.270 1145.240 17.410 ;
        RECT 1144.640 2.400 1144.780 17.270 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1165.710 207.640 1166.030 207.700 ;
        RECT 1174.910 207.640 1175.230 207.700 ;
        RECT 1165.710 207.500 1175.230 207.640 ;
        RECT 1165.710 207.440 1166.030 207.500 ;
        RECT 1174.910 207.440 1175.230 207.500 ;
        RECT 1162.490 17.580 1162.810 17.640 ;
        RECT 1165.710 17.580 1166.030 17.640 ;
        RECT 1162.490 17.440 1166.030 17.580 ;
        RECT 1162.490 17.380 1162.810 17.440 ;
        RECT 1165.710 17.380 1166.030 17.440 ;
      LAYER via ;
        RECT 1165.740 207.440 1166.000 207.700 ;
        RECT 1174.940 207.440 1175.200 207.700 ;
        RECT 1162.520 17.380 1162.780 17.640 ;
        RECT 1165.740 17.380 1166.000 17.640 ;
      LAYER met2 ;
        RECT 1174.980 220.000 1175.260 224.000 ;
        RECT 1175.000 207.730 1175.140 220.000 ;
        RECT 1165.740 207.410 1166.000 207.730 ;
        RECT 1174.940 207.410 1175.200 207.730 ;
        RECT 1165.800 17.670 1165.940 207.410 ;
        RECT 1162.520 17.350 1162.780 17.670 ;
        RECT 1165.740 17.350 1166.000 17.670 ;
        RECT 1162.580 2.400 1162.720 17.350 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 682.710 207.300 683.030 207.360 ;
        RECT 777.930 207.300 778.250 207.360 ;
        RECT 682.710 207.160 778.250 207.300 ;
        RECT 682.710 207.100 683.030 207.160 ;
        RECT 777.930 207.100 778.250 207.160 ;
        RECT 680.410 14.520 680.730 14.580 ;
        RECT 682.710 14.520 683.030 14.580 ;
        RECT 680.410 14.380 683.030 14.520 ;
        RECT 680.410 14.320 680.730 14.380 ;
        RECT 682.710 14.320 683.030 14.380 ;
      LAYER via ;
        RECT 682.740 207.100 683.000 207.360 ;
        RECT 777.960 207.100 778.220 207.360 ;
        RECT 680.440 14.320 680.700 14.580 ;
        RECT 682.740 14.320 683.000 14.580 ;
      LAYER met2 ;
        RECT 778.000 220.000 778.280 224.000 ;
        RECT 778.020 207.390 778.160 220.000 ;
        RECT 682.740 207.070 683.000 207.390 ;
        RECT 777.960 207.070 778.220 207.390 ;
        RECT 682.800 14.610 682.940 207.070 ;
        RECT 680.440 14.290 680.700 14.610 ;
        RECT 682.740 14.290 683.000 14.610 ;
        RECT 680.500 2.400 680.640 14.290 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1179.970 17.920 1180.290 17.980 ;
        RECT 1186.870 17.920 1187.190 17.980 ;
        RECT 1179.970 17.780 1187.190 17.920 ;
        RECT 1179.970 17.720 1180.290 17.780 ;
        RECT 1186.870 17.720 1187.190 17.780 ;
      LAYER via ;
        RECT 1180.000 17.720 1180.260 17.980 ;
        RECT 1186.900 17.720 1187.160 17.980 ;
      LAYER met2 ;
        RECT 1189.700 220.730 1189.980 224.000 ;
        RECT 1186.960 220.590 1189.980 220.730 ;
        RECT 1186.960 18.010 1187.100 220.590 ;
        RECT 1189.700 220.000 1189.980 220.590 ;
        RECT 1180.000 17.690 1180.260 18.010 ;
        RECT 1186.900 17.690 1187.160 18.010 ;
        RECT 1180.060 2.400 1180.200 17.690 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1200.210 213.760 1200.530 213.820 ;
        RECT 1204.350 213.760 1204.670 213.820 ;
        RECT 1200.210 213.620 1204.670 213.760 ;
        RECT 1200.210 213.560 1200.530 213.620 ;
        RECT 1204.350 213.560 1204.670 213.620 ;
        RECT 1197.910 17.580 1198.230 17.640 ;
        RECT 1200.210 17.580 1200.530 17.640 ;
        RECT 1197.910 17.440 1200.530 17.580 ;
        RECT 1197.910 17.380 1198.230 17.440 ;
        RECT 1200.210 17.380 1200.530 17.440 ;
      LAYER via ;
        RECT 1200.240 213.560 1200.500 213.820 ;
        RECT 1204.380 213.560 1204.640 213.820 ;
        RECT 1197.940 17.380 1198.200 17.640 ;
        RECT 1200.240 17.380 1200.500 17.640 ;
      LAYER met2 ;
        RECT 1204.420 220.000 1204.700 224.000 ;
        RECT 1204.440 213.850 1204.580 220.000 ;
        RECT 1200.240 213.530 1200.500 213.850 ;
        RECT 1204.380 213.530 1204.640 213.850 ;
        RECT 1200.300 17.670 1200.440 213.530 ;
        RECT 1197.940 17.350 1198.200 17.670 ;
        RECT 1200.240 17.350 1200.500 17.670 ;
        RECT 1198.000 2.400 1198.140 17.350 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1218.680 220.730 1218.960 224.000 ;
        RECT 1214.560 220.590 1218.960 220.730 ;
        RECT 1214.560 24.210 1214.700 220.590 ;
        RECT 1218.680 220.000 1218.960 220.590 ;
        RECT 1214.560 24.070 1216.080 24.210 ;
        RECT 1215.940 2.400 1216.080 24.070 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1229.725 144.925 1229.895 193.035 ;
        RECT 1230.185 48.365 1230.355 96.475 ;
      LAYER mcon ;
        RECT 1229.725 192.865 1229.895 193.035 ;
        RECT 1230.185 96.305 1230.355 96.475 ;
      LAYER met1 ;
        RECT 1229.665 193.020 1229.955 193.065 ;
        RECT 1230.110 193.020 1230.430 193.080 ;
        RECT 1229.665 192.880 1230.430 193.020 ;
        RECT 1229.665 192.835 1229.955 192.880 ;
        RECT 1230.110 192.820 1230.430 192.880 ;
        RECT 1229.650 145.080 1229.970 145.140 ;
        RECT 1229.455 144.940 1229.970 145.080 ;
        RECT 1229.650 144.880 1229.970 144.940 ;
        RECT 1229.190 110.400 1229.510 110.460 ;
        RECT 1230.110 110.400 1230.430 110.460 ;
        RECT 1229.190 110.260 1230.430 110.400 ;
        RECT 1229.190 110.200 1229.510 110.260 ;
        RECT 1230.110 110.200 1230.430 110.260 ;
        RECT 1230.110 96.460 1230.430 96.520 ;
        RECT 1229.915 96.320 1230.430 96.460 ;
        RECT 1230.110 96.260 1230.430 96.320 ;
        RECT 1230.110 48.520 1230.430 48.580 ;
        RECT 1229.915 48.380 1230.430 48.520 ;
        RECT 1230.110 48.320 1230.430 48.380 ;
        RECT 1230.110 20.640 1230.430 20.700 ;
        RECT 1233.790 20.640 1234.110 20.700 ;
        RECT 1230.110 20.500 1234.110 20.640 ;
        RECT 1230.110 20.440 1230.430 20.500 ;
        RECT 1233.790 20.440 1234.110 20.500 ;
      LAYER via ;
        RECT 1230.140 192.820 1230.400 193.080 ;
        RECT 1229.680 144.880 1229.940 145.140 ;
        RECT 1229.220 110.200 1229.480 110.460 ;
        RECT 1230.140 110.200 1230.400 110.460 ;
        RECT 1230.140 96.260 1230.400 96.520 ;
        RECT 1230.140 48.320 1230.400 48.580 ;
        RECT 1230.140 20.440 1230.400 20.700 ;
        RECT 1233.820 20.440 1234.080 20.700 ;
      LAYER met2 ;
        RECT 1233.400 221.410 1233.680 224.000 ;
        RECT 1230.660 221.270 1233.680 221.410 ;
        RECT 1230.660 207.130 1230.800 221.270 ;
        RECT 1233.400 220.000 1233.680 221.270 ;
        RECT 1230.200 206.990 1230.800 207.130 ;
        RECT 1230.200 193.110 1230.340 206.990 ;
        RECT 1230.140 192.790 1230.400 193.110 ;
        RECT 1229.680 144.850 1229.940 145.170 ;
        RECT 1229.740 110.570 1229.880 144.850 ;
        RECT 1229.280 110.490 1229.880 110.570 ;
        RECT 1229.220 110.430 1229.880 110.490 ;
        RECT 1229.220 110.170 1229.480 110.430 ;
        RECT 1230.140 110.170 1230.400 110.490 ;
        RECT 1230.200 96.550 1230.340 110.170 ;
        RECT 1230.140 96.230 1230.400 96.550 ;
        RECT 1230.140 48.290 1230.400 48.610 ;
        RECT 1230.200 20.730 1230.340 48.290 ;
        RECT 1230.140 20.410 1230.400 20.730 ;
        RECT 1233.820 20.410 1234.080 20.730 ;
        RECT 1233.880 2.400 1234.020 20.410 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1248.510 20.640 1248.830 20.700 ;
        RECT 1251.730 20.640 1252.050 20.700 ;
        RECT 1248.510 20.500 1252.050 20.640 ;
        RECT 1248.510 20.440 1248.830 20.500 ;
        RECT 1251.730 20.440 1252.050 20.500 ;
      LAYER via ;
        RECT 1248.540 20.440 1248.800 20.700 ;
        RECT 1251.760 20.440 1252.020 20.700 ;
      LAYER met2 ;
        RECT 1248.120 220.730 1248.400 224.000 ;
        RECT 1248.120 220.590 1248.740 220.730 ;
        RECT 1248.120 220.000 1248.400 220.590 ;
        RECT 1248.600 20.730 1248.740 220.590 ;
        RECT 1248.540 20.410 1248.800 20.730 ;
        RECT 1251.760 20.410 1252.020 20.730 ;
        RECT 1251.820 2.400 1251.960 20.410 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1262.770 20.640 1263.090 20.700 ;
        RECT 1269.210 20.640 1269.530 20.700 ;
        RECT 1262.770 20.500 1269.530 20.640 ;
        RECT 1262.770 20.440 1263.090 20.500 ;
        RECT 1269.210 20.440 1269.530 20.500 ;
      LAYER via ;
        RECT 1262.800 20.440 1263.060 20.700 ;
        RECT 1269.240 20.440 1269.500 20.700 ;
      LAYER met2 ;
        RECT 1262.840 220.000 1263.120 224.000 ;
        RECT 1262.860 20.730 1263.000 220.000 ;
        RECT 1262.800 20.410 1263.060 20.730 ;
        RECT 1269.240 20.410 1269.500 20.730 ;
        RECT 1269.300 2.400 1269.440 20.410 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1277.490 207.300 1277.810 207.360 ;
        RECT 1283.470 207.300 1283.790 207.360 ;
        RECT 1277.490 207.160 1283.790 207.300 ;
        RECT 1277.490 207.100 1277.810 207.160 ;
        RECT 1283.470 207.100 1283.790 207.160 ;
        RECT 1283.470 2.960 1283.790 3.020 ;
        RECT 1287.150 2.960 1287.470 3.020 ;
        RECT 1283.470 2.820 1287.470 2.960 ;
        RECT 1283.470 2.760 1283.790 2.820 ;
        RECT 1287.150 2.760 1287.470 2.820 ;
      LAYER via ;
        RECT 1277.520 207.100 1277.780 207.360 ;
        RECT 1283.500 207.100 1283.760 207.360 ;
        RECT 1283.500 2.760 1283.760 3.020 ;
        RECT 1287.180 2.760 1287.440 3.020 ;
      LAYER met2 ;
        RECT 1277.560 220.000 1277.840 224.000 ;
        RECT 1277.580 207.390 1277.720 220.000 ;
        RECT 1277.520 207.070 1277.780 207.390 ;
        RECT 1283.500 207.070 1283.760 207.390 ;
        RECT 1283.560 3.050 1283.700 207.070 ;
        RECT 1283.500 2.730 1283.760 3.050 ;
        RECT 1287.180 2.730 1287.440 3.050 ;
        RECT 1287.240 2.400 1287.380 2.730 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1292.210 207.300 1292.530 207.360 ;
        RECT 1296.810 207.300 1297.130 207.360 ;
        RECT 1292.210 207.160 1297.130 207.300 ;
        RECT 1292.210 207.100 1292.530 207.160 ;
        RECT 1296.810 207.100 1297.130 207.160 ;
        RECT 1296.810 17.240 1297.130 17.300 ;
        RECT 1305.090 17.240 1305.410 17.300 ;
        RECT 1296.810 17.100 1305.410 17.240 ;
        RECT 1296.810 17.040 1297.130 17.100 ;
        RECT 1305.090 17.040 1305.410 17.100 ;
      LAYER via ;
        RECT 1292.240 207.100 1292.500 207.360 ;
        RECT 1296.840 207.100 1297.100 207.360 ;
        RECT 1296.840 17.040 1297.100 17.300 ;
        RECT 1305.120 17.040 1305.380 17.300 ;
      LAYER met2 ;
        RECT 1292.280 220.000 1292.560 224.000 ;
        RECT 1292.300 207.390 1292.440 220.000 ;
        RECT 1292.240 207.070 1292.500 207.390 ;
        RECT 1296.840 207.070 1297.100 207.390 ;
        RECT 1296.900 17.330 1297.040 207.070 ;
        RECT 1296.840 17.010 1297.100 17.330 ;
        RECT 1305.120 17.010 1305.380 17.330 ;
        RECT 1305.180 2.400 1305.320 17.010 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1310.610 15.540 1310.930 15.600 ;
        RECT 1323.030 15.540 1323.350 15.600 ;
        RECT 1310.610 15.400 1323.350 15.540 ;
        RECT 1310.610 15.340 1310.930 15.400 ;
        RECT 1323.030 15.340 1323.350 15.400 ;
      LAYER via ;
        RECT 1310.640 15.340 1310.900 15.600 ;
        RECT 1323.060 15.340 1323.320 15.600 ;
      LAYER met2 ;
        RECT 1307.000 220.730 1307.280 224.000 ;
        RECT 1307.000 220.590 1310.840 220.730 ;
        RECT 1307.000 220.000 1307.280 220.590 ;
        RECT 1310.700 15.630 1310.840 220.590 ;
        RECT 1310.640 15.310 1310.900 15.630 ;
        RECT 1323.060 15.310 1323.320 15.630 ;
        RECT 1323.120 2.400 1323.260 15.310 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1321.650 207.640 1321.970 207.700 ;
        RECT 1334.990 207.640 1335.310 207.700 ;
        RECT 1321.650 207.500 1335.310 207.640 ;
        RECT 1321.650 207.440 1321.970 207.500 ;
        RECT 1334.990 207.440 1335.310 207.500 ;
        RECT 1334.990 20.640 1335.310 20.700 ;
        RECT 1340.510 20.640 1340.830 20.700 ;
        RECT 1334.990 20.500 1340.830 20.640 ;
        RECT 1334.990 20.440 1335.310 20.500 ;
        RECT 1340.510 20.440 1340.830 20.500 ;
      LAYER via ;
        RECT 1321.680 207.440 1321.940 207.700 ;
        RECT 1335.020 207.440 1335.280 207.700 ;
        RECT 1335.020 20.440 1335.280 20.700 ;
        RECT 1340.540 20.440 1340.800 20.700 ;
      LAYER met2 ;
        RECT 1321.720 220.000 1322.000 224.000 ;
        RECT 1321.740 207.730 1321.880 220.000 ;
        RECT 1321.680 207.410 1321.940 207.730 ;
        RECT 1335.020 207.410 1335.280 207.730 ;
        RECT 1335.080 20.730 1335.220 207.410 ;
        RECT 1335.020 20.410 1335.280 20.730 ;
        RECT 1340.540 20.410 1340.800 20.730 ;
        RECT 1340.600 2.400 1340.740 20.410 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 703.410 208.660 703.730 208.720 ;
        RECT 792.650 208.660 792.970 208.720 ;
        RECT 703.410 208.520 792.970 208.660 ;
        RECT 703.410 208.460 703.730 208.520 ;
        RECT 792.650 208.460 792.970 208.520 ;
        RECT 698.350 17.580 698.670 17.640 ;
        RECT 703.410 17.580 703.730 17.640 ;
        RECT 698.350 17.440 703.730 17.580 ;
        RECT 698.350 17.380 698.670 17.440 ;
        RECT 703.410 17.380 703.730 17.440 ;
      LAYER via ;
        RECT 703.440 208.460 703.700 208.720 ;
        RECT 792.680 208.460 792.940 208.720 ;
        RECT 698.380 17.380 698.640 17.640 ;
        RECT 703.440 17.380 703.700 17.640 ;
      LAYER met2 ;
        RECT 792.720 220.000 793.000 224.000 ;
        RECT 792.740 208.750 792.880 220.000 ;
        RECT 703.440 208.430 703.700 208.750 ;
        RECT 792.680 208.430 792.940 208.750 ;
        RECT 703.500 17.670 703.640 208.430 ;
        RECT 698.380 17.350 698.640 17.670 ;
        RECT 703.440 17.350 703.700 17.670 ;
        RECT 698.440 2.400 698.580 17.350 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1338.210 18.600 1338.530 18.660 ;
        RECT 1358.450 18.600 1358.770 18.660 ;
        RECT 1338.210 18.460 1358.770 18.600 ;
        RECT 1338.210 18.400 1338.530 18.460 ;
        RECT 1358.450 18.400 1358.770 18.460 ;
      LAYER via ;
        RECT 1338.240 18.400 1338.500 18.660 ;
        RECT 1358.480 18.400 1358.740 18.660 ;
      LAYER met2 ;
        RECT 1336.440 220.730 1336.720 224.000 ;
        RECT 1336.440 220.590 1338.440 220.730 ;
        RECT 1336.440 220.000 1336.720 220.590 ;
        RECT 1338.300 18.690 1338.440 220.590 ;
        RECT 1338.240 18.370 1338.500 18.690 ;
        RECT 1358.480 18.370 1358.740 18.690 ;
        RECT 1358.540 2.400 1358.680 18.370 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1351.550 17.240 1351.870 17.300 ;
        RECT 1376.390 17.240 1376.710 17.300 ;
        RECT 1351.550 17.100 1376.710 17.240 ;
        RECT 1351.550 17.040 1351.870 17.100 ;
        RECT 1376.390 17.040 1376.710 17.100 ;
      LAYER via ;
        RECT 1351.580 17.040 1351.840 17.300 ;
        RECT 1376.420 17.040 1376.680 17.300 ;
      LAYER met2 ;
        RECT 1351.160 220.730 1351.440 224.000 ;
        RECT 1351.160 220.590 1351.780 220.730 ;
        RECT 1351.160 220.000 1351.440 220.590 ;
        RECT 1351.640 17.330 1351.780 220.590 ;
        RECT 1351.580 17.010 1351.840 17.330 ;
        RECT 1376.420 17.010 1376.680 17.330 ;
        RECT 1376.480 2.400 1376.620 17.010 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1365.810 19.280 1366.130 19.340 ;
        RECT 1394.330 19.280 1394.650 19.340 ;
        RECT 1365.810 19.140 1394.650 19.280 ;
        RECT 1365.810 19.080 1366.130 19.140 ;
        RECT 1394.330 19.080 1394.650 19.140 ;
      LAYER via ;
        RECT 1365.840 19.080 1366.100 19.340 ;
        RECT 1394.360 19.080 1394.620 19.340 ;
      LAYER met2 ;
        RECT 1365.880 220.000 1366.160 224.000 ;
        RECT 1365.900 19.370 1366.040 220.000 ;
        RECT 1365.840 19.050 1366.100 19.370 ;
        RECT 1394.360 19.050 1394.620 19.370 ;
        RECT 1394.420 2.400 1394.560 19.050 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1380.530 207.300 1380.850 207.360 ;
        RECT 1386.510 207.300 1386.830 207.360 ;
        RECT 1380.530 207.160 1386.830 207.300 ;
        RECT 1380.530 207.100 1380.850 207.160 ;
        RECT 1386.510 207.100 1386.830 207.160 ;
        RECT 1386.510 18.940 1386.830 19.000 ;
        RECT 1412.270 18.940 1412.590 19.000 ;
        RECT 1386.510 18.800 1412.590 18.940 ;
        RECT 1386.510 18.740 1386.830 18.800 ;
        RECT 1412.270 18.740 1412.590 18.800 ;
      LAYER via ;
        RECT 1380.560 207.100 1380.820 207.360 ;
        RECT 1386.540 207.100 1386.800 207.360 ;
        RECT 1386.540 18.740 1386.800 19.000 ;
        RECT 1412.300 18.740 1412.560 19.000 ;
      LAYER met2 ;
        RECT 1380.600 220.000 1380.880 224.000 ;
        RECT 1380.620 207.390 1380.760 220.000 ;
        RECT 1380.560 207.070 1380.820 207.390 ;
        RECT 1386.540 207.070 1386.800 207.390 ;
        RECT 1386.600 19.030 1386.740 207.070 ;
        RECT 1386.540 18.710 1386.800 19.030 ;
        RECT 1412.300 18.710 1412.560 19.030 ;
        RECT 1412.360 2.400 1412.500 18.710 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1395.250 207.300 1395.570 207.360 ;
        RECT 1400.310 207.300 1400.630 207.360 ;
        RECT 1395.250 207.160 1400.630 207.300 ;
        RECT 1395.250 207.100 1395.570 207.160 ;
        RECT 1400.310 207.100 1400.630 207.160 ;
        RECT 1400.310 17.580 1400.630 17.640 ;
        RECT 1429.750 17.580 1430.070 17.640 ;
        RECT 1400.310 17.440 1430.070 17.580 ;
        RECT 1400.310 17.380 1400.630 17.440 ;
        RECT 1429.750 17.380 1430.070 17.440 ;
      LAYER via ;
        RECT 1395.280 207.100 1395.540 207.360 ;
        RECT 1400.340 207.100 1400.600 207.360 ;
        RECT 1400.340 17.380 1400.600 17.640 ;
        RECT 1429.780 17.380 1430.040 17.640 ;
      LAYER met2 ;
        RECT 1395.320 220.000 1395.600 224.000 ;
        RECT 1395.340 207.390 1395.480 220.000 ;
        RECT 1395.280 207.070 1395.540 207.390 ;
        RECT 1400.340 207.070 1400.600 207.390 ;
        RECT 1400.400 17.670 1400.540 207.070 ;
        RECT 1400.340 17.350 1400.600 17.670 ;
        RECT 1429.780 17.350 1430.040 17.670 ;
        RECT 1429.840 2.400 1429.980 17.350 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1409.970 207.300 1410.290 207.360 ;
        RECT 1414.110 207.300 1414.430 207.360 ;
        RECT 1409.970 207.160 1414.430 207.300 ;
        RECT 1409.970 207.100 1410.290 207.160 ;
        RECT 1414.110 207.100 1414.430 207.160 ;
        RECT 1414.110 15.200 1414.430 15.260 ;
        RECT 1447.690 15.200 1448.010 15.260 ;
        RECT 1414.110 15.060 1448.010 15.200 ;
        RECT 1414.110 15.000 1414.430 15.060 ;
        RECT 1447.690 15.000 1448.010 15.060 ;
      LAYER via ;
        RECT 1410.000 207.100 1410.260 207.360 ;
        RECT 1414.140 207.100 1414.400 207.360 ;
        RECT 1414.140 15.000 1414.400 15.260 ;
        RECT 1447.720 15.000 1447.980 15.260 ;
      LAYER met2 ;
        RECT 1410.040 220.000 1410.320 224.000 ;
        RECT 1410.060 207.390 1410.200 220.000 ;
        RECT 1410.000 207.070 1410.260 207.390 ;
        RECT 1414.140 207.070 1414.400 207.390 ;
        RECT 1414.200 15.290 1414.340 207.070 ;
        RECT 1414.140 14.970 1414.400 15.290 ;
        RECT 1447.720 14.970 1447.980 15.290 ;
        RECT 1447.780 2.400 1447.920 14.970 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1427.910 19.280 1428.230 19.340 ;
        RECT 1465.630 19.280 1465.950 19.340 ;
        RECT 1427.910 19.140 1465.950 19.280 ;
        RECT 1427.910 19.080 1428.230 19.140 ;
        RECT 1465.630 19.080 1465.950 19.140 ;
      LAYER via ;
        RECT 1427.940 19.080 1428.200 19.340 ;
        RECT 1465.660 19.080 1465.920 19.340 ;
      LAYER met2 ;
        RECT 1424.760 220.730 1425.040 224.000 ;
        RECT 1424.760 220.590 1428.140 220.730 ;
        RECT 1424.760 220.000 1425.040 220.590 ;
        RECT 1428.000 19.370 1428.140 220.590 ;
        RECT 1427.940 19.050 1428.200 19.370 ;
        RECT 1465.660 19.050 1465.920 19.370 ;
        RECT 1465.720 2.400 1465.860 19.050 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1441.710 17.580 1442.030 17.640 ;
        RECT 1483.570 17.580 1483.890 17.640 ;
        RECT 1441.710 17.440 1483.890 17.580 ;
        RECT 1441.710 17.380 1442.030 17.440 ;
        RECT 1483.570 17.380 1483.890 17.440 ;
      LAYER via ;
        RECT 1441.740 17.380 1442.000 17.640 ;
        RECT 1483.600 17.380 1483.860 17.640 ;
      LAYER met2 ;
        RECT 1439.480 220.730 1439.760 224.000 ;
        RECT 1439.480 220.590 1441.940 220.730 ;
        RECT 1439.480 220.000 1439.760 220.590 ;
        RECT 1441.800 17.670 1441.940 220.590 ;
        RECT 1441.740 17.350 1442.000 17.670 ;
        RECT 1483.600 17.350 1483.860 17.670 ;
        RECT 1483.660 2.400 1483.800 17.350 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1455.050 18.260 1455.370 18.320 ;
        RECT 1501.510 18.260 1501.830 18.320 ;
        RECT 1455.050 18.120 1501.830 18.260 ;
        RECT 1455.050 18.060 1455.370 18.120 ;
        RECT 1501.510 18.060 1501.830 18.120 ;
      LAYER via ;
        RECT 1455.080 18.060 1455.340 18.320 ;
        RECT 1501.540 18.060 1501.800 18.320 ;
      LAYER met2 ;
        RECT 1454.200 220.730 1454.480 224.000 ;
        RECT 1454.200 220.590 1455.280 220.730 ;
        RECT 1454.200 220.000 1454.480 220.590 ;
        RECT 1455.140 18.350 1455.280 220.590 ;
        RECT 1455.080 18.030 1455.340 18.350 ;
        RECT 1501.540 18.030 1501.800 18.350 ;
        RECT 1501.600 2.400 1501.740 18.030 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1469.310 19.620 1469.630 19.680 ;
        RECT 1518.990 19.620 1519.310 19.680 ;
        RECT 1469.310 19.480 1519.310 19.620 ;
        RECT 1469.310 19.420 1469.630 19.480 ;
        RECT 1518.990 19.420 1519.310 19.480 ;
      LAYER via ;
        RECT 1469.340 19.420 1469.600 19.680 ;
        RECT 1519.020 19.420 1519.280 19.680 ;
      LAYER met2 ;
        RECT 1468.460 220.730 1468.740 224.000 ;
        RECT 1468.460 220.590 1469.540 220.730 ;
        RECT 1468.460 220.000 1468.740 220.590 ;
        RECT 1469.400 19.710 1469.540 220.590 ;
        RECT 1469.340 19.390 1469.600 19.710 ;
        RECT 1519.020 19.390 1519.280 19.710 ;
        RECT 1519.080 2.400 1519.220 19.390 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 717.210 210.700 717.530 210.760 ;
        RECT 807.370 210.700 807.690 210.760 ;
        RECT 717.210 210.560 807.690 210.700 ;
        RECT 717.210 210.500 717.530 210.560 ;
        RECT 807.370 210.500 807.690 210.560 ;
      LAYER via ;
        RECT 717.240 210.500 717.500 210.760 ;
        RECT 807.400 210.500 807.660 210.760 ;
      LAYER met2 ;
        RECT 807.440 220.000 807.720 224.000 ;
        RECT 807.460 210.790 807.600 220.000 ;
        RECT 717.240 210.470 717.500 210.790 ;
        RECT 807.400 210.470 807.660 210.790 ;
        RECT 717.300 16.730 717.440 210.470 ;
        RECT 716.380 16.590 717.440 16.730 ;
        RECT 716.380 2.400 716.520 16.590 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1483.110 17.240 1483.430 17.300 ;
        RECT 1536.930 17.240 1537.250 17.300 ;
        RECT 1483.110 17.100 1537.250 17.240 ;
        RECT 1483.110 17.040 1483.430 17.100 ;
        RECT 1536.930 17.040 1537.250 17.100 ;
      LAYER via ;
        RECT 1483.140 17.040 1483.400 17.300 ;
        RECT 1536.960 17.040 1537.220 17.300 ;
      LAYER met2 ;
        RECT 1483.180 220.000 1483.460 224.000 ;
        RECT 1483.200 17.330 1483.340 220.000 ;
        RECT 1483.140 17.010 1483.400 17.330 ;
        RECT 1536.960 17.010 1537.220 17.330 ;
        RECT 1537.020 2.400 1537.160 17.010 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1497.830 207.300 1498.150 207.360 ;
        RECT 1503.810 207.300 1504.130 207.360 ;
        RECT 1497.830 207.160 1504.130 207.300 ;
        RECT 1497.830 207.100 1498.150 207.160 ;
        RECT 1503.810 207.100 1504.130 207.160 ;
        RECT 1503.810 18.260 1504.130 18.320 ;
        RECT 1554.870 18.260 1555.190 18.320 ;
        RECT 1503.810 18.120 1555.190 18.260 ;
        RECT 1503.810 18.060 1504.130 18.120 ;
        RECT 1554.870 18.060 1555.190 18.120 ;
      LAYER via ;
        RECT 1497.860 207.100 1498.120 207.360 ;
        RECT 1503.840 207.100 1504.100 207.360 ;
        RECT 1503.840 18.060 1504.100 18.320 ;
        RECT 1554.900 18.060 1555.160 18.320 ;
      LAYER met2 ;
        RECT 1497.900 220.000 1498.180 224.000 ;
        RECT 1497.920 207.390 1498.060 220.000 ;
        RECT 1497.860 207.070 1498.120 207.390 ;
        RECT 1503.840 207.070 1504.100 207.390 ;
        RECT 1503.900 18.350 1504.040 207.070 ;
        RECT 1503.840 18.030 1504.100 18.350 ;
        RECT 1554.900 18.030 1555.160 18.350 ;
        RECT 1554.960 2.400 1555.100 18.030 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1512.550 207.300 1512.870 207.360 ;
        RECT 1517.610 207.300 1517.930 207.360 ;
        RECT 1512.550 207.160 1517.930 207.300 ;
        RECT 1512.550 207.100 1512.870 207.160 ;
        RECT 1517.610 207.100 1517.930 207.160 ;
        RECT 1517.610 20.640 1517.930 20.700 ;
        RECT 1571.890 20.640 1572.210 20.700 ;
        RECT 1517.610 20.500 1572.210 20.640 ;
        RECT 1517.610 20.440 1517.930 20.500 ;
        RECT 1571.890 20.440 1572.210 20.500 ;
      LAYER via ;
        RECT 1512.580 207.100 1512.840 207.360 ;
        RECT 1517.640 207.100 1517.900 207.360 ;
        RECT 1517.640 20.440 1517.900 20.700 ;
        RECT 1571.920 20.440 1572.180 20.700 ;
      LAYER met2 ;
        RECT 1512.620 220.000 1512.900 224.000 ;
        RECT 1512.640 207.390 1512.780 220.000 ;
        RECT 1512.580 207.070 1512.840 207.390 ;
        RECT 1517.640 207.070 1517.900 207.390 ;
        RECT 1517.700 20.730 1517.840 207.070 ;
        RECT 1517.640 20.410 1517.900 20.730 ;
        RECT 1571.920 20.410 1572.180 20.730 ;
        RECT 1571.980 18.090 1572.120 20.410 ;
        RECT 1571.980 17.950 1573.040 18.090 ;
        RECT 1572.900 2.400 1573.040 17.950 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1527.270 207.300 1527.590 207.360 ;
        RECT 1531.410 207.300 1531.730 207.360 ;
        RECT 1527.270 207.160 1531.730 207.300 ;
        RECT 1527.270 207.100 1527.590 207.160 ;
        RECT 1531.410 207.100 1531.730 207.160 ;
        RECT 1531.410 16.900 1531.730 16.960 ;
        RECT 1590.290 16.900 1590.610 16.960 ;
        RECT 1531.410 16.760 1590.610 16.900 ;
        RECT 1531.410 16.700 1531.730 16.760 ;
        RECT 1590.290 16.700 1590.610 16.760 ;
      LAYER via ;
        RECT 1527.300 207.100 1527.560 207.360 ;
        RECT 1531.440 207.100 1531.700 207.360 ;
        RECT 1531.440 16.700 1531.700 16.960 ;
        RECT 1590.320 16.700 1590.580 16.960 ;
      LAYER met2 ;
        RECT 1527.340 220.000 1527.620 224.000 ;
        RECT 1527.360 207.390 1527.500 220.000 ;
        RECT 1527.300 207.070 1527.560 207.390 ;
        RECT 1531.440 207.070 1531.700 207.390 ;
        RECT 1531.500 16.990 1531.640 207.070 ;
        RECT 1531.440 16.670 1531.700 16.990 ;
        RECT 1590.320 16.670 1590.580 16.990 ;
        RECT 1590.380 2.400 1590.520 16.670 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1545.210 17.920 1545.530 17.980 ;
        RECT 1608.230 17.920 1608.550 17.980 ;
        RECT 1545.210 17.780 1608.550 17.920 ;
        RECT 1545.210 17.720 1545.530 17.780 ;
        RECT 1608.230 17.720 1608.550 17.780 ;
      LAYER via ;
        RECT 1545.240 17.720 1545.500 17.980 ;
        RECT 1608.260 17.720 1608.520 17.980 ;
      LAYER met2 ;
        RECT 1542.060 220.730 1542.340 224.000 ;
        RECT 1542.060 220.590 1545.440 220.730 ;
        RECT 1542.060 220.000 1542.340 220.590 ;
        RECT 1545.300 18.010 1545.440 220.590 ;
        RECT 1545.240 17.690 1545.500 18.010 ;
        RECT 1608.260 17.690 1608.520 18.010 ;
        RECT 1608.320 2.400 1608.460 17.690 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1559.010 18.260 1559.330 18.320 ;
        RECT 1626.170 18.260 1626.490 18.320 ;
        RECT 1559.010 18.120 1626.490 18.260 ;
        RECT 1559.010 18.060 1559.330 18.120 ;
        RECT 1626.170 18.060 1626.490 18.120 ;
      LAYER via ;
        RECT 1559.040 18.060 1559.300 18.320 ;
        RECT 1626.200 18.060 1626.460 18.320 ;
      LAYER met2 ;
        RECT 1556.780 220.730 1557.060 224.000 ;
        RECT 1556.780 220.590 1559.240 220.730 ;
        RECT 1556.780 220.000 1557.060 220.590 ;
        RECT 1559.100 18.350 1559.240 220.590 ;
        RECT 1559.040 18.030 1559.300 18.350 ;
        RECT 1626.200 18.030 1626.460 18.350 ;
        RECT 1626.260 2.400 1626.400 18.030 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1572.350 18.940 1572.670 19.000 ;
        RECT 1644.110 18.940 1644.430 19.000 ;
        RECT 1572.350 18.800 1644.430 18.940 ;
        RECT 1572.350 18.740 1572.670 18.800 ;
        RECT 1644.110 18.740 1644.430 18.800 ;
      LAYER via ;
        RECT 1572.380 18.740 1572.640 19.000 ;
        RECT 1644.140 18.740 1644.400 19.000 ;
      LAYER met2 ;
        RECT 1571.500 220.730 1571.780 224.000 ;
        RECT 1571.500 220.590 1572.580 220.730 ;
        RECT 1571.500 220.000 1571.780 220.590 ;
        RECT 1572.440 19.030 1572.580 220.590 ;
        RECT 1572.380 18.710 1572.640 19.030 ;
        RECT 1644.140 18.710 1644.400 19.030 ;
        RECT 1644.200 2.400 1644.340 18.710 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1586.610 16.560 1586.930 16.620 ;
        RECT 1662.050 16.560 1662.370 16.620 ;
        RECT 1586.610 16.420 1662.370 16.560 ;
        RECT 1586.610 16.360 1586.930 16.420 ;
        RECT 1662.050 16.360 1662.370 16.420 ;
      LAYER via ;
        RECT 1586.640 16.360 1586.900 16.620 ;
        RECT 1662.080 16.360 1662.340 16.620 ;
      LAYER met2 ;
        RECT 1586.220 220.730 1586.500 224.000 ;
        RECT 1586.220 220.590 1586.840 220.730 ;
        RECT 1586.220 220.000 1586.500 220.590 ;
        RECT 1586.700 16.650 1586.840 220.590 ;
        RECT 1586.640 16.330 1586.900 16.650 ;
        RECT 1662.080 16.330 1662.340 16.650 ;
        RECT 1662.140 2.400 1662.280 16.330 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1600.870 207.300 1601.190 207.360 ;
        RECT 1607.310 207.300 1607.630 207.360 ;
        RECT 1600.870 207.160 1607.630 207.300 ;
        RECT 1600.870 207.100 1601.190 207.160 ;
        RECT 1607.310 207.100 1607.630 207.160 ;
        RECT 1607.310 14.520 1607.630 14.580 ;
        RECT 1679.530 14.520 1679.850 14.580 ;
        RECT 1607.310 14.380 1679.850 14.520 ;
        RECT 1607.310 14.320 1607.630 14.380 ;
        RECT 1679.530 14.320 1679.850 14.380 ;
      LAYER via ;
        RECT 1600.900 207.100 1601.160 207.360 ;
        RECT 1607.340 207.100 1607.600 207.360 ;
        RECT 1607.340 14.320 1607.600 14.580 ;
        RECT 1679.560 14.320 1679.820 14.580 ;
      LAYER met2 ;
        RECT 1600.940 220.000 1601.220 224.000 ;
        RECT 1600.960 207.390 1601.100 220.000 ;
        RECT 1600.900 207.070 1601.160 207.390 ;
        RECT 1607.340 207.070 1607.600 207.390 ;
        RECT 1607.400 14.610 1607.540 207.070 ;
        RECT 1607.340 14.290 1607.600 14.610 ;
        RECT 1679.560 14.290 1679.820 14.610 ;
        RECT 1679.620 2.400 1679.760 14.290 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1615.590 207.300 1615.910 207.360 ;
        RECT 1621.110 207.300 1621.430 207.360 ;
        RECT 1615.590 207.160 1621.430 207.300 ;
        RECT 1615.590 207.100 1615.910 207.160 ;
        RECT 1621.110 207.100 1621.430 207.160 ;
        RECT 1621.110 16.220 1621.430 16.280 ;
        RECT 1697.470 16.220 1697.790 16.280 ;
        RECT 1621.110 16.080 1697.790 16.220 ;
        RECT 1621.110 16.020 1621.430 16.080 ;
        RECT 1697.470 16.020 1697.790 16.080 ;
      LAYER via ;
        RECT 1615.620 207.100 1615.880 207.360 ;
        RECT 1621.140 207.100 1621.400 207.360 ;
        RECT 1621.140 16.020 1621.400 16.280 ;
        RECT 1697.500 16.020 1697.760 16.280 ;
      LAYER met2 ;
        RECT 1615.660 220.000 1615.940 224.000 ;
        RECT 1615.680 207.390 1615.820 220.000 ;
        RECT 1615.620 207.070 1615.880 207.390 ;
        RECT 1621.140 207.070 1621.400 207.390 ;
        RECT 1621.200 16.310 1621.340 207.070 ;
        RECT 1621.140 15.990 1621.400 16.310 ;
        RECT 1697.500 15.990 1697.760 16.310 ;
        RECT 1697.560 2.400 1697.700 15.990 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 737.910 211.040 738.230 211.100 ;
        RECT 822.090 211.040 822.410 211.100 ;
        RECT 737.910 210.900 822.410 211.040 ;
        RECT 737.910 210.840 738.230 210.900 ;
        RECT 822.090 210.840 822.410 210.900 ;
        RECT 734.230 17.580 734.550 17.640 ;
        RECT 737.910 17.580 738.230 17.640 ;
        RECT 734.230 17.440 738.230 17.580 ;
        RECT 734.230 17.380 734.550 17.440 ;
        RECT 737.910 17.380 738.230 17.440 ;
      LAYER via ;
        RECT 737.940 210.840 738.200 211.100 ;
        RECT 822.120 210.840 822.380 211.100 ;
        RECT 734.260 17.380 734.520 17.640 ;
        RECT 737.940 17.380 738.200 17.640 ;
      LAYER met2 ;
        RECT 822.160 220.000 822.440 224.000 ;
        RECT 822.180 211.130 822.320 220.000 ;
        RECT 737.940 210.810 738.200 211.130 ;
        RECT 822.120 210.810 822.380 211.130 ;
        RECT 738.000 17.670 738.140 210.810 ;
        RECT 734.260 17.350 734.520 17.670 ;
        RECT 737.940 17.350 738.200 17.670 ;
        RECT 734.320 2.400 734.460 17.350 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1630.310 207.300 1630.630 207.360 ;
        RECT 1634.450 207.300 1634.770 207.360 ;
        RECT 1630.310 207.160 1634.770 207.300 ;
        RECT 1630.310 207.100 1630.630 207.160 ;
        RECT 1634.450 207.100 1634.770 207.160 ;
        RECT 1634.450 18.260 1634.770 18.320 ;
        RECT 1715.410 18.260 1715.730 18.320 ;
        RECT 1634.450 18.120 1715.730 18.260 ;
        RECT 1634.450 18.060 1634.770 18.120 ;
        RECT 1715.410 18.060 1715.730 18.120 ;
      LAYER via ;
        RECT 1630.340 207.100 1630.600 207.360 ;
        RECT 1634.480 207.100 1634.740 207.360 ;
        RECT 1634.480 18.060 1634.740 18.320 ;
        RECT 1715.440 18.060 1715.700 18.320 ;
      LAYER met2 ;
        RECT 1630.380 220.000 1630.660 224.000 ;
        RECT 1630.400 207.390 1630.540 220.000 ;
        RECT 1630.340 207.070 1630.600 207.390 ;
        RECT 1634.480 207.070 1634.740 207.390 ;
        RECT 1634.540 18.350 1634.680 207.070 ;
        RECT 1634.480 18.030 1634.740 18.350 ;
        RECT 1715.440 18.030 1715.700 18.350 ;
        RECT 1715.500 2.400 1715.640 18.030 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1645.030 207.300 1645.350 207.360 ;
        RECT 1648.710 207.300 1649.030 207.360 ;
        RECT 1645.030 207.160 1649.030 207.300 ;
        RECT 1645.030 207.100 1645.350 207.160 ;
        RECT 1648.710 207.100 1649.030 207.160 ;
        RECT 1648.710 16.900 1649.030 16.960 ;
        RECT 1733.350 16.900 1733.670 16.960 ;
        RECT 1648.710 16.760 1733.670 16.900 ;
        RECT 1648.710 16.700 1649.030 16.760 ;
        RECT 1733.350 16.700 1733.670 16.760 ;
      LAYER via ;
        RECT 1645.060 207.100 1645.320 207.360 ;
        RECT 1648.740 207.100 1649.000 207.360 ;
        RECT 1648.740 16.700 1649.000 16.960 ;
        RECT 1733.380 16.700 1733.640 16.960 ;
      LAYER met2 ;
        RECT 1645.100 220.000 1645.380 224.000 ;
        RECT 1645.120 207.390 1645.260 220.000 ;
        RECT 1645.060 207.070 1645.320 207.390 ;
        RECT 1648.740 207.070 1649.000 207.390 ;
        RECT 1648.800 16.990 1648.940 207.070 ;
        RECT 1648.740 16.670 1649.000 16.990 ;
        RECT 1733.380 16.670 1733.640 16.990 ;
        RECT 1733.440 2.400 1733.580 16.670 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1662.510 15.200 1662.830 15.260 ;
        RECT 1751.290 15.200 1751.610 15.260 ;
        RECT 1662.510 15.060 1751.610 15.200 ;
        RECT 1662.510 15.000 1662.830 15.060 ;
        RECT 1751.290 15.000 1751.610 15.060 ;
      LAYER via ;
        RECT 1662.540 15.000 1662.800 15.260 ;
        RECT 1751.320 15.000 1751.580 15.260 ;
      LAYER met2 ;
        RECT 1659.820 220.730 1660.100 224.000 ;
        RECT 1659.820 220.590 1662.740 220.730 ;
        RECT 1659.820 220.000 1660.100 220.590 ;
        RECT 1662.600 15.290 1662.740 220.590 ;
        RECT 1662.540 14.970 1662.800 15.290 ;
        RECT 1751.320 14.970 1751.580 15.290 ;
        RECT 1751.380 2.400 1751.520 14.970 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1676.310 18.940 1676.630 19.000 ;
        RECT 1768.770 18.940 1769.090 19.000 ;
        RECT 1676.310 18.800 1769.090 18.940 ;
        RECT 1676.310 18.740 1676.630 18.800 ;
        RECT 1768.770 18.740 1769.090 18.800 ;
      LAYER via ;
        RECT 1676.340 18.740 1676.600 19.000 ;
        RECT 1768.800 18.740 1769.060 19.000 ;
      LAYER met2 ;
        RECT 1674.540 220.730 1674.820 224.000 ;
        RECT 1674.540 220.590 1676.540 220.730 ;
        RECT 1674.540 220.000 1674.820 220.590 ;
        RECT 1676.400 19.030 1676.540 220.590 ;
        RECT 1676.340 18.710 1676.600 19.030 ;
        RECT 1768.800 18.710 1769.060 19.030 ;
        RECT 1768.860 2.400 1769.000 18.710 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1689.650 17.240 1689.970 17.300 ;
        RECT 1786.710 17.240 1787.030 17.300 ;
        RECT 1689.650 17.100 1787.030 17.240 ;
        RECT 1689.650 17.040 1689.970 17.100 ;
        RECT 1786.710 17.040 1787.030 17.100 ;
      LAYER via ;
        RECT 1689.680 17.040 1689.940 17.300 ;
        RECT 1786.740 17.040 1787.000 17.300 ;
      LAYER met2 ;
        RECT 1689.260 220.730 1689.540 224.000 ;
        RECT 1689.260 220.590 1689.880 220.730 ;
        RECT 1689.260 220.000 1689.540 220.590 ;
        RECT 1689.740 17.330 1689.880 220.590 ;
        RECT 1689.680 17.010 1689.940 17.330 ;
        RECT 1786.740 17.010 1787.000 17.330 ;
        RECT 1786.800 2.400 1786.940 17.010 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.910 17.580 1704.230 17.640 ;
        RECT 1804.650 17.580 1804.970 17.640 ;
        RECT 1703.910 17.440 1804.970 17.580 ;
        RECT 1703.910 17.380 1704.230 17.440 ;
        RECT 1804.650 17.380 1804.970 17.440 ;
      LAYER via ;
        RECT 1703.940 17.380 1704.200 17.640 ;
        RECT 1804.680 17.380 1804.940 17.640 ;
      LAYER met2 ;
        RECT 1703.980 220.730 1704.260 224.000 ;
        RECT 1703.540 220.590 1704.260 220.730 ;
        RECT 1703.540 26.250 1703.680 220.590 ;
        RECT 1703.980 220.000 1704.260 220.590 ;
        RECT 1703.540 26.110 1704.140 26.250 ;
        RECT 1704.000 17.670 1704.140 26.110 ;
        RECT 1703.940 17.350 1704.200 17.670 ;
        RECT 1804.680 17.350 1804.940 17.670 ;
        RECT 1804.740 2.400 1804.880 17.350 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1718.170 207.300 1718.490 207.360 ;
        RECT 1724.610 207.300 1724.930 207.360 ;
        RECT 1718.170 207.160 1724.930 207.300 ;
        RECT 1718.170 207.100 1718.490 207.160 ;
        RECT 1724.610 207.100 1724.930 207.160 ;
        RECT 1724.610 20.300 1724.930 20.360 ;
        RECT 1822.590 20.300 1822.910 20.360 ;
        RECT 1724.610 20.160 1822.910 20.300 ;
        RECT 1724.610 20.100 1724.930 20.160 ;
        RECT 1822.590 20.100 1822.910 20.160 ;
      LAYER via ;
        RECT 1718.200 207.100 1718.460 207.360 ;
        RECT 1724.640 207.100 1724.900 207.360 ;
        RECT 1724.640 20.100 1724.900 20.360 ;
        RECT 1822.620 20.100 1822.880 20.360 ;
      LAYER met2 ;
        RECT 1718.240 220.000 1718.520 224.000 ;
        RECT 1718.260 207.390 1718.400 220.000 ;
        RECT 1718.200 207.070 1718.460 207.390 ;
        RECT 1724.640 207.070 1724.900 207.390 ;
        RECT 1724.700 20.390 1724.840 207.070 ;
        RECT 1724.640 20.070 1724.900 20.390 ;
        RECT 1822.620 20.070 1822.880 20.390 ;
        RECT 1822.680 2.400 1822.820 20.070 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1732.890 207.300 1733.210 207.360 ;
        RECT 1738.410 207.300 1738.730 207.360 ;
        RECT 1732.890 207.160 1738.730 207.300 ;
        RECT 1732.890 207.100 1733.210 207.160 ;
        RECT 1738.410 207.100 1738.730 207.160 ;
        RECT 1738.410 16.900 1738.730 16.960 ;
        RECT 1840.070 16.900 1840.390 16.960 ;
        RECT 1738.410 16.760 1840.390 16.900 ;
        RECT 1738.410 16.700 1738.730 16.760 ;
        RECT 1840.070 16.700 1840.390 16.760 ;
      LAYER via ;
        RECT 1732.920 207.100 1733.180 207.360 ;
        RECT 1738.440 207.100 1738.700 207.360 ;
        RECT 1738.440 16.700 1738.700 16.960 ;
        RECT 1840.100 16.700 1840.360 16.960 ;
      LAYER met2 ;
        RECT 1732.960 220.000 1733.240 224.000 ;
        RECT 1732.980 207.390 1733.120 220.000 ;
        RECT 1732.920 207.070 1733.180 207.390 ;
        RECT 1738.440 207.070 1738.700 207.390 ;
        RECT 1738.500 16.990 1738.640 207.070 ;
        RECT 1738.440 16.670 1738.700 16.990 ;
        RECT 1840.100 16.670 1840.360 16.990 ;
        RECT 1840.160 2.400 1840.300 16.670 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1747.610 207.300 1747.930 207.360 ;
        RECT 1752.210 207.300 1752.530 207.360 ;
        RECT 1747.610 207.160 1752.530 207.300 ;
        RECT 1747.610 207.100 1747.930 207.160 ;
        RECT 1752.210 207.100 1752.530 207.160 ;
        RECT 1752.210 19.960 1752.530 20.020 ;
        RECT 1858.010 19.960 1858.330 20.020 ;
        RECT 1752.210 19.820 1858.330 19.960 ;
        RECT 1752.210 19.760 1752.530 19.820 ;
        RECT 1858.010 19.760 1858.330 19.820 ;
      LAYER via ;
        RECT 1747.640 207.100 1747.900 207.360 ;
        RECT 1752.240 207.100 1752.500 207.360 ;
        RECT 1752.240 19.760 1752.500 20.020 ;
        RECT 1858.040 19.760 1858.300 20.020 ;
      LAYER met2 ;
        RECT 1747.680 220.000 1747.960 224.000 ;
        RECT 1747.700 207.390 1747.840 220.000 ;
        RECT 1747.640 207.070 1747.900 207.390 ;
        RECT 1752.240 207.070 1752.500 207.390 ;
        RECT 1752.300 20.050 1752.440 207.070 ;
        RECT 1752.240 19.730 1752.500 20.050 ;
        RECT 1858.040 19.730 1858.300 20.050 ;
        RECT 1858.100 2.400 1858.240 19.730 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1766.010 15.200 1766.330 15.260 ;
        RECT 1875.950 15.200 1876.270 15.260 ;
        RECT 1766.010 15.060 1876.270 15.200 ;
        RECT 1766.010 15.000 1766.330 15.060 ;
        RECT 1875.950 15.000 1876.270 15.060 ;
      LAYER via ;
        RECT 1766.040 15.000 1766.300 15.260 ;
        RECT 1875.980 15.000 1876.240 15.260 ;
      LAYER met2 ;
        RECT 1762.400 220.730 1762.680 224.000 ;
        RECT 1762.400 220.590 1766.240 220.730 ;
        RECT 1762.400 220.000 1762.680 220.590 ;
        RECT 1766.100 15.290 1766.240 220.590 ;
        RECT 1766.040 14.970 1766.300 15.290 ;
        RECT 1875.980 14.970 1876.240 15.290 ;
        RECT 1876.040 2.400 1876.180 14.970 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 758.150 213.420 758.470 213.480 ;
        RECT 836.810 213.420 837.130 213.480 ;
        RECT 758.150 213.280 837.130 213.420 ;
        RECT 758.150 213.220 758.470 213.280 ;
        RECT 836.810 213.220 837.130 213.280 ;
        RECT 752.170 17.920 752.490 17.980 ;
        RECT 758.150 17.920 758.470 17.980 ;
        RECT 752.170 17.780 758.470 17.920 ;
        RECT 752.170 17.720 752.490 17.780 ;
        RECT 758.150 17.720 758.470 17.780 ;
      LAYER via ;
        RECT 758.180 213.220 758.440 213.480 ;
        RECT 836.840 213.220 837.100 213.480 ;
        RECT 752.200 17.720 752.460 17.980 ;
        RECT 758.180 17.720 758.440 17.980 ;
      LAYER met2 ;
        RECT 836.880 220.000 837.160 224.000 ;
        RECT 836.900 213.510 837.040 220.000 ;
        RECT 758.180 213.190 758.440 213.510 ;
        RECT 836.840 213.190 837.100 213.510 ;
        RECT 758.240 18.010 758.380 213.190 ;
        RECT 752.200 17.690 752.460 18.010 ;
        RECT 758.180 17.690 758.440 18.010 ;
        RECT 752.260 2.400 752.400 17.690 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1779.810 19.280 1780.130 19.340 ;
        RECT 1893.890 19.280 1894.210 19.340 ;
        RECT 1779.810 19.140 1894.210 19.280 ;
        RECT 1779.810 19.080 1780.130 19.140 ;
        RECT 1893.890 19.080 1894.210 19.140 ;
      LAYER via ;
        RECT 1779.840 19.080 1780.100 19.340 ;
        RECT 1893.920 19.080 1894.180 19.340 ;
      LAYER met2 ;
        RECT 1777.120 220.730 1777.400 224.000 ;
        RECT 1777.120 220.590 1780.040 220.730 ;
        RECT 1777.120 220.000 1777.400 220.590 ;
        RECT 1779.900 19.370 1780.040 220.590 ;
        RECT 1779.840 19.050 1780.100 19.370 ;
        RECT 1893.920 19.050 1894.180 19.370 ;
        RECT 1893.980 2.400 1894.120 19.050 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1793.150 17.240 1793.470 17.300 ;
        RECT 1911.830 17.240 1912.150 17.300 ;
        RECT 1793.150 17.100 1912.150 17.240 ;
        RECT 1793.150 17.040 1793.470 17.100 ;
        RECT 1911.830 17.040 1912.150 17.100 ;
      LAYER via ;
        RECT 1793.180 17.040 1793.440 17.300 ;
        RECT 1911.860 17.040 1912.120 17.300 ;
      LAYER met2 ;
        RECT 1791.840 220.730 1792.120 224.000 ;
        RECT 1791.840 220.590 1793.380 220.730 ;
        RECT 1791.840 220.000 1792.120 220.590 ;
        RECT 1793.240 17.330 1793.380 220.590 ;
        RECT 1793.180 17.010 1793.440 17.330 ;
        RECT 1911.860 17.010 1912.120 17.330 ;
        RECT 1911.920 2.400 1912.060 17.010 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1806.950 17.920 1807.270 17.980 ;
        RECT 1929.310 17.920 1929.630 17.980 ;
        RECT 1806.950 17.780 1929.630 17.920 ;
        RECT 1806.950 17.720 1807.270 17.780 ;
        RECT 1929.310 17.720 1929.630 17.780 ;
      LAYER via ;
        RECT 1806.980 17.720 1807.240 17.980 ;
        RECT 1929.340 17.720 1929.600 17.980 ;
      LAYER met2 ;
        RECT 1806.560 220.730 1806.840 224.000 ;
        RECT 1806.560 220.590 1807.180 220.730 ;
        RECT 1806.560 220.000 1806.840 220.590 ;
        RECT 1807.040 18.010 1807.180 220.590 ;
        RECT 1806.980 17.690 1807.240 18.010 ;
        RECT 1929.340 17.690 1929.600 18.010 ;
        RECT 1929.400 2.400 1929.540 17.690 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1820.750 17.580 1821.070 17.640 ;
        RECT 1947.250 17.580 1947.570 17.640 ;
        RECT 1820.750 17.440 1947.570 17.580 ;
        RECT 1820.750 17.380 1821.070 17.440 ;
        RECT 1947.250 17.380 1947.570 17.440 ;
      LAYER via ;
        RECT 1820.780 17.380 1821.040 17.640 ;
        RECT 1947.280 17.380 1947.540 17.640 ;
      LAYER met2 ;
        RECT 1821.280 220.730 1821.560 224.000 ;
        RECT 1820.840 220.590 1821.560 220.730 ;
        RECT 1820.840 17.670 1820.980 220.590 ;
        RECT 1821.280 220.000 1821.560 220.590 ;
        RECT 1820.780 17.350 1821.040 17.670 ;
        RECT 1947.280 17.350 1947.540 17.670 ;
        RECT 1947.340 2.400 1947.480 17.350 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1835.930 207.300 1836.250 207.360 ;
        RECT 1841.910 207.300 1842.230 207.360 ;
        RECT 1835.930 207.160 1842.230 207.300 ;
        RECT 1835.930 207.100 1836.250 207.160 ;
        RECT 1841.910 207.100 1842.230 207.160 ;
        RECT 1841.910 20.640 1842.230 20.700 ;
        RECT 1965.190 20.640 1965.510 20.700 ;
        RECT 1841.910 20.500 1965.510 20.640 ;
        RECT 1841.910 20.440 1842.230 20.500 ;
        RECT 1965.190 20.440 1965.510 20.500 ;
      LAYER via ;
        RECT 1835.960 207.100 1836.220 207.360 ;
        RECT 1841.940 207.100 1842.200 207.360 ;
        RECT 1841.940 20.440 1842.200 20.700 ;
        RECT 1965.220 20.440 1965.480 20.700 ;
      LAYER met2 ;
        RECT 1836.000 220.000 1836.280 224.000 ;
        RECT 1836.020 207.390 1836.160 220.000 ;
        RECT 1835.960 207.070 1836.220 207.390 ;
        RECT 1841.940 207.070 1842.200 207.390 ;
        RECT 1842.000 20.730 1842.140 207.070 ;
        RECT 1841.940 20.410 1842.200 20.730 ;
        RECT 1965.220 20.410 1965.480 20.730 ;
        RECT 1965.280 2.400 1965.420 20.410 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1850.650 207.300 1850.970 207.360 ;
        RECT 1855.710 207.300 1856.030 207.360 ;
        RECT 1850.650 207.160 1856.030 207.300 ;
        RECT 1850.650 207.100 1850.970 207.160 ;
        RECT 1855.710 207.100 1856.030 207.160 ;
        RECT 1855.710 20.300 1856.030 20.360 ;
        RECT 1983.130 20.300 1983.450 20.360 ;
        RECT 1855.710 20.160 1983.450 20.300 ;
        RECT 1855.710 20.100 1856.030 20.160 ;
        RECT 1983.130 20.100 1983.450 20.160 ;
      LAYER via ;
        RECT 1850.680 207.100 1850.940 207.360 ;
        RECT 1855.740 207.100 1856.000 207.360 ;
        RECT 1855.740 20.100 1856.000 20.360 ;
        RECT 1983.160 20.100 1983.420 20.360 ;
      LAYER met2 ;
        RECT 1850.720 220.000 1851.000 224.000 ;
        RECT 1850.740 207.390 1850.880 220.000 ;
        RECT 1850.680 207.070 1850.940 207.390 ;
        RECT 1855.740 207.070 1856.000 207.390 ;
        RECT 1855.800 20.390 1855.940 207.070 ;
        RECT 1855.740 20.070 1856.000 20.390 ;
        RECT 1983.160 20.070 1983.420 20.390 ;
        RECT 1983.220 2.400 1983.360 20.070 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1979.525 16.745 1979.695 19.975 ;
      LAYER mcon ;
        RECT 1979.525 19.805 1979.695 19.975 ;
      LAYER met1 ;
        RECT 1865.370 207.300 1865.690 207.360 ;
        RECT 1869.510 207.300 1869.830 207.360 ;
        RECT 1865.370 207.160 1869.830 207.300 ;
        RECT 1865.370 207.100 1865.690 207.160 ;
        RECT 1869.510 207.100 1869.830 207.160 ;
        RECT 1869.510 19.960 1869.830 20.020 ;
        RECT 1979.465 19.960 1979.755 20.005 ;
        RECT 1869.510 19.820 1979.755 19.960 ;
        RECT 1869.510 19.760 1869.830 19.820 ;
        RECT 1979.465 19.775 1979.755 19.820 ;
        RECT 1979.465 16.900 1979.755 16.945 ;
        RECT 2001.070 16.900 2001.390 16.960 ;
        RECT 1979.465 16.760 2001.390 16.900 ;
        RECT 1979.465 16.715 1979.755 16.760 ;
        RECT 2001.070 16.700 2001.390 16.760 ;
      LAYER via ;
        RECT 1865.400 207.100 1865.660 207.360 ;
        RECT 1869.540 207.100 1869.800 207.360 ;
        RECT 1869.540 19.760 1869.800 20.020 ;
        RECT 2001.100 16.700 2001.360 16.960 ;
      LAYER met2 ;
        RECT 1865.440 220.000 1865.720 224.000 ;
        RECT 1865.460 207.390 1865.600 220.000 ;
        RECT 1865.400 207.070 1865.660 207.390 ;
        RECT 1869.540 207.070 1869.800 207.390 ;
        RECT 1869.600 20.050 1869.740 207.070 ;
        RECT 1869.540 19.730 1869.800 20.050 ;
        RECT 2001.100 16.670 2001.360 16.990 ;
        RECT 2001.160 2.400 2001.300 16.670 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1883.310 16.220 1883.630 16.280 ;
        RECT 2018.550 16.220 2018.870 16.280 ;
        RECT 1883.310 16.080 2018.870 16.220 ;
        RECT 1883.310 16.020 1883.630 16.080 ;
        RECT 2018.550 16.020 2018.870 16.080 ;
      LAYER via ;
        RECT 1883.340 16.020 1883.600 16.280 ;
        RECT 2018.580 16.020 2018.840 16.280 ;
      LAYER met2 ;
        RECT 1880.160 220.730 1880.440 224.000 ;
        RECT 1880.160 220.590 1883.540 220.730 ;
        RECT 1880.160 220.000 1880.440 220.590 ;
        RECT 1883.400 16.310 1883.540 220.590 ;
        RECT 1883.340 15.990 1883.600 16.310 ;
        RECT 2018.580 15.990 2018.840 16.310 ;
        RECT 2018.640 2.400 2018.780 15.990 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1897.110 19.280 1897.430 19.340 ;
        RECT 2036.490 19.280 2036.810 19.340 ;
        RECT 1897.110 19.140 2036.810 19.280 ;
        RECT 1897.110 19.080 1897.430 19.140 ;
        RECT 2036.490 19.080 2036.810 19.140 ;
      LAYER via ;
        RECT 1897.140 19.080 1897.400 19.340 ;
        RECT 2036.520 19.080 2036.780 19.340 ;
      LAYER met2 ;
        RECT 1894.880 220.730 1895.160 224.000 ;
        RECT 1894.880 220.590 1897.340 220.730 ;
        RECT 1894.880 220.000 1895.160 220.590 ;
        RECT 1897.200 19.370 1897.340 220.590 ;
        RECT 1897.140 19.050 1897.400 19.370 ;
        RECT 2036.520 19.050 2036.780 19.370 ;
        RECT 2036.580 2.400 2036.720 19.050 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1910.450 18.600 1910.770 18.660 ;
        RECT 2054.430 18.600 2054.750 18.660 ;
        RECT 1910.450 18.460 2054.750 18.600 ;
        RECT 1910.450 18.400 1910.770 18.460 ;
        RECT 2054.430 18.400 2054.750 18.460 ;
      LAYER via ;
        RECT 1910.480 18.400 1910.740 18.660 ;
        RECT 2054.460 18.400 2054.720 18.660 ;
      LAYER met2 ;
        RECT 1909.600 220.730 1909.880 224.000 ;
        RECT 1909.600 220.590 1910.680 220.730 ;
        RECT 1909.600 220.000 1909.880 220.590 ;
        RECT 1910.540 18.690 1910.680 220.590 ;
        RECT 1910.480 18.370 1910.740 18.690 ;
        RECT 2054.460 18.370 2054.720 18.690 ;
        RECT 2054.520 2.400 2054.660 18.370 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 772.410 213.760 772.730 213.820 ;
        RECT 851.530 213.760 851.850 213.820 ;
        RECT 772.410 213.620 851.850 213.760 ;
        RECT 772.410 213.560 772.730 213.620 ;
        RECT 851.530 213.560 851.850 213.620 ;
        RECT 769.650 17.580 769.970 17.640 ;
        RECT 772.410 17.580 772.730 17.640 ;
        RECT 769.650 17.440 772.730 17.580 ;
        RECT 769.650 17.380 769.970 17.440 ;
        RECT 772.410 17.380 772.730 17.440 ;
      LAYER via ;
        RECT 772.440 213.560 772.700 213.820 ;
        RECT 851.560 213.560 851.820 213.820 ;
        RECT 769.680 17.380 769.940 17.640 ;
        RECT 772.440 17.380 772.700 17.640 ;
      LAYER met2 ;
        RECT 851.600 220.000 851.880 224.000 ;
        RECT 851.620 213.850 851.760 220.000 ;
        RECT 772.440 213.530 772.700 213.850 ;
        RECT 851.560 213.530 851.820 213.850 ;
        RECT 772.500 17.670 772.640 213.530 ;
        RECT 769.680 17.350 769.940 17.670 ;
        RECT 772.440 17.350 772.700 17.670 ;
        RECT 769.740 2.400 769.880 17.350 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1924.250 17.240 1924.570 17.300 ;
        RECT 2072.370 17.240 2072.690 17.300 ;
        RECT 1924.250 17.100 2072.690 17.240 ;
        RECT 1924.250 17.040 1924.570 17.100 ;
        RECT 2072.370 17.040 2072.690 17.100 ;
      LAYER via ;
        RECT 1924.280 17.040 1924.540 17.300 ;
        RECT 2072.400 17.040 2072.660 17.300 ;
      LAYER met2 ;
        RECT 1924.320 220.000 1924.600 224.000 ;
        RECT 1924.340 17.330 1924.480 220.000 ;
        RECT 1924.280 17.010 1924.540 17.330 ;
        RECT 2072.400 17.010 2072.660 17.330 ;
        RECT 2072.460 2.400 2072.600 17.010 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1938.970 207.300 1939.290 207.360 ;
        RECT 1945.410 207.300 1945.730 207.360 ;
        RECT 1938.970 207.160 1945.730 207.300 ;
        RECT 1938.970 207.100 1939.290 207.160 ;
        RECT 1945.410 207.100 1945.730 207.160 ;
        RECT 1945.410 15.200 1945.730 15.260 ;
        RECT 2089.850 15.200 2090.170 15.260 ;
        RECT 1945.410 15.060 2090.170 15.200 ;
        RECT 1945.410 15.000 1945.730 15.060 ;
        RECT 2089.850 15.000 2090.170 15.060 ;
      LAYER via ;
        RECT 1939.000 207.100 1939.260 207.360 ;
        RECT 1945.440 207.100 1945.700 207.360 ;
        RECT 1945.440 15.000 1945.700 15.260 ;
        RECT 2089.880 15.000 2090.140 15.260 ;
      LAYER met2 ;
        RECT 1939.040 220.000 1939.320 224.000 ;
        RECT 1939.060 207.390 1939.200 220.000 ;
        RECT 1939.000 207.070 1939.260 207.390 ;
        RECT 1945.440 207.070 1945.700 207.390 ;
        RECT 1945.500 15.290 1945.640 207.070 ;
        RECT 1945.440 14.970 1945.700 15.290 ;
        RECT 2089.880 14.970 2090.140 15.290 ;
        RECT 2089.940 2.400 2090.080 14.970 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1953.690 207.300 1954.010 207.360 ;
        RECT 1959.210 207.300 1959.530 207.360 ;
        RECT 1953.690 207.160 1959.530 207.300 ;
        RECT 1953.690 207.100 1954.010 207.160 ;
        RECT 1959.210 207.100 1959.530 207.160 ;
        RECT 2107.790 15.880 2108.110 15.940 ;
        RECT 1959.760 15.740 2108.110 15.880 ;
        RECT 1958.750 15.540 1959.070 15.600 ;
        RECT 1959.760 15.540 1959.900 15.740 ;
        RECT 2107.790 15.680 2108.110 15.740 ;
        RECT 1958.750 15.400 1959.900 15.540 ;
        RECT 1958.750 15.340 1959.070 15.400 ;
      LAYER via ;
        RECT 1953.720 207.100 1953.980 207.360 ;
        RECT 1959.240 207.100 1959.500 207.360 ;
        RECT 1958.780 15.340 1959.040 15.600 ;
        RECT 2107.820 15.680 2108.080 15.940 ;
      LAYER met2 ;
        RECT 1953.760 220.000 1954.040 224.000 ;
        RECT 1953.780 207.390 1953.920 220.000 ;
        RECT 1953.720 207.070 1953.980 207.390 ;
        RECT 1959.240 207.070 1959.500 207.390 ;
        RECT 1959.300 23.530 1959.440 207.070 ;
        RECT 1958.840 23.390 1959.440 23.530 ;
        RECT 1958.840 15.630 1958.980 23.390 ;
        RECT 2107.820 15.650 2108.080 15.970 ;
        RECT 1958.780 15.310 1959.040 15.630 ;
        RECT 2107.880 2.400 2108.020 15.650 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1967.950 207.300 1968.270 207.360 ;
        RECT 1973.010 207.300 1973.330 207.360 ;
        RECT 1967.950 207.160 1973.330 207.300 ;
        RECT 1967.950 207.100 1968.270 207.160 ;
        RECT 1973.010 207.100 1973.330 207.160 ;
        RECT 1973.010 20.640 1973.330 20.700 ;
        RECT 2125.730 20.640 2126.050 20.700 ;
        RECT 1973.010 20.500 2126.050 20.640 ;
        RECT 1973.010 20.440 1973.330 20.500 ;
        RECT 2125.730 20.440 2126.050 20.500 ;
      LAYER via ;
        RECT 1967.980 207.100 1968.240 207.360 ;
        RECT 1973.040 207.100 1973.300 207.360 ;
        RECT 1973.040 20.440 1973.300 20.700 ;
        RECT 2125.760 20.440 2126.020 20.700 ;
      LAYER met2 ;
        RECT 1968.020 220.000 1968.300 224.000 ;
        RECT 1968.040 207.390 1968.180 220.000 ;
        RECT 1967.980 207.070 1968.240 207.390 ;
        RECT 1973.040 207.070 1973.300 207.390 ;
        RECT 1973.100 20.730 1973.240 207.070 ;
        RECT 1973.040 20.410 1973.300 20.730 ;
        RECT 2125.760 20.410 2126.020 20.730 ;
        RECT 2125.820 2.400 2125.960 20.410 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1982.670 207.640 1982.990 207.700 ;
        RECT 1982.670 207.500 1997.160 207.640 ;
        RECT 1982.670 207.440 1982.990 207.500 ;
        RECT 1997.020 206.620 1997.160 207.500 ;
        RECT 1997.390 206.620 1997.710 206.680 ;
        RECT 1997.020 206.480 1997.710 206.620 ;
        RECT 1997.390 206.420 1997.710 206.480 ;
        RECT 1997.850 15.540 1998.170 15.600 ;
        RECT 2143.670 15.540 2143.990 15.600 ;
        RECT 1997.850 15.400 2143.990 15.540 ;
        RECT 1997.850 15.340 1998.170 15.400 ;
        RECT 2143.670 15.340 2143.990 15.400 ;
      LAYER via ;
        RECT 1982.700 207.440 1982.960 207.700 ;
        RECT 1997.420 206.420 1997.680 206.680 ;
        RECT 1997.880 15.340 1998.140 15.600 ;
        RECT 2143.700 15.340 2143.960 15.600 ;
      LAYER met2 ;
        RECT 1982.740 220.000 1983.020 224.000 ;
        RECT 1982.760 207.730 1982.900 220.000 ;
        RECT 1982.700 207.410 1982.960 207.730 ;
        RECT 1997.420 206.390 1997.680 206.710 ;
        RECT 1997.480 158.850 1997.620 206.390 ;
        RECT 1997.480 158.710 1998.080 158.850 ;
        RECT 1997.940 134.370 1998.080 158.710 ;
        RECT 1997.480 134.230 1998.080 134.370 ;
        RECT 1997.480 62.290 1997.620 134.230 ;
        RECT 1997.480 62.150 1998.080 62.290 ;
        RECT 1997.940 15.630 1998.080 62.150 ;
        RECT 1997.880 15.310 1998.140 15.630 ;
        RECT 2143.700 15.310 2143.960 15.630 ;
        RECT 2143.760 2.400 2143.900 15.310 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1997.390 213.420 1997.710 213.480 ;
        RECT 2011.190 213.420 2011.510 213.480 ;
        RECT 1997.390 213.280 2011.510 213.420 ;
        RECT 1997.390 213.220 1997.710 213.280 ;
        RECT 2011.190 213.220 2011.510 213.280 ;
        RECT 2011.190 19.620 2011.510 19.680 ;
        RECT 2013.950 19.620 2014.270 19.680 ;
        RECT 2011.190 19.480 2014.270 19.620 ;
        RECT 2011.190 19.420 2011.510 19.480 ;
        RECT 2013.950 19.420 2014.270 19.480 ;
        RECT 2013.950 16.560 2014.270 16.620 ;
        RECT 2161.610 16.560 2161.930 16.620 ;
        RECT 2013.950 16.420 2161.930 16.560 ;
        RECT 2013.950 16.360 2014.270 16.420 ;
        RECT 2161.610 16.360 2161.930 16.420 ;
      LAYER via ;
        RECT 1997.420 213.220 1997.680 213.480 ;
        RECT 2011.220 213.220 2011.480 213.480 ;
        RECT 2011.220 19.420 2011.480 19.680 ;
        RECT 2013.980 19.420 2014.240 19.680 ;
        RECT 2013.980 16.360 2014.240 16.620 ;
        RECT 2161.640 16.360 2161.900 16.620 ;
      LAYER met2 ;
        RECT 1997.460 220.000 1997.740 224.000 ;
        RECT 1997.480 213.510 1997.620 220.000 ;
        RECT 1997.420 213.190 1997.680 213.510 ;
        RECT 2011.220 213.190 2011.480 213.510 ;
        RECT 2011.280 19.710 2011.420 213.190 ;
        RECT 2011.220 19.390 2011.480 19.710 ;
        RECT 2013.980 19.390 2014.240 19.710 ;
        RECT 2014.040 16.650 2014.180 19.390 ;
        RECT 2013.980 16.330 2014.240 16.650 ;
        RECT 2161.640 16.330 2161.900 16.650 ;
        RECT 2161.700 2.400 2161.840 16.330 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2169.890 213.080 2170.210 213.140 ;
        RECT 2042.100 212.940 2170.210 213.080 ;
        RECT 2012.110 212.400 2012.430 212.460 ;
        RECT 2042.100 212.400 2042.240 212.940 ;
        RECT 2169.890 212.880 2170.210 212.940 ;
        RECT 2012.110 212.260 2042.240 212.400 ;
        RECT 2012.110 212.200 2012.430 212.260 ;
        RECT 2169.890 20.640 2170.210 20.700 ;
        RECT 2179.090 20.640 2179.410 20.700 ;
        RECT 2169.890 20.500 2179.410 20.640 ;
        RECT 2169.890 20.440 2170.210 20.500 ;
        RECT 2179.090 20.440 2179.410 20.500 ;
      LAYER via ;
        RECT 2012.140 212.200 2012.400 212.460 ;
        RECT 2169.920 212.880 2170.180 213.140 ;
        RECT 2169.920 20.440 2170.180 20.700 ;
        RECT 2179.120 20.440 2179.380 20.700 ;
      LAYER met2 ;
        RECT 2012.180 220.000 2012.460 224.000 ;
        RECT 2012.200 212.490 2012.340 220.000 ;
        RECT 2169.920 212.850 2170.180 213.170 ;
        RECT 2012.140 212.170 2012.400 212.490 ;
        RECT 2169.980 20.730 2170.120 212.850 ;
        RECT 2169.920 20.410 2170.180 20.730 ;
        RECT 2179.120 20.410 2179.380 20.730 ;
        RECT 2179.180 2.400 2179.320 20.410 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2163.525 14.535 2163.695 15.895 ;
        RECT 2172.265 15.725 2172.895 15.895 ;
        RECT 2172.725 14.705 2172.895 15.725 ;
        RECT 2159.385 14.365 2163.695 14.535 ;
        RECT 2159.385 14.025 2159.555 14.365 ;
        RECT 2173.645 11.305 2173.815 14.875 ;
      LAYER mcon ;
        RECT 2163.525 15.725 2163.695 15.895 ;
        RECT 2173.645 14.705 2173.815 14.875 ;
      LAYER met1 ;
        RECT 2087.090 213.420 2087.410 213.480 ;
        RECT 2034.740 213.280 2087.410 213.420 ;
        RECT 2026.830 213.080 2027.150 213.140 ;
        RECT 2034.740 213.080 2034.880 213.280 ;
        RECT 2087.090 213.220 2087.410 213.280 ;
        RECT 2026.830 212.940 2034.880 213.080 ;
        RECT 2026.830 212.880 2027.150 212.940 ;
        RECT 2163.465 15.880 2163.755 15.925 ;
        RECT 2172.205 15.880 2172.495 15.925 ;
        RECT 2163.465 15.740 2172.495 15.880 ;
        RECT 2163.465 15.695 2163.755 15.740 ;
        RECT 2172.205 15.695 2172.495 15.740 ;
        RECT 2172.665 14.860 2172.955 14.905 ;
        RECT 2173.585 14.860 2173.875 14.905 ;
        RECT 2172.665 14.720 2173.875 14.860 ;
        RECT 2172.665 14.675 2172.955 14.720 ;
        RECT 2173.585 14.675 2173.875 14.720 ;
        RECT 2087.090 14.180 2087.410 14.240 ;
        RECT 2159.325 14.180 2159.615 14.225 ;
        RECT 2087.090 14.040 2159.615 14.180 ;
        RECT 2087.090 13.980 2087.410 14.040 ;
        RECT 2159.325 13.995 2159.615 14.040 ;
        RECT 2173.585 11.460 2173.875 11.505 ;
        RECT 2197.030 11.460 2197.350 11.520 ;
        RECT 2173.585 11.320 2197.350 11.460 ;
        RECT 2173.585 11.275 2173.875 11.320 ;
        RECT 2197.030 11.260 2197.350 11.320 ;
      LAYER via ;
        RECT 2026.860 212.880 2027.120 213.140 ;
        RECT 2087.120 213.220 2087.380 213.480 ;
        RECT 2087.120 13.980 2087.380 14.240 ;
        RECT 2197.060 11.260 2197.320 11.520 ;
      LAYER met2 ;
        RECT 2026.900 220.000 2027.180 224.000 ;
        RECT 2026.920 213.170 2027.060 220.000 ;
        RECT 2087.120 213.190 2087.380 213.510 ;
        RECT 2026.860 212.850 2027.120 213.170 ;
        RECT 2087.180 14.270 2087.320 213.190 ;
        RECT 2087.120 13.950 2087.380 14.270 ;
        RECT 2197.060 11.230 2197.320 11.550 ;
        RECT 2197.120 2.400 2197.260 11.230 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2041.550 210.360 2041.870 210.420 ;
        RECT 2214.970 210.360 2215.290 210.420 ;
        RECT 2041.550 210.220 2215.290 210.360 ;
        RECT 2041.550 210.160 2041.870 210.220 ;
        RECT 2214.970 210.160 2215.290 210.220 ;
      LAYER via ;
        RECT 2041.580 210.160 2041.840 210.420 ;
        RECT 2215.000 210.160 2215.260 210.420 ;
      LAYER met2 ;
        RECT 2041.620 220.000 2041.900 224.000 ;
        RECT 2041.640 210.450 2041.780 220.000 ;
        RECT 2041.580 210.130 2041.840 210.450 ;
        RECT 2215.000 210.130 2215.260 210.450 ;
        RECT 2215.060 2.400 2215.200 210.130 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2056.270 212.740 2056.590 212.800 ;
        RECT 2228.770 212.740 2229.090 212.800 ;
        RECT 2056.270 212.600 2229.090 212.740 ;
        RECT 2056.270 212.540 2056.590 212.600 ;
        RECT 2228.770 212.540 2229.090 212.600 ;
        RECT 2228.770 2.960 2229.090 3.020 ;
        RECT 2232.910 2.960 2233.230 3.020 ;
        RECT 2228.770 2.820 2233.230 2.960 ;
        RECT 2228.770 2.760 2229.090 2.820 ;
        RECT 2232.910 2.760 2233.230 2.820 ;
      LAYER via ;
        RECT 2056.300 212.540 2056.560 212.800 ;
        RECT 2228.800 212.540 2229.060 212.800 ;
        RECT 2228.800 2.760 2229.060 3.020 ;
        RECT 2232.940 2.760 2233.200 3.020 ;
      LAYER met2 ;
        RECT 2056.340 220.000 2056.620 224.000 ;
        RECT 2056.360 212.830 2056.500 220.000 ;
        RECT 2056.300 212.510 2056.560 212.830 ;
        RECT 2228.800 212.510 2229.060 212.830 ;
        RECT 2228.860 3.050 2229.000 212.510 ;
        RECT 2228.800 2.730 2229.060 3.050 ;
        RECT 2232.940 2.730 2233.200 3.050 ;
        RECT 2233.000 2.400 2233.140 2.730 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.110 212.400 793.430 212.460 ;
        RECT 866.250 212.400 866.570 212.460 ;
        RECT 793.110 212.260 866.570 212.400 ;
        RECT 793.110 212.200 793.430 212.260 ;
        RECT 866.250 212.200 866.570 212.260 ;
        RECT 787.590 16.560 787.910 16.620 ;
        RECT 793.110 16.560 793.430 16.620 ;
        RECT 787.590 16.420 793.430 16.560 ;
        RECT 787.590 16.360 787.910 16.420 ;
        RECT 793.110 16.360 793.430 16.420 ;
      LAYER via ;
        RECT 793.140 212.200 793.400 212.460 ;
        RECT 866.280 212.200 866.540 212.460 ;
        RECT 787.620 16.360 787.880 16.620 ;
        RECT 793.140 16.360 793.400 16.620 ;
      LAYER met2 ;
        RECT 866.320 220.000 866.600 224.000 ;
        RECT 866.340 212.490 866.480 220.000 ;
        RECT 793.140 212.170 793.400 212.490 ;
        RECT 866.280 212.170 866.540 212.490 ;
        RECT 793.200 16.650 793.340 212.170 ;
        RECT 787.620 16.330 787.880 16.650 ;
        RECT 793.140 16.330 793.400 16.650 ;
        RECT 787.680 2.400 787.820 16.330 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2158.925 13.345 2159.095 14.875 ;
      LAYER mcon ;
        RECT 2158.925 14.705 2159.095 14.875 ;
      LAYER met1 ;
        RECT 2070.990 213.760 2071.310 213.820 ;
        RECT 2114.690 213.760 2115.010 213.820 ;
        RECT 2070.990 213.620 2115.010 213.760 ;
        RECT 2070.990 213.560 2071.310 213.620 ;
        RECT 2114.690 213.560 2115.010 213.620 ;
        RECT 2114.690 14.860 2115.010 14.920 ;
        RECT 2158.865 14.860 2159.155 14.905 ;
        RECT 2114.690 14.720 2159.155 14.860 ;
        RECT 2114.690 14.660 2115.010 14.720 ;
        RECT 2158.865 14.675 2159.155 14.720 ;
        RECT 2250.850 14.180 2251.170 14.240 ;
        RECT 2159.860 14.040 2251.170 14.180 ;
        RECT 2158.865 13.500 2159.155 13.545 ;
        RECT 2159.860 13.500 2160.000 14.040 ;
        RECT 2250.850 13.980 2251.170 14.040 ;
        RECT 2158.865 13.360 2160.000 13.500 ;
        RECT 2158.865 13.315 2159.155 13.360 ;
      LAYER via ;
        RECT 2071.020 213.560 2071.280 213.820 ;
        RECT 2114.720 213.560 2114.980 213.820 ;
        RECT 2114.720 14.660 2114.980 14.920 ;
        RECT 2250.880 13.980 2251.140 14.240 ;
      LAYER met2 ;
        RECT 2071.060 220.000 2071.340 224.000 ;
        RECT 2071.080 213.850 2071.220 220.000 ;
        RECT 2071.020 213.530 2071.280 213.850 ;
        RECT 2114.720 213.530 2114.980 213.850 ;
        RECT 2114.780 14.950 2114.920 213.530 ;
        RECT 2114.720 14.630 2114.980 14.950 ;
        RECT 2250.880 13.950 2251.140 14.270 ;
        RECT 2250.940 2.400 2251.080 13.950 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2085.710 212.400 2086.030 212.460 ;
        RECT 2259.590 212.400 2259.910 212.460 ;
        RECT 2085.710 212.260 2259.910 212.400 ;
        RECT 2085.710 212.200 2086.030 212.260 ;
        RECT 2259.590 212.200 2259.910 212.260 ;
        RECT 2259.590 19.620 2259.910 19.680 ;
        RECT 2268.330 19.620 2268.650 19.680 ;
        RECT 2259.590 19.480 2268.650 19.620 ;
        RECT 2259.590 19.420 2259.910 19.480 ;
        RECT 2268.330 19.420 2268.650 19.480 ;
      LAYER via ;
        RECT 2085.740 212.200 2086.000 212.460 ;
        RECT 2259.620 212.200 2259.880 212.460 ;
        RECT 2259.620 19.420 2259.880 19.680 ;
        RECT 2268.360 19.420 2268.620 19.680 ;
      LAYER met2 ;
        RECT 2085.780 220.000 2086.060 224.000 ;
        RECT 2085.800 212.490 2085.940 220.000 ;
        RECT 2085.740 212.170 2086.000 212.490 ;
        RECT 2259.620 212.170 2259.880 212.490 ;
        RECT 2259.680 19.710 2259.820 212.170 ;
        RECT 2259.620 19.390 2259.880 19.710 ;
        RECT 2268.360 19.390 2268.620 19.710 ;
        RECT 2268.420 2.400 2268.560 19.390 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2268.865 18.445 2269.035 19.635 ;
      LAYER mcon ;
        RECT 2268.865 19.465 2269.035 19.635 ;
      LAYER met1 ;
        RECT 2100.430 207.300 2100.750 207.360 ;
        RECT 2104.110 207.300 2104.430 207.360 ;
        RECT 2100.430 207.160 2104.430 207.300 ;
        RECT 2100.430 207.100 2100.750 207.160 ;
        RECT 2104.110 207.100 2104.430 207.160 ;
        RECT 2268.805 19.620 2269.095 19.665 ;
        RECT 2286.270 19.620 2286.590 19.680 ;
        RECT 2268.805 19.480 2286.590 19.620 ;
        RECT 2268.805 19.435 2269.095 19.480 ;
        RECT 2286.270 19.420 2286.590 19.480 ;
        RECT 2268.805 18.600 2269.095 18.645 ;
        RECT 2259.220 18.460 2269.095 18.600 ;
        RECT 2104.110 18.260 2104.430 18.320 ;
        RECT 2259.220 18.260 2259.360 18.460 ;
        RECT 2268.805 18.415 2269.095 18.460 ;
        RECT 2104.110 18.120 2259.360 18.260 ;
        RECT 2104.110 18.060 2104.430 18.120 ;
      LAYER via ;
        RECT 2100.460 207.100 2100.720 207.360 ;
        RECT 2104.140 207.100 2104.400 207.360 ;
        RECT 2286.300 19.420 2286.560 19.680 ;
        RECT 2104.140 18.060 2104.400 18.320 ;
      LAYER met2 ;
        RECT 2100.500 220.000 2100.780 224.000 ;
        RECT 2100.520 207.390 2100.660 220.000 ;
        RECT 2100.460 207.070 2100.720 207.390 ;
        RECT 2104.140 207.070 2104.400 207.390 ;
        RECT 2104.200 18.350 2104.340 207.070 ;
        RECT 2286.300 19.390 2286.560 19.710 ;
        RECT 2104.140 18.030 2104.400 18.350 ;
        RECT 2286.360 2.400 2286.500 19.390 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2115.150 211.380 2115.470 211.440 ;
        RECT 2298.230 211.380 2298.550 211.440 ;
        RECT 2115.150 211.240 2298.550 211.380 ;
        RECT 2115.150 211.180 2115.470 211.240 ;
        RECT 2298.230 211.180 2298.550 211.240 ;
        RECT 2298.230 17.240 2298.550 17.300 ;
        RECT 2304.210 17.240 2304.530 17.300 ;
        RECT 2298.230 17.100 2304.530 17.240 ;
        RECT 2298.230 17.040 2298.550 17.100 ;
        RECT 2304.210 17.040 2304.530 17.100 ;
      LAYER via ;
        RECT 2115.180 211.180 2115.440 211.440 ;
        RECT 2298.260 211.180 2298.520 211.440 ;
        RECT 2298.260 17.040 2298.520 17.300 ;
        RECT 2304.240 17.040 2304.500 17.300 ;
      LAYER met2 ;
        RECT 2115.220 220.000 2115.500 224.000 ;
        RECT 2115.240 211.470 2115.380 220.000 ;
        RECT 2115.180 211.150 2115.440 211.470 ;
        RECT 2298.260 211.150 2298.520 211.470 ;
        RECT 2298.320 17.330 2298.460 211.150 ;
        RECT 2298.260 17.010 2298.520 17.330 ;
        RECT 2304.240 17.010 2304.500 17.330 ;
        RECT 2304.300 2.400 2304.440 17.010 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2129.870 211.040 2130.190 211.100 ;
        RECT 2314.790 211.040 2315.110 211.100 ;
        RECT 2129.870 210.900 2315.110 211.040 ;
        RECT 2129.870 210.840 2130.190 210.900 ;
        RECT 2314.790 210.840 2315.110 210.900 ;
        RECT 2314.790 17.580 2315.110 17.640 ;
        RECT 2322.150 17.580 2322.470 17.640 ;
        RECT 2314.790 17.440 2322.470 17.580 ;
        RECT 2314.790 17.380 2315.110 17.440 ;
        RECT 2322.150 17.380 2322.470 17.440 ;
      LAYER via ;
        RECT 2129.900 210.840 2130.160 211.100 ;
        RECT 2314.820 210.840 2315.080 211.100 ;
        RECT 2314.820 17.380 2315.080 17.640 ;
        RECT 2322.180 17.380 2322.440 17.640 ;
      LAYER met2 ;
        RECT 2129.940 220.000 2130.220 224.000 ;
        RECT 2129.960 211.130 2130.100 220.000 ;
        RECT 2129.900 210.810 2130.160 211.130 ;
        RECT 2314.820 210.810 2315.080 211.130 ;
        RECT 2314.880 17.670 2315.020 210.810 ;
        RECT 2314.820 17.350 2315.080 17.670 ;
        RECT 2322.180 17.350 2322.440 17.670 ;
        RECT 2322.240 2.400 2322.380 17.350 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2144.590 211.720 2144.910 211.780 ;
        RECT 2321.690 211.720 2322.010 211.780 ;
        RECT 2144.590 211.580 2322.010 211.720 ;
        RECT 2144.590 211.520 2144.910 211.580 ;
        RECT 2321.690 211.520 2322.010 211.580 ;
        RECT 2321.690 17.240 2322.010 17.300 ;
        RECT 2339.630 17.240 2339.950 17.300 ;
        RECT 2321.690 17.100 2339.950 17.240 ;
        RECT 2321.690 17.040 2322.010 17.100 ;
        RECT 2339.630 17.040 2339.950 17.100 ;
      LAYER via ;
        RECT 2144.620 211.520 2144.880 211.780 ;
        RECT 2321.720 211.520 2321.980 211.780 ;
        RECT 2321.720 17.040 2321.980 17.300 ;
        RECT 2339.660 17.040 2339.920 17.300 ;
      LAYER met2 ;
        RECT 2144.660 220.000 2144.940 224.000 ;
        RECT 2144.680 211.810 2144.820 220.000 ;
        RECT 2144.620 211.490 2144.880 211.810 ;
        RECT 2321.720 211.490 2321.980 211.810 ;
        RECT 2321.780 17.330 2321.920 211.490 ;
        RECT 2321.720 17.010 2321.980 17.330 ;
        RECT 2339.660 17.010 2339.920 17.330 ;
        RECT 2339.720 2.400 2339.860 17.010 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2173.645 15.385 2173.815 16.915 ;
      LAYER mcon ;
        RECT 2173.645 16.745 2173.815 16.915 ;
      LAYER met1 ;
        RECT 2173.585 16.900 2173.875 16.945 ;
        RECT 2357.570 16.900 2357.890 16.960 ;
        RECT 2173.585 16.760 2357.890 16.900 ;
        RECT 2173.585 16.715 2173.875 16.760 ;
        RECT 2357.570 16.700 2357.890 16.760 ;
        RECT 2158.850 15.540 2159.170 15.600 ;
        RECT 2173.585 15.540 2173.875 15.585 ;
        RECT 2158.850 15.400 2173.875 15.540 ;
        RECT 2158.850 15.340 2159.170 15.400 ;
        RECT 2173.585 15.355 2173.875 15.400 ;
      LAYER via ;
        RECT 2357.600 16.700 2357.860 16.960 ;
        RECT 2158.880 15.340 2159.140 15.600 ;
      LAYER met2 ;
        RECT 2159.380 220.730 2159.660 224.000 ;
        RECT 2158.940 220.590 2159.660 220.730 ;
        RECT 2158.940 15.630 2159.080 220.590 ;
        RECT 2159.380 220.000 2159.660 220.590 ;
        RECT 2357.600 16.670 2357.860 16.990 ;
        RECT 2158.880 15.310 2159.140 15.630 ;
        RECT 2357.660 2.400 2357.800 16.670 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2174.030 208.660 2174.350 208.720 ;
        RECT 2335.490 208.660 2335.810 208.720 ;
        RECT 2174.030 208.520 2335.810 208.660 ;
        RECT 2174.030 208.460 2174.350 208.520 ;
        RECT 2335.490 208.460 2335.810 208.520 ;
        RECT 2335.490 15.540 2335.810 15.600 ;
        RECT 2375.510 15.540 2375.830 15.600 ;
        RECT 2335.490 15.400 2375.830 15.540 ;
        RECT 2335.490 15.340 2335.810 15.400 ;
        RECT 2375.510 15.340 2375.830 15.400 ;
      LAYER via ;
        RECT 2174.060 208.460 2174.320 208.720 ;
        RECT 2335.520 208.460 2335.780 208.720 ;
        RECT 2335.520 15.340 2335.780 15.600 ;
        RECT 2375.540 15.340 2375.800 15.600 ;
      LAYER met2 ;
        RECT 2174.100 220.000 2174.380 224.000 ;
        RECT 2174.120 208.750 2174.260 220.000 ;
        RECT 2174.060 208.430 2174.320 208.750 ;
        RECT 2335.520 208.430 2335.780 208.750 ;
        RECT 2335.580 15.630 2335.720 208.430 ;
        RECT 2335.520 15.310 2335.780 15.630 ;
        RECT 2375.540 15.310 2375.800 15.630 ;
        RECT 2375.600 2.400 2375.740 15.310 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2210.905 16.235 2211.075 16.575 ;
        RECT 2210.905 16.065 2212.455 16.235 ;
      LAYER mcon ;
        RECT 2210.905 16.405 2211.075 16.575 ;
        RECT 2212.285 16.065 2212.455 16.235 ;
      LAYER met1 ;
        RECT 2188.750 207.300 2189.070 207.360 ;
        RECT 2193.810 207.300 2194.130 207.360 ;
        RECT 2188.750 207.160 2194.130 207.300 ;
        RECT 2188.750 207.100 2189.070 207.160 ;
        RECT 2193.810 207.100 2194.130 207.160 ;
        RECT 2193.810 16.560 2194.130 16.620 ;
        RECT 2210.845 16.560 2211.135 16.605 ;
        RECT 2193.810 16.420 2211.135 16.560 ;
        RECT 2193.810 16.360 2194.130 16.420 ;
        RECT 2210.845 16.375 2211.135 16.420 ;
        RECT 2212.225 16.220 2212.515 16.265 ;
        RECT 2393.450 16.220 2393.770 16.280 ;
        RECT 2212.225 16.080 2393.770 16.220 ;
        RECT 2212.225 16.035 2212.515 16.080 ;
        RECT 2393.450 16.020 2393.770 16.080 ;
      LAYER via ;
        RECT 2188.780 207.100 2189.040 207.360 ;
        RECT 2193.840 207.100 2194.100 207.360 ;
        RECT 2193.840 16.360 2194.100 16.620 ;
        RECT 2393.480 16.020 2393.740 16.280 ;
      LAYER met2 ;
        RECT 2188.820 220.000 2189.100 224.000 ;
        RECT 2188.840 207.390 2188.980 220.000 ;
        RECT 2188.780 207.070 2189.040 207.390 ;
        RECT 2193.840 207.070 2194.100 207.390 ;
        RECT 2193.900 16.650 2194.040 207.070 ;
        RECT 2193.840 16.330 2194.100 16.650 ;
        RECT 2393.480 15.990 2393.740 16.310 ;
        RECT 2393.540 2.400 2393.680 15.990 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2346.145 14.705 2346.315 17.255 ;
      LAYER mcon ;
        RECT 2346.145 17.085 2346.315 17.255 ;
      LAYER met1 ;
        RECT 2203.470 208.320 2203.790 208.380 ;
        RECT 2342.390 208.320 2342.710 208.380 ;
        RECT 2203.470 208.180 2342.710 208.320 ;
        RECT 2203.470 208.120 2203.790 208.180 ;
        RECT 2342.390 208.120 2342.710 208.180 ;
        RECT 2342.390 17.240 2342.710 17.300 ;
        RECT 2346.085 17.240 2346.375 17.285 ;
        RECT 2342.390 17.100 2346.375 17.240 ;
        RECT 2342.390 17.040 2342.710 17.100 ;
        RECT 2346.085 17.055 2346.375 17.100 ;
        RECT 2346.085 14.860 2346.375 14.905 ;
        RECT 2411.390 14.860 2411.710 14.920 ;
        RECT 2346.085 14.720 2411.710 14.860 ;
        RECT 2346.085 14.675 2346.375 14.720 ;
        RECT 2411.390 14.660 2411.710 14.720 ;
      LAYER via ;
        RECT 2203.500 208.120 2203.760 208.380 ;
        RECT 2342.420 208.120 2342.680 208.380 ;
        RECT 2342.420 17.040 2342.680 17.300 ;
        RECT 2411.420 14.660 2411.680 14.920 ;
      LAYER met2 ;
        RECT 2203.540 220.000 2203.820 224.000 ;
        RECT 2203.560 208.410 2203.700 220.000 ;
        RECT 2203.500 208.090 2203.760 208.410 ;
        RECT 2342.420 208.090 2342.680 208.410 ;
        RECT 2342.480 17.330 2342.620 208.090 ;
        RECT 2342.420 17.010 2342.680 17.330 ;
        RECT 2411.420 14.630 2411.680 14.950 ;
        RECT 2411.480 2.400 2411.620 14.630 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 806.910 208.660 807.230 208.720 ;
        RECT 880.970 208.660 881.290 208.720 ;
        RECT 806.910 208.520 881.290 208.660 ;
        RECT 806.910 208.460 807.230 208.520 ;
        RECT 880.970 208.460 881.290 208.520 ;
      LAYER via ;
        RECT 806.940 208.460 807.200 208.720 ;
        RECT 881.000 208.460 881.260 208.720 ;
      LAYER met2 ;
        RECT 881.040 220.000 881.320 224.000 ;
        RECT 881.060 208.750 881.200 220.000 ;
        RECT 806.940 208.430 807.200 208.750 ;
        RECT 881.000 208.430 881.260 208.750 ;
        RECT 807.000 17.410 807.140 208.430 ;
        RECT 805.620 17.270 807.140 17.410 ;
        RECT 805.620 2.400 805.760 17.270 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 17.580 3.150 17.640 ;
        RECT 2.830 17.440 197.180 17.580 ;
        RECT 2.830 17.380 3.150 17.440 ;
        RECT 197.040 17.240 197.180 17.440 ;
        RECT 214.430 17.240 214.750 17.300 ;
        RECT 197.040 17.100 214.750 17.240 ;
        RECT 214.430 17.040 214.750 17.100 ;
      LAYER via ;
        RECT 2.860 17.380 3.120 17.640 ;
        RECT 214.460 17.040 214.720 17.300 ;
      LAYER met2 ;
        RECT 220.020 220.730 220.300 224.000 ;
        RECT 214.520 220.590 220.300 220.730 ;
        RECT 2.860 17.350 3.120 17.670 ;
        RECT 2.920 2.400 3.060 17.350 ;
        RECT 214.520 17.330 214.660 220.590 ;
        RECT 220.020 220.000 220.300 220.590 ;
        RECT 214.460 17.010 214.720 17.330 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 17.240 8.670 17.300 ;
        RECT 8.350 17.100 179.700 17.240 ;
        RECT 8.350 17.040 8.670 17.100 ;
        RECT 179.560 16.220 179.700 17.100 ;
        RECT 221.330 16.220 221.650 16.280 ;
        RECT 179.560 16.080 221.650 16.220 ;
        RECT 221.330 16.020 221.650 16.080 ;
      LAYER via ;
        RECT 8.380 17.040 8.640 17.300 ;
        RECT 221.360 16.020 221.620 16.280 ;
      LAYER met2 ;
        RECT 224.620 220.730 224.900 224.000 ;
        RECT 221.420 220.590 224.900 220.730 ;
        RECT 8.380 17.010 8.640 17.330 ;
        RECT 8.440 2.400 8.580 17.010 ;
        RECT 221.420 16.310 221.560 220.590 ;
        RECT 224.620 220.000 224.900 220.590 ;
        RECT 221.360 15.990 221.620 16.310 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 110.100 18.460 134.620 18.600 ;
        RECT 14.330 17.920 14.650 17.980 ;
        RECT 110.100 17.920 110.240 18.460 ;
        RECT 14.330 17.780 110.240 17.920 ;
        RECT 134.480 17.920 134.620 18.460 ;
        RECT 228.230 18.260 228.550 18.320 ;
        RECT 203.480 18.120 228.550 18.260 ;
        RECT 203.480 17.920 203.620 18.120 ;
        RECT 228.230 18.060 228.550 18.120 ;
        RECT 134.480 17.780 203.620 17.920 ;
        RECT 14.330 17.720 14.650 17.780 ;
      LAYER via ;
        RECT 14.360 17.720 14.620 17.980 ;
        RECT 228.260 18.060 228.520 18.320 ;
      LAYER met2 ;
        RECT 229.680 220.730 229.960 224.000 ;
        RECT 228.320 220.590 229.960 220.730 ;
        RECT 228.320 18.350 228.460 220.590 ;
        RECT 229.680 220.000 229.960 220.590 ;
        RECT 228.260 18.030 228.520 18.350 ;
        RECT 14.360 17.690 14.620 18.010 ;
        RECT 14.420 2.400 14.560 17.690 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 24.040 38.570 24.100 ;
        RECT 248.930 24.040 249.250 24.100 ;
        RECT 38.250 23.900 249.250 24.040 ;
        RECT 38.250 23.840 38.570 23.900 ;
        RECT 248.930 23.840 249.250 23.900 ;
      LAYER via ;
        RECT 38.280 23.840 38.540 24.100 ;
        RECT 248.960 23.840 249.220 24.100 ;
      LAYER met2 ;
        RECT 249.000 220.000 249.280 224.000 ;
        RECT 249.020 24.130 249.160 220.000 ;
        RECT 38.280 23.810 38.540 24.130 ;
        RECT 248.960 23.810 249.220 24.130 ;
        RECT 38.340 2.400 38.480 23.810 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 240.650 16.900 240.970 16.960 ;
        RECT 414.990 16.900 415.310 16.960 ;
        RECT 240.650 16.760 415.310 16.900 ;
        RECT 240.650 16.700 240.970 16.760 ;
        RECT 414.990 16.700 415.310 16.760 ;
      LAYER via ;
        RECT 240.680 16.700 240.940 16.960 ;
        RECT 415.020 16.700 415.280 16.960 ;
      LAYER met2 ;
        RECT 415.520 220.730 415.800 224.000 ;
        RECT 415.080 220.590 415.800 220.730 ;
        RECT 415.080 16.990 415.220 220.590 ;
        RECT 415.520 220.000 415.800 220.590 ;
        RECT 240.680 16.670 240.940 16.990 ;
        RECT 415.020 16.670 415.280 16.990 ;
        RECT 240.740 2.400 240.880 16.670 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 412.305 16.405 412.475 17.935 ;
      LAYER mcon ;
        RECT 412.305 17.765 412.475 17.935 ;
      LAYER met1 ;
        RECT 412.245 17.920 412.535 17.965 ;
        RECT 376.440 17.780 412.535 17.920 ;
        RECT 258.130 17.580 258.450 17.640 ;
        RECT 376.440 17.580 376.580 17.780 ;
        RECT 412.245 17.735 412.535 17.780 ;
        RECT 258.130 17.440 376.580 17.580 ;
        RECT 258.130 17.380 258.450 17.440 ;
        RECT 428.330 16.900 428.650 16.960 ;
        RECT 415.540 16.760 428.650 16.900 ;
        RECT 412.245 16.560 412.535 16.605 ;
        RECT 415.540 16.560 415.680 16.760 ;
        RECT 428.330 16.700 428.650 16.760 ;
        RECT 412.245 16.420 415.680 16.560 ;
        RECT 412.245 16.375 412.535 16.420 ;
      LAYER via ;
        RECT 258.160 17.380 258.420 17.640 ;
        RECT 428.360 16.700 428.620 16.960 ;
      LAYER met2 ;
        RECT 430.240 220.730 430.520 224.000 ;
        RECT 428.420 220.590 430.520 220.730 ;
        RECT 258.160 17.350 258.420 17.670 ;
        RECT 258.220 2.400 258.360 17.350 ;
        RECT 428.420 16.990 428.560 220.590 ;
        RECT 430.240 220.000 430.520 220.590 ;
        RECT 428.360 16.670 428.620 16.990 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 412.765 17.765 412.935 19.295 ;
      LAYER mcon ;
        RECT 412.765 19.125 412.935 19.295 ;
      LAYER met1 ;
        RECT 276.070 19.280 276.390 19.340 ;
        RECT 412.705 19.280 412.995 19.325 ;
        RECT 276.070 19.140 412.995 19.280 ;
        RECT 276.070 19.080 276.390 19.140 ;
        RECT 412.705 19.095 412.995 19.140 ;
        RECT 412.705 17.920 412.995 17.965 ;
        RECT 441.670 17.920 441.990 17.980 ;
        RECT 412.705 17.780 441.990 17.920 ;
        RECT 412.705 17.735 412.995 17.780 ;
        RECT 441.670 17.720 441.990 17.780 ;
      LAYER via ;
        RECT 276.100 19.080 276.360 19.340 ;
        RECT 441.700 17.720 441.960 17.980 ;
      LAYER met2 ;
        RECT 444.960 220.730 445.240 224.000 ;
        RECT 441.760 220.590 445.240 220.730 ;
        RECT 276.100 19.050 276.360 19.370 ;
        RECT 276.160 2.400 276.300 19.050 ;
        RECT 441.760 18.010 441.900 220.590 ;
        RECT 444.960 220.000 445.240 220.590 ;
        RECT 441.700 17.690 441.960 18.010 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 18.260 294.330 18.320 ;
        RECT 455.470 18.260 455.790 18.320 ;
        RECT 294.010 18.120 455.790 18.260 ;
        RECT 294.010 18.060 294.330 18.120 ;
        RECT 455.470 18.060 455.790 18.120 ;
      LAYER via ;
        RECT 294.040 18.060 294.300 18.320 ;
        RECT 455.500 18.060 455.760 18.320 ;
      LAYER met2 ;
        RECT 459.680 220.730 459.960 224.000 ;
        RECT 455.560 220.590 459.960 220.730 ;
        RECT 455.560 18.350 455.700 220.590 ;
        RECT 459.680 220.000 459.960 220.590 ;
        RECT 294.040 18.030 294.300 18.350 ;
        RECT 455.500 18.030 455.760 18.350 ;
        RECT 294.100 2.400 294.240 18.030 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 19.620 312.270 19.680 ;
        RECT 469.730 19.620 470.050 19.680 ;
        RECT 311.950 19.480 470.050 19.620 ;
        RECT 311.950 19.420 312.270 19.480 ;
        RECT 469.730 19.420 470.050 19.480 ;
      LAYER via ;
        RECT 311.980 19.420 312.240 19.680 ;
        RECT 469.760 19.420 470.020 19.680 ;
      LAYER met2 ;
        RECT 474.400 220.730 474.680 224.000 ;
        RECT 469.820 220.590 474.680 220.730 ;
        RECT 469.820 19.710 469.960 220.590 ;
        RECT 474.400 220.000 474.680 220.590 ;
        RECT 311.980 19.390 312.240 19.710 ;
        RECT 469.760 19.390 470.020 19.710 ;
        RECT 312.040 2.400 312.180 19.390 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 483.070 145.080 483.390 145.140 ;
        RECT 487.670 145.080 487.990 145.140 ;
        RECT 483.070 144.940 487.990 145.080 ;
        RECT 483.070 144.880 483.390 144.940 ;
        RECT 487.670 144.880 487.990 144.940 ;
        RECT 483.070 96.800 483.390 96.860 ;
        RECT 483.530 96.800 483.850 96.860 ;
        RECT 483.070 96.660 483.850 96.800 ;
        RECT 483.070 96.600 483.390 96.660 ;
        RECT 483.530 96.600 483.850 96.660 ;
        RECT 329.890 19.960 330.210 20.020 ;
        RECT 483.990 19.960 484.310 20.020 ;
        RECT 329.890 19.820 484.310 19.960 ;
        RECT 329.890 19.760 330.210 19.820 ;
        RECT 483.990 19.760 484.310 19.820 ;
      LAYER via ;
        RECT 483.100 144.880 483.360 145.140 ;
        RECT 487.700 144.880 487.960 145.140 ;
        RECT 483.100 96.600 483.360 96.860 ;
        RECT 483.560 96.600 483.820 96.860 ;
        RECT 329.920 19.760 330.180 20.020 ;
        RECT 484.020 19.760 484.280 20.020 ;
      LAYER met2 ;
        RECT 489.120 220.730 489.400 224.000 ;
        RECT 487.760 220.590 489.400 220.730 ;
        RECT 487.760 145.170 487.900 220.590 ;
        RECT 489.120 220.000 489.400 220.590 ;
        RECT 483.100 144.850 483.360 145.170 ;
        RECT 487.700 144.850 487.960 145.170 ;
        RECT 483.160 96.890 483.300 144.850 ;
        RECT 483.100 96.570 483.360 96.890 ;
        RECT 483.560 96.570 483.820 96.890 ;
        RECT 483.620 96.290 483.760 96.570 ;
        RECT 483.620 96.150 484.220 96.290 ;
        RECT 484.080 20.050 484.220 96.150 ;
        RECT 329.920 19.730 330.180 20.050 ;
        RECT 484.020 19.730 484.280 20.050 ;
        RECT 329.980 2.400 330.120 19.730 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 20.300 347.690 20.360 ;
        RECT 504.230 20.300 504.550 20.360 ;
        RECT 347.370 20.160 504.550 20.300 ;
        RECT 347.370 20.100 347.690 20.160 ;
        RECT 504.230 20.100 504.550 20.160 ;
      LAYER via ;
        RECT 347.400 20.100 347.660 20.360 ;
        RECT 504.260 20.100 504.520 20.360 ;
      LAYER met2 ;
        RECT 503.840 220.730 504.120 224.000 ;
        RECT 503.840 220.590 504.460 220.730 ;
        RECT 503.840 220.000 504.120 220.590 ;
        RECT 504.320 20.390 504.460 220.590 ;
        RECT 347.400 20.070 347.660 20.390 ;
        RECT 504.260 20.070 504.520 20.390 ;
        RECT 347.460 2.400 347.600 20.070 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 24.040 365.630 24.100 ;
        RECT 518.030 24.040 518.350 24.100 ;
        RECT 365.310 23.900 518.350 24.040 ;
        RECT 365.310 23.840 365.630 23.900 ;
        RECT 518.030 23.840 518.350 23.900 ;
      LAYER via ;
        RECT 365.340 23.840 365.600 24.100 ;
        RECT 518.060 23.840 518.320 24.100 ;
      LAYER met2 ;
        RECT 518.560 220.730 518.840 224.000 ;
        RECT 518.120 220.590 518.840 220.730 ;
        RECT 518.120 24.130 518.260 220.590 ;
        RECT 518.560 220.000 518.840 220.590 ;
        RECT 365.340 23.810 365.600 24.130 ;
        RECT 518.060 23.810 518.320 24.130 ;
        RECT 365.400 2.400 365.540 23.810 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 18.600 383.570 18.660 ;
        RECT 531.370 18.600 531.690 18.660 ;
        RECT 383.250 18.460 531.690 18.600 ;
        RECT 383.250 18.400 383.570 18.460 ;
        RECT 531.370 18.400 531.690 18.460 ;
      LAYER via ;
        RECT 383.280 18.400 383.540 18.660 ;
        RECT 531.400 18.400 531.660 18.660 ;
      LAYER met2 ;
        RECT 533.280 220.730 533.560 224.000 ;
        RECT 531.460 220.590 533.560 220.730 ;
        RECT 531.460 18.690 531.600 220.590 ;
        RECT 533.280 220.000 533.560 220.590 ;
        RECT 383.280 18.370 383.540 18.690 ;
        RECT 531.400 18.370 531.660 18.690 ;
        RECT 383.340 2.400 383.480 18.370 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 18.940 401.510 19.000 ;
        RECT 545.170 18.940 545.490 19.000 ;
        RECT 401.190 18.800 545.490 18.940 ;
        RECT 401.190 18.740 401.510 18.800 ;
        RECT 545.170 18.740 545.490 18.800 ;
      LAYER via ;
        RECT 401.220 18.740 401.480 19.000 ;
        RECT 545.200 18.740 545.460 19.000 ;
      LAYER met2 ;
        RECT 548.000 220.730 548.280 224.000 ;
        RECT 545.260 220.590 548.280 220.730 ;
        RECT 545.260 19.030 545.400 220.590 ;
        RECT 548.000 220.000 548.280 220.590 ;
        RECT 401.220 18.710 401.480 19.030 ;
        RECT 545.200 18.710 545.460 19.030 ;
        RECT 401.280 2.400 401.420 18.710 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 266.485 144.925 266.655 193.035 ;
      LAYER mcon ;
        RECT 266.485 192.865 266.655 193.035 ;
      LAYER met1 ;
        RECT 266.425 193.020 266.715 193.065 ;
        RECT 266.870 193.020 267.190 193.080 ;
        RECT 266.425 192.880 267.190 193.020 ;
        RECT 266.425 192.835 266.715 192.880 ;
        RECT 266.870 192.820 267.190 192.880 ;
        RECT 266.410 145.080 266.730 145.140 ;
        RECT 266.215 144.940 266.730 145.080 ;
        RECT 266.410 144.880 266.730 144.940 ;
        RECT 262.730 110.740 263.050 110.800 ;
        RECT 266.410 110.740 266.730 110.800 ;
        RECT 262.730 110.600 266.730 110.740 ;
        RECT 262.730 110.540 263.050 110.600 ;
        RECT 266.410 110.540 266.730 110.600 ;
        RECT 62.170 24.380 62.490 24.440 ;
        RECT 263.190 24.380 263.510 24.440 ;
        RECT 62.170 24.240 263.510 24.380 ;
        RECT 62.170 24.180 62.490 24.240 ;
        RECT 263.190 24.180 263.510 24.240 ;
      LAYER via ;
        RECT 266.900 192.820 267.160 193.080 ;
        RECT 266.440 144.880 266.700 145.140 ;
        RECT 262.760 110.540 263.020 110.800 ;
        RECT 266.440 110.540 266.700 110.800 ;
        RECT 62.200 24.180 62.460 24.440 ;
        RECT 263.220 24.180 263.480 24.440 ;
      LAYER met2 ;
        RECT 268.780 220.730 269.060 224.000 ;
        RECT 266.960 220.590 269.060 220.730 ;
        RECT 266.960 193.110 267.100 220.590 ;
        RECT 268.780 220.000 269.060 220.590 ;
        RECT 266.900 192.790 267.160 193.110 ;
        RECT 266.440 144.850 266.700 145.170 ;
        RECT 266.500 110.830 266.640 144.850 ;
        RECT 262.760 110.510 263.020 110.830 ;
        RECT 266.440 110.510 266.700 110.830 ;
        RECT 262.820 62.290 262.960 110.510 ;
        RECT 262.820 62.150 263.420 62.290 ;
        RECT 263.280 24.470 263.420 62.150 ;
        RECT 62.200 24.150 62.460 24.470 ;
        RECT 263.220 24.150 263.480 24.470 ;
        RECT 62.260 2.400 62.400 24.150 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 471.660 17.100 521.020 17.240 ;
        RECT 419.130 16.560 419.450 16.620 ;
        RECT 471.660 16.560 471.800 17.100 ;
        RECT 520.880 16.900 521.020 17.100 ;
        RECT 559.430 16.900 559.750 16.960 ;
        RECT 520.880 16.760 559.750 16.900 ;
        RECT 559.430 16.700 559.750 16.760 ;
        RECT 419.130 16.420 471.800 16.560 ;
        RECT 419.130 16.360 419.450 16.420 ;
      LAYER via ;
        RECT 419.160 16.360 419.420 16.620 ;
        RECT 559.460 16.700 559.720 16.960 ;
      LAYER met2 ;
        RECT 562.720 220.730 563.000 224.000 ;
        RECT 559.520 220.590 563.000 220.730 ;
        RECT 559.520 16.990 559.660 220.590 ;
        RECT 562.720 220.000 563.000 220.590 ;
        RECT 559.460 16.670 559.720 16.990 ;
        RECT 419.160 16.330 419.420 16.650 ;
        RECT 419.220 2.400 419.360 16.330 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 573.230 17.580 573.550 17.640 ;
        RECT 456.020 17.440 573.550 17.580 ;
        RECT 456.020 17.240 456.160 17.440 ;
        RECT 573.230 17.380 573.550 17.440 ;
        RECT 449.120 17.100 456.160 17.240 ;
        RECT 436.610 16.900 436.930 16.960 ;
        RECT 449.120 16.900 449.260 17.100 ;
        RECT 436.610 16.760 449.260 16.900 ;
        RECT 436.610 16.700 436.930 16.760 ;
      LAYER via ;
        RECT 573.260 17.380 573.520 17.640 ;
        RECT 436.640 16.700 436.900 16.960 ;
      LAYER met2 ;
        RECT 577.440 220.730 577.720 224.000 ;
        RECT 573.320 220.590 577.720 220.730 ;
        RECT 573.320 17.670 573.460 220.590 ;
        RECT 577.440 220.000 577.720 220.590 ;
        RECT 573.260 17.350 573.520 17.670 ;
        RECT 436.640 16.670 436.900 16.990 ;
        RECT 436.700 2.400 436.840 16.670 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 588.485 48.365 588.655 137.955 ;
      LAYER mcon ;
        RECT 588.485 137.785 588.655 137.955 ;
      LAYER met1 ;
        RECT 587.030 137.940 587.350 138.000 ;
        RECT 588.425 137.940 588.715 137.985 ;
        RECT 587.030 137.800 588.715 137.940 ;
        RECT 587.030 137.740 587.350 137.800 ;
        RECT 588.425 137.755 588.715 137.800 ;
        RECT 588.410 48.520 588.730 48.580 ;
        RECT 588.215 48.380 588.730 48.520 ;
        RECT 588.410 48.320 588.730 48.380 ;
        RECT 588.410 17.920 588.730 17.980 ;
        RECT 455.560 17.780 588.730 17.920 ;
        RECT 454.550 17.580 454.870 17.640 ;
        RECT 455.560 17.580 455.700 17.780 ;
        RECT 588.410 17.720 588.730 17.780 ;
        RECT 454.550 17.440 455.700 17.580 ;
        RECT 454.550 17.380 454.870 17.440 ;
      LAYER via ;
        RECT 587.060 137.740 587.320 138.000 ;
        RECT 588.440 48.320 588.700 48.580 ;
        RECT 454.580 17.380 454.840 17.640 ;
        RECT 588.440 17.720 588.700 17.980 ;
      LAYER met2 ;
        RECT 592.160 220.730 592.440 224.000 ;
        RECT 590.800 220.590 592.440 220.730 ;
        RECT 590.800 146.045 590.940 220.590 ;
        RECT 592.160 220.000 592.440 220.590 ;
        RECT 590.730 145.675 591.010 146.045 ;
        RECT 587.050 144.995 587.330 145.365 ;
        RECT 587.120 138.030 587.260 144.995 ;
        RECT 587.060 137.710 587.320 138.030 ;
        RECT 588.440 48.290 588.700 48.610 ;
        RECT 588.500 18.010 588.640 48.290 ;
        RECT 588.440 17.690 588.700 18.010 ;
        RECT 454.580 17.350 454.840 17.670 ;
        RECT 454.640 2.400 454.780 17.350 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 590.730 145.720 591.010 146.000 ;
        RECT 587.050 145.040 587.330 145.320 ;
      LAYER met3 ;
        RECT 590.705 146.010 591.035 146.025 ;
        RECT 586.350 145.710 591.035 146.010 ;
        RECT 586.350 145.330 586.650 145.710 ;
        RECT 590.705 145.695 591.035 145.710 ;
        RECT 587.025 145.330 587.355 145.345 ;
        RECT 586.350 145.030 587.355 145.330 ;
        RECT 587.025 145.015 587.355 145.030 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 602.285 61.965 602.455 137.955 ;
        RECT 579.745 18.445 579.915 22.015 ;
      LAYER mcon ;
        RECT 602.285 137.785 602.455 137.955 ;
        RECT 579.745 21.845 579.915 22.015 ;
      LAYER met1 ;
        RECT 600.830 137.940 601.150 138.000 ;
        RECT 602.225 137.940 602.515 137.985 ;
        RECT 600.830 137.800 602.515 137.940 ;
        RECT 600.830 137.740 601.150 137.800 ;
        RECT 602.225 137.755 602.515 137.800 ;
        RECT 602.210 62.120 602.530 62.180 ;
        RECT 602.015 61.980 602.530 62.120 ;
        RECT 602.210 61.920 602.530 61.980 ;
        RECT 579.685 22.000 579.975 22.045 ;
        RECT 602.210 22.000 602.530 22.060 ;
        RECT 579.685 21.860 602.530 22.000 ;
        RECT 579.685 21.815 579.975 21.860 ;
        RECT 602.210 21.800 602.530 21.860 ;
        RECT 579.685 18.600 579.975 18.645 ;
        RECT 531.920 18.460 579.975 18.600 ;
        RECT 472.490 18.260 472.810 18.320 ;
        RECT 531.920 18.260 532.060 18.460 ;
        RECT 579.685 18.415 579.975 18.460 ;
        RECT 472.490 18.120 532.060 18.260 ;
        RECT 472.490 18.060 472.810 18.120 ;
      LAYER via ;
        RECT 600.860 137.740 601.120 138.000 ;
        RECT 602.240 61.920 602.500 62.180 ;
        RECT 602.240 21.800 602.500 22.060 ;
        RECT 472.520 18.060 472.780 18.320 ;
      LAYER met2 ;
        RECT 606.880 220.730 607.160 224.000 ;
        RECT 605.520 220.590 607.160 220.730 ;
        RECT 605.520 139.245 605.660 220.590 ;
        RECT 606.880 220.000 607.160 220.590 ;
        RECT 605.450 138.875 605.730 139.245 ;
        RECT 600.850 138.195 601.130 138.565 ;
        RECT 600.920 138.030 601.060 138.195 ;
        RECT 600.860 137.710 601.120 138.030 ;
        RECT 602.240 61.890 602.500 62.210 ;
        RECT 602.300 22.090 602.440 61.890 ;
        RECT 602.240 21.770 602.500 22.090 ;
        RECT 472.520 18.030 472.780 18.350 ;
        RECT 472.580 2.400 472.720 18.030 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 605.450 138.920 605.730 139.200 ;
        RECT 600.850 138.240 601.130 138.520 ;
      LAYER met3 ;
        RECT 605.425 139.210 605.755 139.225 ;
        RECT 600.150 138.910 605.755 139.210 ;
        RECT 600.150 138.530 600.450 138.910 ;
        RECT 605.425 138.895 605.755 138.910 ;
        RECT 600.825 138.530 601.155 138.545 ;
        RECT 600.150 138.230 601.155 138.530 ;
        RECT 600.825 138.215 601.155 138.230 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 490.430 19.620 490.750 19.680 ;
        RECT 621.530 19.620 621.850 19.680 ;
        RECT 490.430 19.480 621.850 19.620 ;
        RECT 490.430 19.420 490.750 19.480 ;
        RECT 621.530 19.420 621.850 19.480 ;
      LAYER via ;
        RECT 490.460 19.420 490.720 19.680 ;
        RECT 621.560 19.420 621.820 19.680 ;
      LAYER met2 ;
        RECT 621.600 220.000 621.880 224.000 ;
        RECT 621.620 19.710 621.760 220.000 ;
        RECT 490.460 19.390 490.720 19.710 ;
        RECT 621.560 19.390 621.820 19.710 ;
        RECT 490.520 2.400 490.660 19.390 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 19.280 508.230 19.340 ;
        RECT 635.330 19.280 635.650 19.340 ;
        RECT 507.910 19.140 635.650 19.280 ;
        RECT 507.910 19.080 508.230 19.140 ;
        RECT 635.330 19.080 635.650 19.140 ;
      LAYER via ;
        RECT 507.940 19.080 508.200 19.340 ;
        RECT 635.360 19.080 635.620 19.340 ;
      LAYER met2 ;
        RECT 635.860 220.730 636.140 224.000 ;
        RECT 635.420 220.590 636.140 220.730 ;
        RECT 635.420 19.370 635.560 220.590 ;
        RECT 635.860 220.000 636.140 220.590 ;
        RECT 507.940 19.050 508.200 19.370 ;
        RECT 635.360 19.050 635.620 19.370 ;
        RECT 508.000 2.400 508.140 19.050 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 565.945 208.845 566.115 210.715 ;
        RECT 585.265 210.545 585.435 212.075 ;
        RECT 602.285 211.225 602.455 212.415 ;
        RECT 613.325 211.225 613.955 211.395 ;
        RECT 613.785 208.845 613.955 211.225 ;
        RECT 620.225 207.825 620.395 209.015 ;
      LAYER mcon ;
        RECT 602.285 212.245 602.455 212.415 ;
        RECT 585.265 211.905 585.435 212.075 ;
        RECT 565.945 210.545 566.115 210.715 ;
        RECT 620.225 208.845 620.395 209.015 ;
      LAYER met1 ;
        RECT 602.225 212.400 602.515 212.445 ;
        RECT 597.240 212.260 602.515 212.400 ;
        RECT 585.205 212.060 585.495 212.105 ;
        RECT 597.240 212.060 597.380 212.260 ;
        RECT 602.225 212.215 602.515 212.260 ;
        RECT 585.205 211.920 597.380 212.060 ;
        RECT 585.205 211.875 585.495 211.920 ;
        RECT 602.225 211.380 602.515 211.425 ;
        RECT 613.265 211.380 613.555 211.425 ;
        RECT 602.225 211.240 613.555 211.380 ;
        RECT 602.225 211.195 602.515 211.240 ;
        RECT 613.265 211.195 613.555 211.240 ;
        RECT 565.885 210.700 566.175 210.745 ;
        RECT 585.205 210.700 585.495 210.745 ;
        RECT 565.885 210.560 585.495 210.700 ;
        RECT 565.885 210.515 566.175 210.560 ;
        RECT 585.205 210.515 585.495 210.560 ;
        RECT 530.910 209.000 531.230 209.060 ;
        RECT 565.885 209.000 566.175 209.045 ;
        RECT 530.910 208.860 566.175 209.000 ;
        RECT 530.910 208.800 531.230 208.860 ;
        RECT 565.885 208.815 566.175 208.860 ;
        RECT 613.725 209.000 614.015 209.045 ;
        RECT 620.165 209.000 620.455 209.045 ;
        RECT 613.725 208.860 620.455 209.000 ;
        RECT 613.725 208.815 614.015 208.860 ;
        RECT 620.165 208.815 620.455 208.860 ;
        RECT 650.510 208.320 650.830 208.380 ;
        RECT 638.640 208.180 650.830 208.320 ;
        RECT 620.165 207.980 620.455 208.025 ;
        RECT 638.640 207.980 638.780 208.180 ;
        RECT 650.510 208.120 650.830 208.180 ;
        RECT 620.165 207.840 638.780 207.980 ;
        RECT 620.165 207.795 620.455 207.840 ;
        RECT 525.850 17.240 526.170 17.300 ;
        RECT 530.910 17.240 531.230 17.300 ;
        RECT 525.850 17.100 531.230 17.240 ;
        RECT 525.850 17.040 526.170 17.100 ;
        RECT 530.910 17.040 531.230 17.100 ;
      LAYER via ;
        RECT 530.940 208.800 531.200 209.060 ;
        RECT 650.540 208.120 650.800 208.380 ;
        RECT 525.880 17.040 526.140 17.300 ;
        RECT 530.940 17.040 531.200 17.300 ;
      LAYER met2 ;
        RECT 650.580 220.000 650.860 224.000 ;
        RECT 530.940 208.770 531.200 209.090 ;
        RECT 531.000 17.330 531.140 208.770 ;
        RECT 650.600 208.410 650.740 220.000 ;
        RECT 650.540 208.090 650.800 208.410 ;
        RECT 525.880 17.010 526.140 17.330 ;
        RECT 530.940 17.010 531.200 17.330 ;
        RECT 525.940 2.400 526.080 17.010 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 544.785 193.205 544.955 210.035 ;
        RECT 544.785 144.925 544.955 192.695 ;
        RECT 543.865 2.805 544.035 48.195 ;
      LAYER mcon ;
        RECT 544.785 209.865 544.955 210.035 ;
        RECT 544.785 192.525 544.955 192.695 ;
        RECT 543.865 48.025 544.035 48.195 ;
      LAYER met1 ;
        RECT 544.725 210.020 545.015 210.065 ;
        RECT 665.230 210.020 665.550 210.080 ;
        RECT 544.725 209.880 665.550 210.020 ;
        RECT 544.725 209.835 545.015 209.880 ;
        RECT 665.230 209.820 665.550 209.880 ;
        RECT 544.710 193.360 545.030 193.420 ;
        RECT 544.515 193.220 545.030 193.360 ;
        RECT 544.710 193.160 545.030 193.220 ;
        RECT 544.710 192.680 545.030 192.740 ;
        RECT 544.515 192.540 545.030 192.680 ;
        RECT 544.710 192.480 545.030 192.540 ;
        RECT 544.710 145.080 545.030 145.140 ;
        RECT 544.515 144.940 545.030 145.080 ;
        RECT 544.710 144.880 545.030 144.940 ;
        RECT 543.790 96.460 544.110 96.520 ;
        RECT 544.710 96.460 545.030 96.520 ;
        RECT 543.790 96.320 545.030 96.460 ;
        RECT 543.790 96.260 544.110 96.320 ;
        RECT 544.710 96.260 545.030 96.320 ;
        RECT 543.805 48.180 544.095 48.225 ;
        RECT 544.710 48.180 545.030 48.240 ;
        RECT 543.805 48.040 545.030 48.180 ;
        RECT 543.805 47.995 544.095 48.040 ;
        RECT 544.710 47.980 545.030 48.040 ;
        RECT 543.790 2.960 544.110 3.020 ;
        RECT 543.595 2.820 544.110 2.960 ;
        RECT 543.790 2.760 544.110 2.820 ;
      LAYER via ;
        RECT 665.260 209.820 665.520 210.080 ;
        RECT 544.740 193.160 545.000 193.420 ;
        RECT 544.740 192.480 545.000 192.740 ;
        RECT 544.740 144.880 545.000 145.140 ;
        RECT 543.820 96.260 544.080 96.520 ;
        RECT 544.740 96.260 545.000 96.520 ;
        RECT 544.740 47.980 545.000 48.240 ;
        RECT 543.820 2.760 544.080 3.020 ;
      LAYER met2 ;
        RECT 665.300 220.000 665.580 224.000 ;
        RECT 665.320 210.110 665.460 220.000 ;
        RECT 665.260 209.790 665.520 210.110 ;
        RECT 544.740 193.130 545.000 193.450 ;
        RECT 544.800 192.770 544.940 193.130 ;
        RECT 544.740 192.450 545.000 192.770 ;
        RECT 544.740 144.850 545.000 145.170 ;
        RECT 544.800 96.550 544.940 144.850 ;
        RECT 543.820 96.230 544.080 96.550 ;
        RECT 544.740 96.230 545.000 96.550 ;
        RECT 543.880 48.805 544.020 96.230 ;
        RECT 543.810 48.435 544.090 48.805 ;
        RECT 544.730 48.435 545.010 48.805 ;
        RECT 544.800 48.270 544.940 48.435 ;
        RECT 544.740 47.950 545.000 48.270 ;
        RECT 543.820 2.730 544.080 3.050 ;
        RECT 543.880 2.400 544.020 2.730 ;
        RECT 543.670 -4.800 544.230 2.400 ;
      LAYER via2 ;
        RECT 543.810 48.480 544.090 48.760 ;
        RECT 544.730 48.480 545.010 48.760 ;
      LAYER met3 ;
        RECT 543.785 48.770 544.115 48.785 ;
        RECT 544.705 48.770 545.035 48.785 ;
        RECT 543.785 48.470 545.035 48.770 ;
        RECT 543.785 48.455 544.115 48.470 ;
        RECT 544.705 48.455 545.035 48.470 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 565.410 207.300 565.730 207.360 ;
        RECT 679.950 207.300 680.270 207.360 ;
        RECT 565.410 207.160 680.270 207.300 ;
        RECT 565.410 207.100 565.730 207.160 ;
        RECT 679.950 207.100 680.270 207.160 ;
        RECT 561.730 20.640 562.050 20.700 ;
        RECT 565.410 20.640 565.730 20.700 ;
        RECT 561.730 20.500 565.730 20.640 ;
        RECT 561.730 20.440 562.050 20.500 ;
        RECT 565.410 20.440 565.730 20.500 ;
      LAYER via ;
        RECT 565.440 207.100 565.700 207.360 ;
        RECT 679.980 207.100 680.240 207.360 ;
        RECT 561.760 20.440 562.020 20.700 ;
        RECT 565.440 20.440 565.700 20.700 ;
      LAYER met2 ;
        RECT 680.020 220.000 680.300 224.000 ;
        RECT 680.040 207.390 680.180 220.000 ;
        RECT 565.440 207.070 565.700 207.390 ;
        RECT 679.980 207.070 680.240 207.390 ;
        RECT 565.500 20.730 565.640 207.070 ;
        RECT 561.760 20.410 562.020 20.730 ;
        RECT 565.440 20.410 565.700 20.730 ;
        RECT 561.820 2.400 561.960 20.410 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 612.405 210.205 612.575 212.415 ;
      LAYER mcon ;
        RECT 612.405 212.245 612.575 212.415 ;
      LAYER met1 ;
        RECT 612.345 212.400 612.635 212.445 ;
        RECT 694.670 212.400 694.990 212.460 ;
        RECT 612.345 212.260 694.990 212.400 ;
        RECT 612.345 212.215 612.635 212.260 ;
        RECT 694.670 212.200 694.990 212.260 ;
        RECT 586.110 210.360 586.430 210.420 ;
        RECT 612.345 210.360 612.635 210.405 ;
        RECT 586.110 210.220 612.635 210.360 ;
        RECT 586.110 210.160 586.430 210.220 ;
        RECT 612.345 210.175 612.635 210.220 ;
        RECT 579.670 20.640 579.990 20.700 ;
        RECT 586.110 20.640 586.430 20.700 ;
        RECT 579.670 20.500 586.430 20.640 ;
        RECT 579.670 20.440 579.990 20.500 ;
        RECT 586.110 20.440 586.430 20.500 ;
      LAYER via ;
        RECT 694.700 212.200 694.960 212.460 ;
        RECT 586.140 210.160 586.400 210.420 ;
        RECT 579.700 20.440 579.960 20.700 ;
        RECT 586.140 20.440 586.400 20.700 ;
      LAYER met2 ;
        RECT 694.740 220.000 695.020 224.000 ;
        RECT 694.760 212.490 694.900 220.000 ;
        RECT 694.700 212.170 694.960 212.490 ;
        RECT 586.140 210.130 586.400 210.450 ;
        RECT 586.200 20.730 586.340 210.130 ;
        RECT 579.700 20.410 579.960 20.730 ;
        RECT 586.140 20.410 586.400 20.730 ;
        RECT 579.760 2.400 579.900 20.410 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 284.350 159.020 284.670 159.080 ;
        RECT 287.110 159.020 287.430 159.080 ;
        RECT 284.350 158.880 287.430 159.020 ;
        RECT 284.350 158.820 284.670 158.880 ;
        RECT 287.110 158.820 287.430 158.880 ;
        RECT 86.090 24.720 86.410 24.780 ;
        RECT 283.430 24.720 283.750 24.780 ;
        RECT 86.090 24.580 283.750 24.720 ;
        RECT 86.090 24.520 86.410 24.580 ;
        RECT 283.430 24.520 283.750 24.580 ;
      LAYER via ;
        RECT 284.380 158.820 284.640 159.080 ;
        RECT 287.140 158.820 287.400 159.080 ;
        RECT 86.120 24.520 86.380 24.780 ;
        RECT 283.460 24.520 283.720 24.780 ;
      LAYER met2 ;
        RECT 288.560 220.730 288.840 224.000 ;
        RECT 287.200 220.590 288.840 220.730 ;
        RECT 287.200 159.110 287.340 220.590 ;
        RECT 288.560 220.000 288.840 220.590 ;
        RECT 284.380 158.790 284.640 159.110 ;
        RECT 287.140 158.790 287.400 159.110 ;
        RECT 284.440 62.290 284.580 158.790 ;
        RECT 283.520 62.150 284.580 62.290 ;
        RECT 283.520 24.810 283.660 62.150 ;
        RECT 86.120 24.490 86.380 24.810 ;
        RECT 283.460 24.490 283.720 24.810 ;
        RECT 86.180 2.400 86.320 24.490 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 599.910 212.060 600.230 212.120 ;
        RECT 709.390 212.060 709.710 212.120 ;
        RECT 599.910 211.920 709.710 212.060 ;
        RECT 599.910 211.860 600.230 211.920 ;
        RECT 709.390 211.860 709.710 211.920 ;
        RECT 597.150 20.640 597.470 20.700 ;
        RECT 599.910 20.640 600.230 20.700 ;
        RECT 597.150 20.500 600.230 20.640 ;
        RECT 597.150 20.440 597.470 20.500 ;
        RECT 599.910 20.440 600.230 20.500 ;
      LAYER via ;
        RECT 599.940 211.860 600.200 212.120 ;
        RECT 709.420 211.860 709.680 212.120 ;
        RECT 597.180 20.440 597.440 20.700 ;
        RECT 599.940 20.440 600.200 20.700 ;
      LAYER met2 ;
        RECT 709.460 220.000 709.740 224.000 ;
        RECT 709.480 212.150 709.620 220.000 ;
        RECT 599.940 211.830 600.200 212.150 ;
        RECT 709.420 211.830 709.680 212.150 ;
        RECT 600.000 20.730 600.140 211.830 ;
        RECT 597.180 20.410 597.440 20.730 ;
        RECT 599.940 20.410 600.200 20.730 ;
        RECT 597.240 2.400 597.380 20.410 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 620.610 209.000 620.930 209.060 ;
        RECT 724.110 209.000 724.430 209.060 ;
        RECT 620.610 208.860 724.430 209.000 ;
        RECT 620.610 208.800 620.930 208.860 ;
        RECT 724.110 208.800 724.430 208.860 ;
        RECT 615.090 18.260 615.410 18.320 ;
        RECT 620.610 18.260 620.930 18.320 ;
        RECT 615.090 18.120 620.930 18.260 ;
        RECT 615.090 18.060 615.410 18.120 ;
        RECT 620.610 18.060 620.930 18.120 ;
      LAYER via ;
        RECT 620.640 208.800 620.900 209.060 ;
        RECT 724.140 208.800 724.400 209.060 ;
        RECT 615.120 18.060 615.380 18.320 ;
        RECT 620.640 18.060 620.900 18.320 ;
      LAYER met2 ;
        RECT 724.180 220.000 724.460 224.000 ;
        RECT 724.200 209.090 724.340 220.000 ;
        RECT 620.640 208.770 620.900 209.090 ;
        RECT 724.140 208.770 724.400 209.090 ;
        RECT 620.700 18.350 620.840 208.770 ;
        RECT 615.120 18.030 615.380 18.350 ;
        RECT 620.640 18.030 620.900 18.350 ;
        RECT 615.180 2.400 615.320 18.030 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 110.010 25.060 110.330 25.120 ;
        RECT 303.670 25.060 303.990 25.120 ;
        RECT 110.010 24.920 303.990 25.060 ;
        RECT 110.010 24.860 110.330 24.920 ;
        RECT 303.670 24.860 303.990 24.920 ;
      LAYER via ;
        RECT 110.040 24.860 110.300 25.120 ;
        RECT 303.700 24.860 303.960 25.120 ;
      LAYER met2 ;
        RECT 307.880 220.730 308.160 224.000 ;
        RECT 303.760 220.590 308.160 220.730 ;
        RECT 303.760 25.150 303.900 220.590 ;
        RECT 307.880 220.000 308.160 220.590 ;
        RECT 110.040 24.830 110.300 25.150 ;
        RECT 303.700 24.830 303.960 25.150 ;
        RECT 110.100 12.650 110.240 24.830 ;
        RECT 109.640 12.510 110.240 12.650 ;
        RECT 109.640 2.400 109.780 12.510 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 133.470 25.400 133.790 25.460 ;
        RECT 324.370 25.400 324.690 25.460 ;
        RECT 133.470 25.260 324.690 25.400 ;
        RECT 133.470 25.200 133.790 25.260 ;
        RECT 324.370 25.200 324.690 25.260 ;
      LAYER via ;
        RECT 133.500 25.200 133.760 25.460 ;
        RECT 324.400 25.200 324.660 25.460 ;
      LAYER met2 ;
        RECT 327.660 220.730 327.940 224.000 ;
        RECT 324.460 220.590 327.940 220.730 ;
        RECT 324.460 25.490 324.600 220.590 ;
        RECT 327.660 220.000 327.940 220.590 ;
        RECT 133.500 25.170 133.760 25.490 ;
        RECT 324.400 25.170 324.660 25.490 ;
        RECT 133.560 2.400 133.700 25.170 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 25.740 151.730 25.800 ;
        RECT 338.170 25.740 338.490 25.800 ;
        RECT 151.410 25.600 338.490 25.740 ;
        RECT 151.410 25.540 151.730 25.600 ;
        RECT 338.170 25.540 338.490 25.600 ;
      LAYER via ;
        RECT 151.440 25.540 151.700 25.800 ;
        RECT 338.200 25.540 338.460 25.800 ;
      LAYER met2 ;
        RECT 342.380 220.730 342.660 224.000 ;
        RECT 338.260 220.590 342.660 220.730 ;
        RECT 338.260 25.830 338.400 220.590 ;
        RECT 342.380 220.000 342.660 220.590 ;
        RECT 151.440 25.510 151.700 25.830 ;
        RECT 338.200 25.510 338.460 25.830 ;
        RECT 151.500 2.400 151.640 25.510 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 169.350 26.080 169.670 26.140 ;
        RECT 352.430 26.080 352.750 26.140 ;
        RECT 169.350 25.940 352.750 26.080 ;
        RECT 169.350 25.880 169.670 25.940 ;
        RECT 352.430 25.880 352.750 25.940 ;
      LAYER via ;
        RECT 169.380 25.880 169.640 26.140 ;
        RECT 352.460 25.880 352.720 26.140 ;
      LAYER met2 ;
        RECT 357.100 220.730 357.380 224.000 ;
        RECT 352.520 220.590 357.380 220.730 ;
        RECT 352.520 26.170 352.660 220.590 ;
        RECT 357.100 220.000 357.380 220.590 ;
        RECT 169.380 25.850 169.640 26.170 ;
        RECT 352.460 25.850 352.720 26.170 ;
        RECT 169.440 2.400 169.580 25.850 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 367.685 144.925 367.855 193.035 ;
      LAYER mcon ;
        RECT 367.685 192.865 367.855 193.035 ;
      LAYER met1 ;
        RECT 367.610 193.020 367.930 193.080 ;
        RECT 367.415 192.880 367.930 193.020 ;
        RECT 367.610 192.820 367.930 192.880 ;
        RECT 367.625 145.080 367.915 145.125 ;
        RECT 368.070 145.080 368.390 145.140 ;
        RECT 367.625 144.940 368.390 145.080 ;
        RECT 367.625 144.895 367.915 144.940 ;
        RECT 368.070 144.880 368.390 144.940 ;
        RECT 186.830 26.420 187.150 26.480 ;
        RECT 366.230 26.420 366.550 26.480 ;
        RECT 186.830 26.280 366.550 26.420 ;
        RECT 186.830 26.220 187.150 26.280 ;
        RECT 366.230 26.220 366.550 26.280 ;
      LAYER via ;
        RECT 367.640 192.820 367.900 193.080 ;
        RECT 368.100 144.880 368.360 145.140 ;
        RECT 186.860 26.220 187.120 26.480 ;
        RECT 366.260 26.220 366.520 26.480 ;
      LAYER met2 ;
        RECT 371.820 220.000 372.100 224.000 ;
        RECT 371.840 194.325 371.980 220.000 ;
        RECT 371.770 193.955 372.050 194.325 ;
        RECT 367.170 193.530 367.450 193.645 ;
        RECT 367.170 193.390 367.840 193.530 ;
        RECT 367.170 193.275 367.450 193.390 ;
        RECT 367.700 193.110 367.840 193.390 ;
        RECT 367.640 192.790 367.900 193.110 ;
        RECT 368.100 144.850 368.360 145.170 ;
        RECT 368.160 110.570 368.300 144.850 ;
        RECT 367.240 110.430 368.300 110.570 ;
        RECT 367.240 62.290 367.380 110.430 ;
        RECT 366.320 62.150 367.380 62.290 ;
        RECT 366.320 26.510 366.460 62.150 ;
        RECT 186.860 26.190 187.120 26.510 ;
        RECT 366.260 26.190 366.520 26.510 ;
        RECT 186.920 2.400 187.060 26.190 ;
        RECT 186.710 -4.800 187.270 2.400 ;
      LAYER via2 ;
        RECT 371.770 194.000 372.050 194.280 ;
        RECT 367.170 193.320 367.450 193.600 ;
      LAYER met3 ;
        RECT 371.745 194.290 372.075 194.305 ;
        RECT 366.470 193.990 372.075 194.290 ;
        RECT 366.470 193.610 366.770 193.990 ;
        RECT 371.745 193.975 372.075 193.990 ;
        RECT 367.145 193.610 367.475 193.625 ;
        RECT 366.470 193.310 367.475 193.610 ;
        RECT 367.145 193.295 367.475 193.310 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 341.005 207.825 341.175 210.035 ;
        RECT 376.885 209.185 377.055 210.035 ;
      LAYER mcon ;
        RECT 341.005 209.865 341.175 210.035 ;
        RECT 376.885 209.865 377.055 210.035 ;
      LAYER met1 ;
        RECT 340.945 210.020 341.235 210.065 ;
        RECT 376.825 210.020 377.115 210.065 ;
        RECT 340.945 209.880 377.115 210.020 ;
        RECT 340.945 209.835 341.235 209.880 ;
        RECT 376.825 209.835 377.115 209.880 ;
        RECT 376.825 209.340 377.115 209.385 ;
        RECT 386.010 209.340 386.330 209.400 ;
        RECT 376.825 209.200 386.330 209.340 ;
        RECT 376.825 209.155 377.115 209.200 ;
        RECT 386.010 209.140 386.330 209.200 ;
        RECT 206.610 207.980 206.930 208.040 ;
        RECT 340.945 207.980 341.235 208.025 ;
        RECT 206.610 207.840 341.235 207.980 ;
        RECT 206.610 207.780 206.930 207.840 ;
        RECT 340.945 207.795 341.235 207.840 ;
        RECT 204.770 2.960 205.090 3.020 ;
        RECT 206.610 2.960 206.930 3.020 ;
        RECT 204.770 2.820 206.930 2.960 ;
        RECT 204.770 2.760 205.090 2.820 ;
        RECT 206.610 2.760 206.930 2.820 ;
      LAYER via ;
        RECT 386.040 209.140 386.300 209.400 ;
        RECT 206.640 207.780 206.900 208.040 ;
        RECT 204.800 2.760 205.060 3.020 ;
        RECT 206.640 2.760 206.900 3.020 ;
      LAYER met2 ;
        RECT 386.080 220.000 386.360 224.000 ;
        RECT 386.100 209.430 386.240 220.000 ;
        RECT 386.040 209.110 386.300 209.430 ;
        RECT 206.640 207.750 206.900 208.070 ;
        RECT 206.700 3.050 206.840 207.750 ;
        RECT 204.800 2.730 205.060 3.050 ;
        RECT 206.640 2.730 206.900 3.050 ;
        RECT 204.860 2.400 205.000 2.730 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 227.310 208.320 227.630 208.380 ;
        RECT 400.730 208.320 401.050 208.380 ;
        RECT 227.310 208.180 401.050 208.320 ;
        RECT 227.310 208.120 227.630 208.180 ;
        RECT 400.730 208.120 401.050 208.180 ;
        RECT 222.710 17.580 223.030 17.640 ;
        RECT 227.310 17.580 227.630 17.640 ;
        RECT 222.710 17.440 227.630 17.580 ;
        RECT 222.710 17.380 223.030 17.440 ;
        RECT 227.310 17.380 227.630 17.440 ;
      LAYER via ;
        RECT 227.340 208.120 227.600 208.380 ;
        RECT 400.760 208.120 401.020 208.380 ;
        RECT 222.740 17.380 223.000 17.640 ;
        RECT 227.340 17.380 227.600 17.640 ;
      LAYER met2 ;
        RECT 400.800 220.000 401.080 224.000 ;
        RECT 400.820 208.410 400.960 220.000 ;
        RECT 227.340 208.090 227.600 208.410 ;
        RECT 400.760 208.090 401.020 208.410 ;
        RECT 227.400 17.670 227.540 208.090 ;
        RECT 222.740 17.350 223.000 17.670 ;
        RECT 227.340 17.350 227.600 17.670 ;
        RECT 222.800 2.400 222.940 17.350 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 210.700 20.630 210.760 ;
        RECT 234.210 210.700 234.530 210.760 ;
        RECT 20.310 210.560 234.530 210.700 ;
        RECT 20.310 210.500 20.630 210.560 ;
        RECT 234.210 210.500 234.530 210.560 ;
      LAYER via ;
        RECT 20.340 210.500 20.600 210.760 ;
        RECT 234.240 210.500 234.500 210.760 ;
      LAYER met2 ;
        RECT 234.280 220.000 234.560 224.000 ;
        RECT 234.300 210.790 234.440 220.000 ;
        RECT 20.340 210.470 20.600 210.790 ;
        RECT 234.240 210.470 234.500 210.790 ;
        RECT 20.400 2.400 20.540 210.470 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.910 212.400 48.230 212.460 ;
        RECT 253.990 212.400 254.310 212.460 ;
        RECT 47.910 212.260 254.310 212.400 ;
        RECT 47.910 212.200 48.230 212.260 ;
        RECT 253.990 212.200 254.310 212.260 ;
        RECT 44.230 16.900 44.550 16.960 ;
        RECT 47.910 16.900 48.230 16.960 ;
        RECT 44.230 16.760 48.230 16.900 ;
        RECT 44.230 16.700 44.550 16.760 ;
        RECT 47.910 16.700 48.230 16.760 ;
      LAYER via ;
        RECT 47.940 212.200 48.200 212.460 ;
        RECT 254.020 212.200 254.280 212.460 ;
        RECT 44.260 16.700 44.520 16.960 ;
        RECT 47.940 16.700 48.200 16.960 ;
      LAYER met2 ;
        RECT 254.060 220.000 254.340 224.000 ;
        RECT 254.080 212.490 254.220 220.000 ;
        RECT 47.940 212.170 48.200 212.490 ;
        RECT 254.020 212.170 254.280 212.490 ;
        RECT 48.000 16.990 48.140 212.170 ;
        RECT 44.260 16.670 44.520 16.990 ;
        RECT 47.940 16.670 48.200 16.990 ;
        RECT 44.320 2.400 44.460 16.670 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 323.065 207.485 323.235 209.695 ;
        RECT 401.265 207.485 401.435 208.335 ;
      LAYER mcon ;
        RECT 323.065 209.525 323.235 209.695 ;
        RECT 401.265 208.165 401.435 208.335 ;
      LAYER met1 ;
        RECT 248.010 210.360 248.330 210.420 ;
        RECT 299.530 210.360 299.850 210.420 ;
        RECT 248.010 210.220 299.850 210.360 ;
        RECT 248.010 210.160 248.330 210.220 ;
        RECT 299.530 210.160 299.850 210.220 ;
        RECT 299.530 209.680 299.850 209.740 ;
        RECT 323.005 209.680 323.295 209.725 ;
        RECT 299.530 209.540 323.295 209.680 ;
        RECT 299.530 209.480 299.850 209.540 ;
        RECT 323.005 209.495 323.295 209.540 ;
        RECT 401.205 208.320 401.495 208.365 ;
        RECT 416.830 208.320 417.150 208.380 ;
        RECT 401.205 208.180 417.150 208.320 ;
        RECT 401.205 208.135 401.495 208.180 ;
        RECT 416.830 208.120 417.150 208.180 ;
        RECT 323.005 207.640 323.295 207.685 ;
        RECT 401.205 207.640 401.495 207.685 ;
        RECT 323.005 207.500 401.495 207.640 ;
        RECT 323.005 207.455 323.295 207.500 ;
        RECT 401.205 207.455 401.495 207.500 ;
      LAYER via ;
        RECT 248.040 210.160 248.300 210.420 ;
        RECT 299.560 210.160 299.820 210.420 ;
        RECT 299.560 209.480 299.820 209.740 ;
        RECT 416.860 208.120 417.120 208.380 ;
      LAYER met2 ;
        RECT 420.580 220.730 420.860 224.000 ;
        RECT 416.920 220.590 420.860 220.730 ;
        RECT 248.040 210.130 248.300 210.450 ;
        RECT 299.560 210.130 299.820 210.450 ;
        RECT 248.100 3.130 248.240 210.130 ;
        RECT 299.620 209.770 299.760 210.130 ;
        RECT 299.560 209.450 299.820 209.770 ;
        RECT 416.920 208.410 417.060 220.590 ;
        RECT 420.580 220.000 420.860 220.590 ;
        RECT 416.860 208.090 417.120 208.410 ;
        RECT 246.720 2.990 248.240 3.130 ;
        RECT 246.720 2.400 246.860 2.990 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 268.710 211.040 269.030 211.100 ;
        RECT 435.230 211.040 435.550 211.100 ;
        RECT 268.710 210.900 435.550 211.040 ;
        RECT 268.710 210.840 269.030 210.900 ;
        RECT 435.230 210.840 435.550 210.900 ;
        RECT 264.110 17.240 264.430 17.300 ;
        RECT 268.710 17.240 269.030 17.300 ;
        RECT 264.110 17.100 269.030 17.240 ;
        RECT 264.110 17.040 264.430 17.100 ;
        RECT 268.710 17.040 269.030 17.100 ;
      LAYER via ;
        RECT 268.740 210.840 269.000 211.100 ;
        RECT 435.260 210.840 435.520 211.100 ;
        RECT 264.140 17.040 264.400 17.300 ;
        RECT 268.740 17.040 269.000 17.300 ;
      LAYER met2 ;
        RECT 435.300 220.000 435.580 224.000 ;
        RECT 435.320 211.130 435.460 220.000 ;
        RECT 268.740 210.810 269.000 211.130 ;
        RECT 435.260 210.810 435.520 211.130 ;
        RECT 268.800 17.330 268.940 210.810 ;
        RECT 264.140 17.010 264.400 17.330 ;
        RECT 268.740 17.010 269.000 17.330 ;
        RECT 264.200 2.400 264.340 17.010 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 282.125 2.805 282.295 18.275 ;
      LAYER mcon ;
        RECT 282.125 18.105 282.295 18.275 ;
      LAYER met1 ;
        RECT 282.510 211.380 282.830 211.440 ;
        RECT 449.950 211.380 450.270 211.440 ;
        RECT 282.510 211.240 450.270 211.380 ;
        RECT 282.510 211.180 282.830 211.240 ;
        RECT 449.950 211.180 450.270 211.240 ;
        RECT 282.065 18.260 282.355 18.305 ;
        RECT 282.510 18.260 282.830 18.320 ;
        RECT 282.065 18.120 282.830 18.260 ;
        RECT 282.065 18.075 282.355 18.120 ;
        RECT 282.510 18.060 282.830 18.120 ;
        RECT 282.050 2.960 282.370 3.020 ;
        RECT 281.855 2.820 282.370 2.960 ;
        RECT 282.050 2.760 282.370 2.820 ;
      LAYER via ;
        RECT 282.540 211.180 282.800 211.440 ;
        RECT 449.980 211.180 450.240 211.440 ;
        RECT 282.540 18.060 282.800 18.320 ;
        RECT 282.080 2.760 282.340 3.020 ;
      LAYER met2 ;
        RECT 450.020 220.000 450.300 224.000 ;
        RECT 450.040 211.470 450.180 220.000 ;
        RECT 282.540 211.150 282.800 211.470 ;
        RECT 449.980 211.150 450.240 211.470 ;
        RECT 282.600 18.350 282.740 211.150 ;
        RECT 282.540 18.030 282.800 18.350 ;
        RECT 282.080 2.730 282.340 3.050 ;
        RECT 282.140 2.400 282.280 2.730 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 303.210 213.080 303.530 213.140 ;
        RECT 303.210 212.940 331.500 213.080 ;
        RECT 303.210 212.880 303.530 212.940 ;
        RECT 331.360 212.740 331.500 212.940 ;
        RECT 464.670 212.740 464.990 212.800 ;
        RECT 331.360 212.600 464.990 212.740 ;
        RECT 464.670 212.540 464.990 212.600 ;
        RECT 299.990 20.640 300.310 20.700 ;
        RECT 303.210 20.640 303.530 20.700 ;
        RECT 299.990 20.500 303.530 20.640 ;
        RECT 299.990 20.440 300.310 20.500 ;
        RECT 303.210 20.440 303.530 20.500 ;
      LAYER via ;
        RECT 303.240 212.880 303.500 213.140 ;
        RECT 464.700 212.540 464.960 212.800 ;
        RECT 300.020 20.440 300.280 20.700 ;
        RECT 303.240 20.440 303.500 20.700 ;
      LAYER met2 ;
        RECT 464.740 220.000 465.020 224.000 ;
        RECT 303.240 212.850 303.500 213.170 ;
        RECT 303.300 20.730 303.440 212.850 ;
        RECT 464.760 212.830 464.900 220.000 ;
        RECT 464.700 212.510 464.960 212.830 ;
        RECT 300.020 20.410 300.280 20.730 ;
        RECT 303.240 20.410 303.500 20.730 ;
        RECT 300.080 2.400 300.220 20.410 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 323.910 213.420 324.230 213.480 ;
        RECT 479.390 213.420 479.710 213.480 ;
        RECT 323.910 213.280 367.840 213.420 ;
        RECT 323.910 213.220 324.230 213.280 ;
        RECT 367.700 213.080 367.840 213.280 ;
        RECT 371.840 213.280 479.710 213.420 ;
        RECT 371.840 213.080 371.980 213.280 ;
        RECT 479.390 213.220 479.710 213.280 ;
        RECT 367.700 212.940 371.980 213.080 ;
        RECT 317.930 17.240 318.250 17.300 ;
        RECT 323.910 17.240 324.230 17.300 ;
        RECT 317.930 17.100 324.230 17.240 ;
        RECT 317.930 17.040 318.250 17.100 ;
        RECT 323.910 17.040 324.230 17.100 ;
      LAYER via ;
        RECT 323.940 213.220 324.200 213.480 ;
        RECT 479.420 213.220 479.680 213.480 ;
        RECT 317.960 17.040 318.220 17.300 ;
        RECT 323.940 17.040 324.200 17.300 ;
      LAYER met2 ;
        RECT 479.460 220.000 479.740 224.000 ;
        RECT 479.480 213.510 479.620 220.000 ;
        RECT 323.940 213.190 324.200 213.510 ;
        RECT 479.420 213.190 479.680 213.510 ;
        RECT 324.000 17.330 324.140 213.190 ;
        RECT 317.960 17.010 318.220 17.330 ;
        RECT 323.940 17.010 324.200 17.330 ;
        RECT 318.020 2.400 318.160 17.010 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 347.905 207.145 348.075 209.015 ;
        RECT 371.825 208.845 371.995 213.775 ;
      LAYER mcon ;
        RECT 371.825 213.605 371.995 213.775 ;
        RECT 347.905 208.845 348.075 209.015 ;
      LAYER met1 ;
        RECT 371.765 213.760 372.055 213.805 ;
        RECT 494.110 213.760 494.430 213.820 ;
        RECT 371.765 213.620 494.430 213.760 ;
        RECT 371.765 213.575 372.055 213.620 ;
        RECT 494.110 213.560 494.430 213.620 ;
        RECT 347.845 209.000 348.135 209.045 ;
        RECT 371.765 209.000 372.055 209.045 ;
        RECT 347.845 208.860 372.055 209.000 ;
        RECT 347.845 208.815 348.135 208.860 ;
        RECT 371.765 208.815 372.055 208.860 ;
        RECT 337.710 207.300 338.030 207.360 ;
        RECT 347.845 207.300 348.135 207.345 ;
        RECT 337.710 207.160 348.135 207.300 ;
        RECT 337.710 207.100 338.030 207.160 ;
        RECT 347.845 207.115 348.135 207.160 ;
      LAYER via ;
        RECT 494.140 213.560 494.400 213.820 ;
        RECT 337.740 207.100 338.000 207.360 ;
      LAYER met2 ;
        RECT 494.180 220.000 494.460 224.000 ;
        RECT 494.200 213.850 494.340 220.000 ;
        RECT 494.140 213.530 494.400 213.850 ;
        RECT 337.740 207.070 338.000 207.390 ;
        RECT 337.800 3.130 337.940 207.070 ;
        RECT 335.960 2.990 337.940 3.130 ;
        RECT 335.960 2.400 336.100 2.990 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 358.410 207.300 358.730 207.360 ;
        RECT 508.830 207.300 509.150 207.360 ;
        RECT 358.410 207.160 509.150 207.300 ;
        RECT 358.410 207.100 358.730 207.160 ;
        RECT 508.830 207.100 509.150 207.160 ;
        RECT 353.350 16.220 353.670 16.280 ;
        RECT 358.410 16.220 358.730 16.280 ;
        RECT 353.350 16.080 358.730 16.220 ;
        RECT 353.350 16.020 353.670 16.080 ;
        RECT 358.410 16.020 358.730 16.080 ;
      LAYER via ;
        RECT 358.440 207.100 358.700 207.360 ;
        RECT 508.860 207.100 509.120 207.360 ;
        RECT 353.380 16.020 353.640 16.280 ;
        RECT 358.440 16.020 358.700 16.280 ;
      LAYER met2 ;
        RECT 508.900 220.000 509.180 224.000 ;
        RECT 508.920 207.390 509.060 220.000 ;
        RECT 358.440 207.070 358.700 207.390 ;
        RECT 508.860 207.070 509.120 207.390 ;
        RECT 358.500 16.310 358.640 207.070 ;
        RECT 353.380 15.990 353.640 16.310 ;
        RECT 358.440 15.990 358.700 16.310 ;
        RECT 353.440 2.400 353.580 15.990 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 209.000 372.530 209.060 ;
        RECT 523.550 209.000 523.870 209.060 ;
        RECT 372.210 208.860 523.870 209.000 ;
        RECT 372.210 208.800 372.530 208.860 ;
        RECT 523.550 208.800 523.870 208.860 ;
        RECT 371.290 2.960 371.610 3.020 ;
        RECT 372.210 2.960 372.530 3.020 ;
        RECT 371.290 2.820 372.530 2.960 ;
        RECT 371.290 2.760 371.610 2.820 ;
        RECT 372.210 2.760 372.530 2.820 ;
      LAYER via ;
        RECT 372.240 208.800 372.500 209.060 ;
        RECT 523.580 208.800 523.840 209.060 ;
        RECT 371.320 2.760 371.580 3.020 ;
        RECT 372.240 2.760 372.500 3.020 ;
      LAYER met2 ;
        RECT 523.620 220.000 523.900 224.000 ;
        RECT 523.640 209.090 523.780 220.000 ;
        RECT 372.240 208.770 372.500 209.090 ;
        RECT 523.580 208.770 523.840 209.090 ;
        RECT 372.300 3.050 372.440 208.770 ;
        RECT 371.320 2.730 371.580 3.050 ;
        RECT 372.240 2.730 372.500 3.050 ;
        RECT 371.380 2.400 371.520 2.730 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 392.910 209.340 393.230 209.400 ;
        RECT 538.270 209.340 538.590 209.400 ;
        RECT 392.910 209.200 538.590 209.340 ;
        RECT 392.910 209.140 393.230 209.200 ;
        RECT 538.270 209.140 538.590 209.200 ;
        RECT 389.230 15.880 389.550 15.940 ;
        RECT 392.910 15.880 393.230 15.940 ;
        RECT 389.230 15.740 393.230 15.880 ;
        RECT 389.230 15.680 389.550 15.740 ;
        RECT 392.910 15.680 393.230 15.740 ;
      LAYER via ;
        RECT 392.940 209.140 393.200 209.400 ;
        RECT 538.300 209.140 538.560 209.400 ;
        RECT 389.260 15.680 389.520 15.940 ;
        RECT 392.940 15.680 393.200 15.940 ;
      LAYER met2 ;
        RECT 538.340 220.000 538.620 224.000 ;
        RECT 538.360 209.430 538.500 220.000 ;
        RECT 392.940 209.110 393.200 209.430 ;
        RECT 538.300 209.110 538.560 209.430 ;
        RECT 393.000 15.970 393.140 209.110 ;
        RECT 389.260 15.650 389.520 15.970 ;
        RECT 392.940 15.650 393.200 15.970 ;
        RECT 389.320 2.400 389.460 15.650 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 413.610 210.700 413.930 210.760 ;
        RECT 552.530 210.700 552.850 210.760 ;
        RECT 413.610 210.560 552.850 210.700 ;
        RECT 413.610 210.500 413.930 210.560 ;
        RECT 552.530 210.500 552.850 210.560 ;
        RECT 407.170 17.240 407.490 17.300 ;
        RECT 413.610 17.240 413.930 17.300 ;
        RECT 407.170 17.100 413.930 17.240 ;
        RECT 407.170 17.040 407.490 17.100 ;
        RECT 413.610 17.040 413.930 17.100 ;
      LAYER via ;
        RECT 413.640 210.500 413.900 210.760 ;
        RECT 552.560 210.500 552.820 210.760 ;
        RECT 407.200 17.040 407.460 17.300 ;
        RECT 413.640 17.040 413.900 17.300 ;
      LAYER met2 ;
        RECT 552.600 220.000 552.880 224.000 ;
        RECT 552.620 210.790 552.760 220.000 ;
        RECT 413.640 210.470 413.900 210.790 ;
        RECT 552.560 210.470 552.820 210.790 ;
        RECT 413.700 17.330 413.840 210.470 ;
        RECT 407.200 17.010 407.460 17.330 ;
        RECT 413.640 17.010 413.900 17.330 ;
        RECT 407.260 2.400 407.400 17.010 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.150 212.060 68.470 212.120 ;
        RECT 273.770 212.060 274.090 212.120 ;
        RECT 68.150 211.920 274.090 212.060 ;
        RECT 68.150 211.860 68.470 211.920 ;
        RECT 273.770 211.860 274.090 211.920 ;
      LAYER via ;
        RECT 68.180 211.860 68.440 212.120 ;
        RECT 273.800 211.860 274.060 212.120 ;
      LAYER met2 ;
        RECT 273.840 220.000 274.120 224.000 ;
        RECT 273.860 212.150 274.000 220.000 ;
        RECT 68.180 211.830 68.440 212.150 ;
        RECT 273.800 211.830 274.060 212.150 ;
        RECT 68.240 2.400 68.380 211.830 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 210.360 427.730 210.420 ;
        RECT 567.250 210.360 567.570 210.420 ;
        RECT 427.410 210.220 567.570 210.360 ;
        RECT 427.410 210.160 427.730 210.220 ;
        RECT 567.250 210.160 567.570 210.220 ;
        RECT 424.650 20.640 424.970 20.700 ;
        RECT 427.410 20.640 427.730 20.700 ;
        RECT 424.650 20.500 427.730 20.640 ;
        RECT 424.650 20.440 424.970 20.500 ;
        RECT 427.410 20.440 427.730 20.500 ;
      LAYER via ;
        RECT 427.440 210.160 427.700 210.420 ;
        RECT 567.280 210.160 567.540 210.420 ;
        RECT 424.680 20.440 424.940 20.700 ;
        RECT 427.440 20.440 427.700 20.700 ;
      LAYER met2 ;
        RECT 567.320 220.000 567.600 224.000 ;
        RECT 567.340 210.450 567.480 220.000 ;
        RECT 427.440 210.130 427.700 210.450 ;
        RECT 567.280 210.130 567.540 210.450 ;
        RECT 427.500 20.730 427.640 210.130 ;
        RECT 424.680 20.410 424.940 20.730 ;
        RECT 427.440 20.410 427.700 20.730 ;
        RECT 424.740 2.400 424.880 20.410 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 448.110 212.060 448.430 212.120 ;
        RECT 581.970 212.060 582.290 212.120 ;
        RECT 448.110 211.920 582.290 212.060 ;
        RECT 448.110 211.860 448.430 211.920 ;
        RECT 581.970 211.860 582.290 211.920 ;
        RECT 442.590 15.880 442.910 15.940 ;
        RECT 448.110 15.880 448.430 15.940 ;
        RECT 442.590 15.740 448.430 15.880 ;
        RECT 442.590 15.680 442.910 15.740 ;
        RECT 448.110 15.680 448.430 15.740 ;
      LAYER via ;
        RECT 448.140 211.860 448.400 212.120 ;
        RECT 582.000 211.860 582.260 212.120 ;
        RECT 442.620 15.680 442.880 15.940 ;
        RECT 448.140 15.680 448.400 15.940 ;
      LAYER met2 ;
        RECT 582.040 220.000 582.320 224.000 ;
        RECT 582.060 212.150 582.200 220.000 ;
        RECT 448.140 211.830 448.400 212.150 ;
        RECT 582.000 211.830 582.260 212.150 ;
        RECT 448.200 15.970 448.340 211.830 ;
        RECT 442.620 15.650 442.880 15.970 ;
        RECT 448.140 15.650 448.400 15.970 ;
        RECT 442.680 2.400 442.820 15.650 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.910 212.400 462.230 212.460 ;
        RECT 596.690 212.400 597.010 212.460 ;
        RECT 461.910 212.260 597.010 212.400 ;
        RECT 461.910 212.200 462.230 212.260 ;
        RECT 596.690 212.200 597.010 212.260 ;
        RECT 460.530 14.180 460.850 14.240 ;
        RECT 461.910 14.180 462.230 14.240 ;
        RECT 460.530 14.040 462.230 14.180 ;
        RECT 460.530 13.980 460.850 14.040 ;
        RECT 461.910 13.980 462.230 14.040 ;
      LAYER via ;
        RECT 461.940 212.200 462.200 212.460 ;
        RECT 596.720 212.200 596.980 212.460 ;
        RECT 460.560 13.980 460.820 14.240 ;
        RECT 461.940 13.980 462.200 14.240 ;
      LAYER met2 ;
        RECT 596.760 220.000 597.040 224.000 ;
        RECT 596.780 212.490 596.920 220.000 ;
        RECT 461.940 212.170 462.200 212.490 ;
        RECT 596.720 212.170 596.980 212.490 ;
        RECT 462.000 14.270 462.140 212.170 ;
        RECT 460.560 13.950 460.820 14.270 ;
        RECT 461.940 13.950 462.200 14.270 ;
        RECT 460.620 2.400 460.760 13.950 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 212.740 482.930 212.800 ;
        RECT 611.410 212.740 611.730 212.800 ;
        RECT 482.610 212.600 611.730 212.740 ;
        RECT 482.610 212.540 482.930 212.600 ;
        RECT 611.410 212.540 611.730 212.600 ;
        RECT 478.470 16.220 478.790 16.280 ;
        RECT 482.610 16.220 482.930 16.280 ;
        RECT 478.470 16.080 482.930 16.220 ;
        RECT 478.470 16.020 478.790 16.080 ;
        RECT 482.610 16.020 482.930 16.080 ;
      LAYER via ;
        RECT 482.640 212.540 482.900 212.800 ;
        RECT 611.440 212.540 611.700 212.800 ;
        RECT 478.500 16.020 478.760 16.280 ;
        RECT 482.640 16.020 482.900 16.280 ;
      LAYER met2 ;
        RECT 611.480 220.000 611.760 224.000 ;
        RECT 611.500 212.830 611.640 220.000 ;
        RECT 482.640 212.510 482.900 212.830 ;
        RECT 611.440 212.510 611.700 212.830 ;
        RECT 482.700 16.310 482.840 212.510 ;
        RECT 478.500 15.990 478.760 16.310 ;
        RECT 482.640 15.990 482.900 16.310 ;
        RECT 478.560 2.400 478.700 15.990 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 496.410 213.420 496.730 213.480 ;
        RECT 626.130 213.420 626.450 213.480 ;
        RECT 496.410 213.280 626.450 213.420 ;
        RECT 496.410 213.220 496.730 213.280 ;
        RECT 626.130 213.220 626.450 213.280 ;
      LAYER via ;
        RECT 496.440 213.220 496.700 213.480 ;
        RECT 626.160 213.220 626.420 213.480 ;
      LAYER met2 ;
        RECT 626.200 220.000 626.480 224.000 ;
        RECT 626.220 213.510 626.360 220.000 ;
        RECT 496.440 213.190 496.700 213.510 ;
        RECT 626.160 213.190 626.420 213.510 ;
        RECT 496.500 2.400 496.640 213.190 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 619.765 207.825 619.935 209.355 ;
      LAYER mcon ;
        RECT 619.765 209.185 619.935 209.355 ;
      LAYER met1 ;
        RECT 619.705 209.340 619.995 209.385 ;
        RECT 637.630 209.340 637.950 209.400 ;
        RECT 619.705 209.200 637.950 209.340 ;
        RECT 619.705 209.155 619.995 209.200 ;
        RECT 637.630 209.140 637.950 209.200 ;
        RECT 517.110 207.980 517.430 208.040 ;
        RECT 619.705 207.980 619.995 208.025 ;
        RECT 517.110 207.840 619.995 207.980 ;
        RECT 517.110 207.780 517.430 207.840 ;
        RECT 619.705 207.795 619.995 207.840 ;
        RECT 513.890 20.640 514.210 20.700 ;
        RECT 517.110 20.640 517.430 20.700 ;
        RECT 513.890 20.500 517.430 20.640 ;
        RECT 513.890 20.440 514.210 20.500 ;
        RECT 517.110 20.440 517.430 20.500 ;
      LAYER via ;
        RECT 637.660 209.140 637.920 209.400 ;
        RECT 517.140 207.780 517.400 208.040 ;
        RECT 513.920 20.440 514.180 20.700 ;
        RECT 517.140 20.440 517.400 20.700 ;
      LAYER met2 ;
        RECT 640.920 220.730 641.200 224.000 ;
        RECT 637.720 220.590 641.200 220.730 ;
        RECT 637.720 209.430 637.860 220.590 ;
        RECT 640.920 220.000 641.200 220.590 ;
        RECT 637.660 209.110 637.920 209.430 ;
        RECT 517.140 207.750 517.400 208.070 ;
        RECT 517.200 20.730 517.340 207.750 ;
        RECT 513.920 20.410 514.180 20.730 ;
        RECT 517.140 20.410 517.400 20.730 ;
        RECT 513.980 2.400 514.120 20.410 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 537.350 213.080 537.670 213.140 ;
        RECT 655.570 213.080 655.890 213.140 ;
        RECT 537.350 212.940 655.890 213.080 ;
        RECT 537.350 212.880 537.670 212.940 ;
        RECT 655.570 212.880 655.890 212.940 ;
        RECT 531.830 20.640 532.150 20.700 ;
        RECT 537.350 20.640 537.670 20.700 ;
        RECT 531.830 20.500 537.670 20.640 ;
        RECT 531.830 20.440 532.150 20.500 ;
        RECT 537.350 20.440 537.670 20.500 ;
      LAYER via ;
        RECT 537.380 212.880 537.640 213.140 ;
        RECT 655.600 212.880 655.860 213.140 ;
        RECT 531.860 20.440 532.120 20.700 ;
        RECT 537.380 20.440 537.640 20.700 ;
      LAYER met2 ;
        RECT 655.640 220.000 655.920 224.000 ;
        RECT 655.660 213.170 655.800 220.000 ;
        RECT 537.380 212.850 537.640 213.170 ;
        RECT 655.600 212.850 655.860 213.170 ;
        RECT 537.440 20.730 537.580 212.850 ;
        RECT 531.860 20.410 532.120 20.730 ;
        RECT 537.380 20.410 537.640 20.730 ;
        RECT 531.920 2.400 532.060 20.410 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 647.825 213.945 648.915 214.115 ;
        RECT 619.305 209.185 619.475 211.735 ;
        RECT 626.665 211.565 626.835 213.435 ;
        RECT 647.825 213.265 647.995 213.945 ;
      LAYER mcon ;
        RECT 648.745 213.945 648.915 214.115 ;
        RECT 626.665 213.265 626.835 213.435 ;
        RECT 619.305 211.565 619.475 211.735 ;
      LAYER met1 ;
        RECT 648.685 214.100 648.975 214.145 ;
        RECT 648.685 213.960 657.180 214.100 ;
        RECT 648.685 213.915 648.975 213.960 ;
        RECT 626.605 213.420 626.895 213.465 ;
        RECT 647.765 213.420 648.055 213.465 ;
        RECT 626.605 213.280 648.055 213.420 ;
        RECT 657.040 213.420 657.180 213.960 ;
        RECT 670.290 213.420 670.610 213.480 ;
        RECT 657.040 213.280 670.610 213.420 ;
        RECT 626.605 213.235 626.895 213.280 ;
        RECT 647.765 213.235 648.055 213.280 ;
        RECT 670.290 213.220 670.610 213.280 ;
        RECT 619.245 211.720 619.535 211.765 ;
        RECT 626.605 211.720 626.895 211.765 ;
        RECT 619.245 211.580 626.895 211.720 ;
        RECT 619.245 211.535 619.535 211.580 ;
        RECT 626.605 211.535 626.895 211.580 ;
        RECT 551.610 209.340 551.930 209.400 ;
        RECT 619.245 209.340 619.535 209.385 ;
        RECT 551.610 209.200 619.535 209.340 ;
        RECT 551.610 209.140 551.930 209.200 ;
        RECT 619.245 209.155 619.535 209.200 ;
        RECT 549.770 14.180 550.090 14.240 ;
        RECT 551.610 14.180 551.930 14.240 ;
        RECT 549.770 14.040 551.930 14.180 ;
        RECT 549.770 13.980 550.090 14.040 ;
        RECT 551.610 13.980 551.930 14.040 ;
      LAYER via ;
        RECT 670.320 213.220 670.580 213.480 ;
        RECT 551.640 209.140 551.900 209.400 ;
        RECT 549.800 13.980 550.060 14.240 ;
        RECT 551.640 13.980 551.900 14.240 ;
      LAYER met2 ;
        RECT 670.360 220.000 670.640 224.000 ;
        RECT 670.380 213.510 670.520 220.000 ;
        RECT 670.320 213.190 670.580 213.510 ;
        RECT 551.640 209.110 551.900 209.430 ;
        RECT 551.700 14.270 551.840 209.110 ;
        RECT 549.800 13.950 550.060 14.270 ;
        RECT 551.640 13.950 551.900 14.270 ;
        RECT 549.860 2.400 550.000 13.950 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 572.310 207.640 572.630 207.700 ;
        RECT 685.010 207.640 685.330 207.700 ;
        RECT 572.310 207.500 685.330 207.640 ;
        RECT 572.310 207.440 572.630 207.500 ;
        RECT 685.010 207.440 685.330 207.500 ;
        RECT 567.710 20.640 568.030 20.700 ;
        RECT 572.310 20.640 572.630 20.700 ;
        RECT 567.710 20.500 572.630 20.640 ;
        RECT 567.710 20.440 568.030 20.500 ;
        RECT 572.310 20.440 572.630 20.500 ;
      LAYER via ;
        RECT 572.340 207.440 572.600 207.700 ;
        RECT 685.040 207.440 685.300 207.700 ;
        RECT 567.740 20.440 568.000 20.700 ;
        RECT 572.340 20.440 572.600 20.700 ;
      LAYER met2 ;
        RECT 685.080 220.000 685.360 224.000 ;
        RECT 685.100 207.730 685.240 220.000 ;
        RECT 572.340 207.410 572.600 207.730 ;
        RECT 685.040 207.410 685.300 207.730 ;
        RECT 572.400 20.730 572.540 207.410 ;
        RECT 567.740 20.410 568.000 20.730 ;
        RECT 572.340 20.410 572.600 20.730 ;
        RECT 567.800 2.400 567.940 20.410 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 587.580 210.900 627.740 211.040 ;
        RECT 585.650 210.700 585.970 210.760 ;
        RECT 587.580 210.700 587.720 210.900 ;
        RECT 585.650 210.560 587.720 210.700 ;
        RECT 585.650 210.500 585.970 210.560 ;
        RECT 627.600 210.360 627.740 210.900 ;
        RECT 699.730 210.360 700.050 210.420 ;
        RECT 627.600 210.220 700.050 210.360 ;
        RECT 699.730 210.160 700.050 210.220 ;
      LAYER via ;
        RECT 585.680 210.500 585.940 210.760 ;
        RECT 699.760 210.160 700.020 210.420 ;
      LAYER met2 ;
        RECT 699.800 220.000 700.080 224.000 ;
        RECT 585.680 210.470 585.940 210.790 ;
        RECT 585.740 2.400 585.880 210.470 ;
        RECT 699.820 210.450 699.960 220.000 ;
        RECT 699.760 210.130 700.020 210.450 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 96.210 213.080 96.530 213.140 ;
        RECT 293.090 213.080 293.410 213.140 ;
        RECT 96.210 212.940 293.410 213.080 ;
        RECT 96.210 212.880 96.530 212.940 ;
        RECT 293.090 212.880 293.410 212.940 ;
        RECT 91.610 20.640 91.930 20.700 ;
        RECT 96.210 20.640 96.530 20.700 ;
        RECT 91.610 20.500 96.530 20.640 ;
        RECT 91.610 20.440 91.930 20.500 ;
        RECT 96.210 20.440 96.530 20.500 ;
      LAYER via ;
        RECT 96.240 212.880 96.500 213.140 ;
        RECT 293.120 212.880 293.380 213.140 ;
        RECT 91.640 20.440 91.900 20.700 ;
        RECT 96.240 20.440 96.500 20.700 ;
      LAYER met2 ;
        RECT 293.160 220.000 293.440 224.000 ;
        RECT 293.180 213.170 293.320 220.000 ;
        RECT 96.240 212.850 96.500 213.170 ;
        RECT 293.120 212.850 293.380 213.170 ;
        RECT 96.300 20.730 96.440 212.850 ;
        RECT 91.640 20.410 91.900 20.730 ;
        RECT 96.240 20.410 96.500 20.730 ;
        RECT 91.700 2.400 91.840 20.410 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 714.450 212.740 714.770 212.800 ;
        RECT 611.960 212.600 714.770 212.740 ;
        RECT 606.810 212.400 607.130 212.460 ;
        RECT 611.960 212.400 612.100 212.600 ;
        RECT 714.450 212.540 714.770 212.600 ;
        RECT 606.810 212.260 612.100 212.400 ;
        RECT 606.810 212.200 607.130 212.260 ;
        RECT 603.130 16.900 603.450 16.960 ;
        RECT 606.810 16.900 607.130 16.960 ;
        RECT 603.130 16.760 607.130 16.900 ;
        RECT 603.130 16.700 603.450 16.760 ;
        RECT 606.810 16.700 607.130 16.760 ;
      LAYER via ;
        RECT 606.840 212.200 607.100 212.460 ;
        RECT 714.480 212.540 714.740 212.800 ;
        RECT 603.160 16.700 603.420 16.960 ;
        RECT 606.840 16.700 607.100 16.960 ;
      LAYER met2 ;
        RECT 714.520 220.000 714.800 224.000 ;
        RECT 714.540 212.830 714.680 220.000 ;
        RECT 714.480 212.510 714.740 212.830 ;
        RECT 606.840 212.170 607.100 212.490 ;
        RECT 606.900 16.990 607.040 212.170 ;
        RECT 603.160 16.670 603.420 16.990 ;
        RECT 606.840 16.670 607.100 16.990 ;
        RECT 603.220 2.400 603.360 16.670 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 627.050 211.720 627.370 211.780 ;
        RECT 729.170 211.720 729.490 211.780 ;
        RECT 627.050 211.580 729.490 211.720 ;
        RECT 627.050 211.520 627.370 211.580 ;
        RECT 729.170 211.520 729.490 211.580 ;
        RECT 621.070 15.880 621.390 15.940 ;
        RECT 627.050 15.880 627.370 15.940 ;
        RECT 621.070 15.740 627.370 15.880 ;
        RECT 621.070 15.680 621.390 15.740 ;
        RECT 627.050 15.680 627.370 15.740 ;
      LAYER via ;
        RECT 627.080 211.520 627.340 211.780 ;
        RECT 729.200 211.520 729.460 211.780 ;
        RECT 621.100 15.680 621.360 15.940 ;
        RECT 627.080 15.680 627.340 15.940 ;
      LAYER met2 ;
        RECT 729.240 220.000 729.520 224.000 ;
        RECT 729.260 211.810 729.400 220.000 ;
        RECT 627.080 211.490 627.340 211.810 ;
        RECT 729.200 211.490 729.460 211.810 ;
        RECT 627.140 15.970 627.280 211.490 ;
        RECT 621.100 15.650 621.360 15.970 ;
        RECT 627.080 15.650 627.340 15.970 ;
        RECT 621.160 2.400 621.300 15.650 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 116.910 213.420 117.230 213.480 ;
        RECT 312.870 213.420 313.190 213.480 ;
        RECT 116.910 213.280 313.190 213.420 ;
        RECT 116.910 213.220 117.230 213.280 ;
        RECT 312.870 213.220 313.190 213.280 ;
        RECT 115.530 14.180 115.850 14.240 ;
        RECT 116.910 14.180 117.230 14.240 ;
        RECT 115.530 14.040 117.230 14.180 ;
        RECT 115.530 13.980 115.850 14.040 ;
        RECT 116.910 13.980 117.230 14.040 ;
      LAYER via ;
        RECT 116.940 213.220 117.200 213.480 ;
        RECT 312.900 213.220 313.160 213.480 ;
        RECT 115.560 13.980 115.820 14.240 ;
        RECT 116.940 13.980 117.200 14.240 ;
      LAYER met2 ;
        RECT 312.940 220.000 313.220 224.000 ;
        RECT 312.960 213.510 313.100 220.000 ;
        RECT 116.940 213.190 117.200 213.510 ;
        RECT 312.900 213.190 313.160 213.510 ;
        RECT 117.000 14.270 117.140 213.190 ;
        RECT 115.560 13.950 115.820 14.270 ;
        RECT 116.940 13.950 117.200 14.270 ;
        RECT 115.620 2.400 115.760 13.950 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 299.145 209.525 299.315 212.755 ;
      LAYER mcon ;
        RECT 299.145 212.585 299.315 212.755 ;
      LAYER met1 ;
        RECT 299.085 212.740 299.375 212.785 ;
        RECT 330.810 212.740 331.130 212.800 ;
        RECT 299.085 212.600 331.130 212.740 ;
        RECT 299.085 212.555 299.375 212.600 ;
        RECT 330.810 212.540 331.130 212.600 ;
        RECT 144.510 209.680 144.830 209.740 ;
        RECT 299.085 209.680 299.375 209.725 ;
        RECT 144.510 209.540 299.375 209.680 ;
        RECT 144.510 209.480 144.830 209.540 ;
        RECT 299.085 209.495 299.375 209.540 ;
        RECT 139.450 18.600 139.770 18.660 ;
        RECT 144.510 18.600 144.830 18.660 ;
        RECT 139.450 18.460 144.830 18.600 ;
        RECT 139.450 18.400 139.770 18.460 ;
        RECT 144.510 18.400 144.830 18.460 ;
      LAYER via ;
        RECT 330.840 212.540 331.100 212.800 ;
        RECT 144.540 209.480 144.800 209.740 ;
        RECT 139.480 18.400 139.740 18.660 ;
        RECT 144.540 18.400 144.800 18.660 ;
      LAYER met2 ;
        RECT 332.260 220.730 332.540 224.000 ;
        RECT 331.360 220.590 332.540 220.730 ;
        RECT 330.840 212.570 331.100 212.830 ;
        RECT 331.360 212.570 331.500 220.590 ;
        RECT 332.260 220.000 332.540 220.590 ;
        RECT 330.840 212.510 331.500 212.570 ;
        RECT 330.900 212.430 331.500 212.510 ;
        RECT 144.540 209.450 144.800 209.770 ;
        RECT 144.600 18.690 144.740 209.450 ;
        RECT 139.480 18.370 139.740 18.690 ;
        RECT 144.540 18.370 144.800 18.690 ;
        RECT 139.540 2.400 139.680 18.370 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 337.785 209.865 337.955 213.775 ;
        RECT 158.385 144.925 158.555 193.035 ;
        RECT 157.465 2.805 157.635 48.195 ;
      LAYER mcon ;
        RECT 337.785 213.605 337.955 213.775 ;
        RECT 158.385 192.865 158.555 193.035 ;
        RECT 157.465 48.025 157.635 48.195 ;
      LAYER met1 ;
        RECT 345.070 214.100 345.390 214.160 ;
        RECT 344.240 213.960 345.390 214.100 ;
        RECT 337.725 213.760 338.015 213.805 ;
        RECT 344.240 213.760 344.380 213.960 ;
        RECT 345.070 213.900 345.390 213.960 ;
        RECT 337.725 213.620 344.380 213.760 ;
        RECT 337.725 213.575 338.015 213.620 ;
        RECT 158.310 210.020 158.630 210.080 ;
        RECT 337.725 210.020 338.015 210.065 ;
        RECT 158.310 209.880 338.015 210.020 ;
        RECT 158.310 209.820 158.630 209.880 ;
        RECT 337.725 209.835 338.015 209.880 ;
        RECT 158.310 193.020 158.630 193.080 ;
        RECT 158.115 192.880 158.630 193.020 ;
        RECT 158.310 192.820 158.630 192.880 ;
        RECT 158.310 145.080 158.630 145.140 ;
        RECT 158.115 144.940 158.630 145.080 ;
        RECT 158.310 144.880 158.630 144.940 ;
        RECT 157.390 96.460 157.710 96.520 ;
        RECT 158.310 96.460 158.630 96.520 ;
        RECT 157.390 96.320 158.630 96.460 ;
        RECT 157.390 96.260 157.710 96.320 ;
        RECT 158.310 96.260 158.630 96.320 ;
        RECT 157.405 48.180 157.695 48.225 ;
        RECT 158.310 48.180 158.630 48.240 ;
        RECT 157.405 48.040 158.630 48.180 ;
        RECT 157.405 47.995 157.695 48.040 ;
        RECT 158.310 47.980 158.630 48.040 ;
        RECT 157.390 2.960 157.710 3.020 ;
        RECT 157.195 2.820 157.710 2.960 ;
        RECT 157.390 2.760 157.710 2.820 ;
      LAYER via ;
        RECT 345.100 213.900 345.360 214.160 ;
        RECT 158.340 209.820 158.600 210.080 ;
        RECT 158.340 192.820 158.600 193.080 ;
        RECT 158.340 144.880 158.600 145.140 ;
        RECT 157.420 96.260 157.680 96.520 ;
        RECT 158.340 96.260 158.600 96.520 ;
        RECT 158.340 47.980 158.600 48.240 ;
        RECT 157.420 2.760 157.680 3.020 ;
      LAYER met2 ;
        RECT 346.980 220.730 347.260 224.000 ;
        RECT 345.160 220.590 347.260 220.730 ;
        RECT 345.160 214.190 345.300 220.590 ;
        RECT 346.980 220.000 347.260 220.590 ;
        RECT 345.100 213.870 345.360 214.190 ;
        RECT 158.340 209.790 158.600 210.110 ;
        RECT 158.400 193.110 158.540 209.790 ;
        RECT 158.340 192.790 158.600 193.110 ;
        RECT 158.340 144.850 158.600 145.170 ;
        RECT 158.400 96.550 158.540 144.850 ;
        RECT 157.420 96.230 157.680 96.550 ;
        RECT 158.340 96.230 158.600 96.550 ;
        RECT 157.480 48.805 157.620 96.230 ;
        RECT 157.410 48.435 157.690 48.805 ;
        RECT 158.330 48.435 158.610 48.805 ;
        RECT 158.400 48.270 158.540 48.435 ;
        RECT 158.340 47.950 158.600 48.270 ;
        RECT 157.420 2.730 157.680 3.050 ;
        RECT 157.480 2.400 157.620 2.730 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 157.410 48.480 157.690 48.760 ;
        RECT 158.330 48.480 158.610 48.760 ;
      LAYER met3 ;
        RECT 157.385 48.770 157.715 48.785 ;
        RECT 158.305 48.770 158.635 48.785 ;
        RECT 157.385 48.470 158.635 48.770 ;
        RECT 157.385 48.455 157.715 48.470 ;
        RECT 158.305 48.455 158.635 48.470 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 334.105 208.845 334.275 213.095 ;
      LAYER mcon ;
        RECT 334.105 212.925 334.275 213.095 ;
      LAYER met1 ;
        RECT 334.045 213.080 334.335 213.125 ;
        RECT 361.630 213.080 361.950 213.140 ;
        RECT 334.045 212.940 361.950 213.080 ;
        RECT 334.045 212.895 334.335 212.940 ;
        RECT 361.630 212.880 361.950 212.940 ;
        RECT 179.010 209.000 179.330 209.060 ;
        RECT 334.045 209.000 334.335 209.045 ;
        RECT 179.010 208.860 334.335 209.000 ;
        RECT 179.010 208.800 179.330 208.860 ;
        RECT 334.045 208.815 334.335 208.860 ;
        RECT 174.870 16.900 175.190 16.960 ;
        RECT 179.010 16.900 179.330 16.960 ;
        RECT 174.870 16.760 179.330 16.900 ;
        RECT 174.870 16.700 175.190 16.760 ;
        RECT 179.010 16.700 179.330 16.760 ;
      LAYER via ;
        RECT 361.660 212.880 361.920 213.140 ;
        RECT 179.040 208.800 179.300 209.060 ;
        RECT 174.900 16.700 175.160 16.960 ;
        RECT 179.040 16.700 179.300 16.960 ;
      LAYER met2 ;
        RECT 361.700 220.000 361.980 224.000 ;
        RECT 361.720 213.170 361.860 220.000 ;
        RECT 361.660 212.850 361.920 213.170 ;
        RECT 179.040 208.770 179.300 209.090 ;
        RECT 179.100 16.990 179.240 208.770 ;
        RECT 174.900 16.670 175.160 16.990 ;
        RECT 179.040 16.670 179.300 16.990 ;
        RECT 174.960 2.400 175.100 16.670 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.350 209.340 192.670 209.400 ;
        RECT 376.350 209.340 376.670 209.400 ;
        RECT 192.350 209.200 376.670 209.340 ;
        RECT 192.350 209.140 192.670 209.200 ;
        RECT 376.350 209.140 376.670 209.200 ;
      LAYER via ;
        RECT 192.380 209.140 192.640 209.400 ;
        RECT 376.380 209.140 376.640 209.400 ;
      LAYER met2 ;
        RECT 376.420 220.000 376.700 224.000 ;
        RECT 376.440 209.430 376.580 220.000 ;
        RECT 192.380 209.110 192.640 209.430 ;
        RECT 376.380 209.110 376.640 209.430 ;
        RECT 192.440 3.130 192.580 209.110 ;
        RECT 192.440 2.990 193.040 3.130 ;
        RECT 192.900 2.400 193.040 2.990 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 213.510 208.660 213.830 208.720 ;
        RECT 391.070 208.660 391.390 208.720 ;
        RECT 213.510 208.520 391.390 208.660 ;
        RECT 213.510 208.460 213.830 208.520 ;
        RECT 391.070 208.460 391.390 208.520 ;
        RECT 210.750 16.560 211.070 16.620 ;
        RECT 213.510 16.560 213.830 16.620 ;
        RECT 210.750 16.420 213.830 16.560 ;
        RECT 210.750 16.360 211.070 16.420 ;
        RECT 213.510 16.360 213.830 16.420 ;
      LAYER via ;
        RECT 213.540 208.460 213.800 208.720 ;
        RECT 391.100 208.460 391.360 208.720 ;
        RECT 210.780 16.360 211.040 16.620 ;
        RECT 213.540 16.360 213.800 16.620 ;
      LAYER met2 ;
        RECT 391.140 220.000 391.420 224.000 ;
        RECT 391.160 208.750 391.300 220.000 ;
        RECT 213.540 208.430 213.800 208.750 ;
        RECT 391.100 208.430 391.360 208.750 ;
        RECT 213.600 16.650 213.740 208.430 ;
        RECT 210.780 16.330 211.040 16.650 ;
        RECT 213.540 16.330 213.800 16.650 ;
        RECT 210.840 2.400 210.980 16.330 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 234.670 210.700 234.990 210.760 ;
        RECT 405.790 210.700 406.110 210.760 ;
        RECT 234.670 210.560 406.110 210.700 ;
        RECT 234.670 210.500 234.990 210.560 ;
        RECT 405.790 210.500 406.110 210.560 ;
        RECT 228.690 17.580 229.010 17.640 ;
        RECT 234.210 17.580 234.530 17.640 ;
        RECT 228.690 17.440 234.530 17.580 ;
        RECT 228.690 17.380 229.010 17.440 ;
        RECT 234.210 17.380 234.530 17.440 ;
      LAYER via ;
        RECT 234.700 210.500 234.960 210.760 ;
        RECT 405.820 210.500 406.080 210.760 ;
        RECT 228.720 17.380 228.980 17.640 ;
        RECT 234.240 17.380 234.500 17.640 ;
      LAYER met2 ;
        RECT 405.860 220.000 406.140 224.000 ;
        RECT 405.880 210.790 406.020 220.000 ;
        RECT 234.700 210.470 234.960 210.790 ;
        RECT 405.820 210.470 406.080 210.790 ;
        RECT 234.760 209.850 234.900 210.470 ;
        RECT 234.300 209.710 234.900 209.850 ;
        RECT 234.300 17.670 234.440 209.710 ;
        RECT 228.720 17.350 228.980 17.670 ;
        RECT 234.240 17.350 234.500 17.670 ;
        RECT 228.780 2.400 228.920 17.350 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 54.810 211.040 55.130 211.100 ;
        RECT 259.050 211.040 259.370 211.100 ;
        RECT 54.810 210.900 259.370 211.040 ;
        RECT 54.810 210.840 55.130 210.900 ;
        RECT 259.050 210.840 259.370 210.900 ;
        RECT 50.210 16.900 50.530 16.960 ;
        RECT 54.810 16.900 55.130 16.960 ;
        RECT 50.210 16.760 55.130 16.900 ;
        RECT 50.210 16.700 50.530 16.760 ;
        RECT 54.810 16.700 55.130 16.760 ;
      LAYER via ;
        RECT 54.840 210.840 55.100 211.100 ;
        RECT 259.080 210.840 259.340 211.100 ;
        RECT 50.240 16.700 50.500 16.960 ;
        RECT 54.840 16.700 55.100 16.960 ;
      LAYER met2 ;
        RECT 259.120 220.000 259.400 224.000 ;
        RECT 259.140 211.130 259.280 220.000 ;
        RECT 54.840 210.810 55.100 211.130 ;
        RECT 259.080 210.810 259.340 211.130 ;
        RECT 54.900 16.990 55.040 210.810 ;
        RECT 50.240 16.670 50.500 16.990 ;
        RECT 54.840 16.670 55.100 16.990 ;
        RECT 50.300 2.400 50.440 16.670 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 300.065 210.205 300.235 212.415 ;
      LAYER mcon ;
        RECT 300.065 212.245 300.235 212.415 ;
      LAYER met1 ;
        RECT 254.910 212.400 255.230 212.460 ;
        RECT 300.005 212.400 300.295 212.445 ;
        RECT 254.910 212.260 300.295 212.400 ;
        RECT 254.910 212.200 255.230 212.260 ;
        RECT 300.005 212.215 300.295 212.260 ;
        RECT 300.005 210.360 300.295 210.405 ;
        RECT 425.570 210.360 425.890 210.420 ;
        RECT 300.005 210.220 425.890 210.360 ;
        RECT 300.005 210.175 300.295 210.220 ;
        RECT 425.570 210.160 425.890 210.220 ;
        RECT 252.610 17.580 252.930 17.640 ;
        RECT 254.910 17.580 255.230 17.640 ;
        RECT 252.610 17.440 255.230 17.580 ;
        RECT 252.610 17.380 252.930 17.440 ;
        RECT 254.910 17.380 255.230 17.440 ;
      LAYER via ;
        RECT 254.940 212.200 255.200 212.460 ;
        RECT 425.600 210.160 425.860 210.420 ;
        RECT 252.640 17.380 252.900 17.640 ;
        RECT 254.940 17.380 255.200 17.640 ;
      LAYER met2 ;
        RECT 425.640 220.000 425.920 224.000 ;
        RECT 254.940 212.170 255.200 212.490 ;
        RECT 255.000 17.670 255.140 212.170 ;
        RECT 425.660 210.450 425.800 220.000 ;
        RECT 425.600 210.130 425.860 210.450 ;
        RECT 252.640 17.350 252.900 17.670 ;
        RECT 254.940 17.350 255.200 17.670 ;
        RECT 252.700 2.400 252.840 17.350 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 275.610 212.060 275.930 212.120 ;
        RECT 440.290 212.060 440.610 212.120 ;
        RECT 275.610 211.920 440.610 212.060 ;
        RECT 275.610 211.860 275.930 211.920 ;
        RECT 440.290 211.860 440.610 211.920 ;
        RECT 270.090 20.640 270.410 20.700 ;
        RECT 275.610 20.640 275.930 20.700 ;
        RECT 270.090 20.500 275.930 20.640 ;
        RECT 270.090 20.440 270.410 20.500 ;
        RECT 275.610 20.440 275.930 20.500 ;
      LAYER via ;
        RECT 275.640 211.860 275.900 212.120 ;
        RECT 440.320 211.860 440.580 212.120 ;
        RECT 270.120 20.440 270.380 20.700 ;
        RECT 275.640 20.440 275.900 20.700 ;
      LAYER met2 ;
        RECT 440.360 220.000 440.640 224.000 ;
        RECT 440.380 212.150 440.520 220.000 ;
        RECT 275.640 211.830 275.900 212.150 ;
        RECT 440.320 211.830 440.580 212.150 ;
        RECT 275.700 20.730 275.840 211.830 ;
        RECT 270.120 20.410 270.380 20.730 ;
        RECT 275.640 20.410 275.900 20.730 ;
        RECT 270.180 2.400 270.320 20.410 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 300.525 211.565 300.695 212.415 ;
        RECT 288.105 2.805 288.275 14.195 ;
      LAYER mcon ;
        RECT 300.525 212.245 300.695 212.415 ;
        RECT 288.105 14.025 288.275 14.195 ;
      LAYER met1 ;
        RECT 300.465 212.400 300.755 212.445 ;
        RECT 455.010 212.400 455.330 212.460 ;
        RECT 300.465 212.260 455.330 212.400 ;
        RECT 300.465 212.215 300.755 212.260 ;
        RECT 455.010 212.200 455.330 212.260 ;
        RECT 289.410 211.720 289.730 211.780 ;
        RECT 300.465 211.720 300.755 211.765 ;
        RECT 289.410 211.580 300.755 211.720 ;
        RECT 289.410 211.520 289.730 211.580 ;
        RECT 300.465 211.535 300.755 211.580 ;
        RECT 288.045 14.180 288.335 14.225 ;
        RECT 289.410 14.180 289.730 14.240 ;
        RECT 288.045 14.040 289.730 14.180 ;
        RECT 288.045 13.995 288.335 14.040 ;
        RECT 289.410 13.980 289.730 14.040 ;
        RECT 288.030 2.960 288.350 3.020 ;
        RECT 287.835 2.820 288.350 2.960 ;
        RECT 288.030 2.760 288.350 2.820 ;
      LAYER via ;
        RECT 455.040 212.200 455.300 212.460 ;
        RECT 289.440 211.520 289.700 211.780 ;
        RECT 289.440 13.980 289.700 14.240 ;
        RECT 288.060 2.760 288.320 3.020 ;
      LAYER met2 ;
        RECT 455.080 220.000 455.360 224.000 ;
        RECT 455.100 212.490 455.240 220.000 ;
        RECT 455.040 212.170 455.300 212.490 ;
        RECT 289.440 211.490 289.700 211.810 ;
        RECT 289.500 14.270 289.640 211.490 ;
        RECT 289.440 13.950 289.700 14.270 ;
        RECT 288.060 2.730 288.320 3.050 ;
        RECT 288.120 2.400 288.260 2.730 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 310.110 211.720 310.430 211.780 ;
        RECT 469.270 211.720 469.590 211.780 ;
        RECT 310.110 211.580 469.590 211.720 ;
        RECT 310.110 211.520 310.430 211.580 ;
        RECT 469.270 211.520 469.590 211.580 ;
        RECT 305.970 17.240 306.290 17.300 ;
        RECT 310.110 17.240 310.430 17.300 ;
        RECT 305.970 17.100 310.430 17.240 ;
        RECT 305.970 17.040 306.290 17.100 ;
        RECT 310.110 17.040 310.430 17.100 ;
      LAYER via ;
        RECT 310.140 211.520 310.400 211.780 ;
        RECT 469.300 211.520 469.560 211.780 ;
        RECT 306.000 17.040 306.260 17.300 ;
        RECT 310.140 17.040 310.400 17.300 ;
      LAYER met2 ;
        RECT 469.340 220.000 469.620 224.000 ;
        RECT 469.360 211.810 469.500 220.000 ;
        RECT 310.140 211.490 310.400 211.810 ;
        RECT 469.300 211.490 469.560 211.810 ;
        RECT 310.200 17.330 310.340 211.490 ;
        RECT 306.000 17.010 306.260 17.330 ;
        RECT 310.140 17.010 310.400 17.330 ;
        RECT 306.060 2.400 306.200 17.010 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 347.445 208.845 347.615 209.695 ;
      LAYER mcon ;
        RECT 347.445 209.525 347.615 209.695 ;
      LAYER met1 ;
        RECT 347.385 209.680 347.675 209.725 ;
        RECT 483.990 209.680 484.310 209.740 ;
        RECT 347.385 209.540 484.310 209.680 ;
        RECT 347.385 209.495 347.675 209.540 ;
        RECT 483.990 209.480 484.310 209.540 ;
        RECT 334.490 209.000 334.810 209.060 ;
        RECT 347.385 209.000 347.675 209.045 ;
        RECT 334.490 208.860 347.675 209.000 ;
        RECT 334.490 208.800 334.810 208.860 ;
        RECT 347.385 208.815 347.675 208.860 ;
        RECT 323.910 15.540 324.230 15.600 ;
        RECT 334.490 15.540 334.810 15.600 ;
        RECT 323.910 15.400 334.810 15.540 ;
        RECT 323.910 15.340 324.230 15.400 ;
        RECT 334.490 15.340 334.810 15.400 ;
      LAYER via ;
        RECT 484.020 209.480 484.280 209.740 ;
        RECT 334.520 208.800 334.780 209.060 ;
        RECT 323.940 15.340 324.200 15.600 ;
        RECT 334.520 15.340 334.780 15.600 ;
      LAYER met2 ;
        RECT 484.060 220.000 484.340 224.000 ;
        RECT 484.080 209.770 484.220 220.000 ;
        RECT 484.020 209.450 484.280 209.770 ;
        RECT 334.520 208.770 334.780 209.090 ;
        RECT 334.580 15.630 334.720 208.770 ;
        RECT 323.940 15.310 324.200 15.630 ;
        RECT 334.520 15.310 334.780 15.630 ;
        RECT 324.000 2.400 324.140 15.310 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 372.285 212.925 372.455 214.115 ;
      LAYER mcon ;
        RECT 372.285 213.945 372.455 214.115 ;
      LAYER met1 ;
        RECT 372.225 214.100 372.515 214.145 ;
        RECT 371.380 213.960 372.515 214.100 ;
        RECT 344.610 213.760 344.930 213.820 ;
        RECT 371.380 213.760 371.520 213.960 ;
        RECT 372.225 213.915 372.515 213.960 ;
        RECT 344.610 213.620 371.520 213.760 ;
        RECT 344.610 213.560 344.930 213.620 ;
        RECT 372.225 213.080 372.515 213.125 ;
        RECT 498.710 213.080 499.030 213.140 ;
        RECT 372.225 212.940 499.030 213.080 ;
        RECT 372.225 212.895 372.515 212.940 ;
        RECT 498.710 212.880 499.030 212.940 ;
        RECT 341.390 17.240 341.710 17.300 ;
        RECT 344.610 17.240 344.930 17.300 ;
        RECT 341.390 17.100 344.930 17.240 ;
        RECT 341.390 17.040 341.710 17.100 ;
        RECT 344.610 17.040 344.930 17.100 ;
      LAYER via ;
        RECT 344.640 213.560 344.900 213.820 ;
        RECT 498.740 212.880 499.000 213.140 ;
        RECT 341.420 17.040 341.680 17.300 ;
        RECT 344.640 17.040 344.900 17.300 ;
      LAYER met2 ;
        RECT 498.780 220.000 499.060 224.000 ;
        RECT 344.640 213.530 344.900 213.850 ;
        RECT 344.700 17.330 344.840 213.530 ;
        RECT 498.800 213.170 498.940 220.000 ;
        RECT 498.740 212.850 499.000 213.170 ;
        RECT 341.420 17.010 341.680 17.330 ;
        RECT 344.640 17.010 344.900 17.330 ;
        RECT 341.480 2.400 341.620 17.010 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 368.990 207.980 369.310 208.040 ;
        RECT 513.430 207.980 513.750 208.040 ;
        RECT 368.990 207.840 513.750 207.980 ;
        RECT 368.990 207.780 369.310 207.840 ;
        RECT 513.430 207.780 513.750 207.840 ;
        RECT 359.330 20.640 359.650 20.700 ;
        RECT 368.990 20.640 369.310 20.700 ;
        RECT 359.330 20.500 369.310 20.640 ;
        RECT 359.330 20.440 359.650 20.500 ;
        RECT 368.990 20.440 369.310 20.500 ;
      LAYER via ;
        RECT 369.020 207.780 369.280 208.040 ;
        RECT 513.460 207.780 513.720 208.040 ;
        RECT 359.360 20.440 359.620 20.700 ;
        RECT 369.020 20.440 369.280 20.700 ;
      LAYER met2 ;
        RECT 513.500 220.000 513.780 224.000 ;
        RECT 513.520 208.070 513.660 220.000 ;
        RECT 369.020 207.750 369.280 208.070 ;
        RECT 513.460 207.750 513.720 208.070 ;
        RECT 369.080 20.730 369.220 207.750 ;
        RECT 359.360 20.410 359.620 20.730 ;
        RECT 369.020 20.410 369.280 20.730 ;
        RECT 359.420 2.400 359.560 20.410 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 378.725 138.125 378.895 186.235 ;
        RECT 377.345 48.365 377.515 104.975 ;
      LAYER mcon ;
        RECT 378.725 186.065 378.895 186.235 ;
        RECT 377.345 104.805 377.515 104.975 ;
      LAYER met1 ;
        RECT 379.110 210.020 379.430 210.080 ;
        RECT 528.150 210.020 528.470 210.080 ;
        RECT 379.110 209.880 528.470 210.020 ;
        RECT 379.110 209.820 379.430 209.880 ;
        RECT 528.150 209.820 528.470 209.880 ;
        RECT 378.650 193.020 378.970 193.080 ;
        RECT 379.110 193.020 379.430 193.080 ;
        RECT 378.650 192.880 379.430 193.020 ;
        RECT 378.650 192.820 378.970 192.880 ;
        RECT 379.110 192.820 379.430 192.880 ;
        RECT 378.650 186.220 378.970 186.280 ;
        RECT 378.650 186.080 379.165 186.220 ;
        RECT 378.650 186.020 378.970 186.080 ;
        RECT 378.665 138.280 378.955 138.325 ;
        RECT 379.110 138.280 379.430 138.340 ;
        RECT 378.665 138.140 379.430 138.280 ;
        RECT 378.665 138.095 378.955 138.140 ;
        RECT 379.110 138.080 379.430 138.140 ;
        RECT 377.285 104.960 377.575 105.005 ;
        RECT 379.110 104.960 379.430 105.020 ;
        RECT 377.285 104.820 379.430 104.960 ;
        RECT 377.285 104.775 377.575 104.820 ;
        RECT 379.110 104.760 379.430 104.820 ;
        RECT 377.270 48.520 377.590 48.580 ;
        RECT 377.075 48.380 377.590 48.520 ;
        RECT 377.270 48.320 377.590 48.380 ;
      LAYER via ;
        RECT 379.140 209.820 379.400 210.080 ;
        RECT 528.180 209.820 528.440 210.080 ;
        RECT 378.680 192.820 378.940 193.080 ;
        RECT 379.140 192.820 379.400 193.080 ;
        RECT 378.680 186.020 378.940 186.280 ;
        RECT 379.140 138.080 379.400 138.340 ;
        RECT 379.140 104.760 379.400 105.020 ;
        RECT 377.300 48.320 377.560 48.580 ;
      LAYER met2 ;
        RECT 528.220 220.000 528.500 224.000 ;
        RECT 528.240 210.110 528.380 220.000 ;
        RECT 379.140 209.790 379.400 210.110 ;
        RECT 528.180 209.790 528.440 210.110 ;
        RECT 379.200 193.110 379.340 209.790 ;
        RECT 378.680 192.790 378.940 193.110 ;
        RECT 379.140 192.790 379.400 193.110 ;
        RECT 378.740 186.310 378.880 192.790 ;
        RECT 378.680 185.990 378.940 186.310 ;
        RECT 379.140 138.050 379.400 138.370 ;
        RECT 379.200 105.050 379.340 138.050 ;
        RECT 379.140 104.730 379.400 105.050 ;
        RECT 377.300 48.290 377.560 48.610 ;
        RECT 377.360 2.400 377.500 48.290 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 399.810 208.660 400.130 208.720 ;
        RECT 542.870 208.660 543.190 208.720 ;
        RECT 399.810 208.520 543.190 208.660 ;
        RECT 399.810 208.460 400.130 208.520 ;
        RECT 542.870 208.460 543.190 208.520 ;
        RECT 395.210 18.940 395.530 19.000 ;
        RECT 399.810 18.940 400.130 19.000 ;
        RECT 395.210 18.800 400.130 18.940 ;
        RECT 395.210 18.740 395.530 18.800 ;
        RECT 399.810 18.740 400.130 18.800 ;
      LAYER via ;
        RECT 399.840 208.460 400.100 208.720 ;
        RECT 542.900 208.460 543.160 208.720 ;
        RECT 395.240 18.740 395.500 19.000 ;
        RECT 399.840 18.740 400.100 19.000 ;
      LAYER met2 ;
        RECT 542.940 220.000 543.220 224.000 ;
        RECT 542.960 208.750 543.100 220.000 ;
        RECT 399.840 208.430 400.100 208.750 ;
        RECT 542.900 208.430 543.160 208.750 ;
        RECT 399.900 19.030 400.040 208.430 ;
        RECT 395.240 18.710 395.500 19.030 ;
        RECT 399.840 18.710 400.100 19.030 ;
        RECT 395.300 2.400 395.440 18.710 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 417.290 208.320 417.610 208.380 ;
        RECT 557.590 208.320 557.910 208.380 ;
        RECT 417.290 208.180 557.910 208.320 ;
        RECT 417.290 208.120 417.610 208.180 ;
        RECT 557.590 208.120 557.910 208.180 ;
        RECT 413.150 19.280 413.470 19.340 ;
        RECT 417.290 19.280 417.610 19.340 ;
        RECT 413.150 19.140 417.610 19.280 ;
        RECT 413.150 19.080 413.470 19.140 ;
        RECT 417.290 19.080 417.610 19.140 ;
      LAYER via ;
        RECT 417.320 208.120 417.580 208.380 ;
        RECT 557.620 208.120 557.880 208.380 ;
        RECT 413.180 19.080 413.440 19.340 ;
        RECT 417.320 19.080 417.580 19.340 ;
      LAYER met2 ;
        RECT 557.660 220.000 557.940 224.000 ;
        RECT 557.680 208.410 557.820 220.000 ;
        RECT 417.320 208.090 417.580 208.410 ;
        RECT 557.620 208.090 557.880 208.410 ;
        RECT 417.380 19.370 417.520 208.090 ;
        RECT 413.180 19.050 413.440 19.370 ;
        RECT 417.320 19.050 417.580 19.370 ;
        RECT 413.240 2.400 413.380 19.050 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 251.690 207.640 252.010 207.700 ;
        RECT 278.370 207.640 278.690 207.700 ;
        RECT 251.690 207.500 278.690 207.640 ;
        RECT 251.690 207.440 252.010 207.500 ;
        RECT 278.370 207.440 278.690 207.500 ;
        RECT 74.130 19.280 74.450 19.340 ;
        RECT 251.690 19.280 252.010 19.340 ;
        RECT 74.130 19.140 252.010 19.280 ;
        RECT 74.130 19.080 74.450 19.140 ;
        RECT 251.690 19.080 252.010 19.140 ;
      LAYER via ;
        RECT 251.720 207.440 251.980 207.700 ;
        RECT 278.400 207.440 278.660 207.700 ;
        RECT 74.160 19.080 74.420 19.340 ;
        RECT 251.720 19.080 251.980 19.340 ;
      LAYER met2 ;
        RECT 278.440 220.000 278.720 224.000 ;
        RECT 278.460 207.730 278.600 220.000 ;
        RECT 251.720 207.410 251.980 207.730 ;
        RECT 278.400 207.410 278.660 207.730 ;
        RECT 251.780 19.370 251.920 207.410 ;
        RECT 74.160 19.050 74.420 19.370 ;
        RECT 251.720 19.050 251.980 19.370 ;
        RECT 74.220 2.400 74.360 19.050 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 434.310 207.640 434.630 207.700 ;
        RECT 570.470 207.640 570.790 207.700 ;
        RECT 434.310 207.500 570.790 207.640 ;
        RECT 434.310 207.440 434.630 207.500 ;
        RECT 570.470 207.440 570.790 207.500 ;
        RECT 430.630 20.640 430.950 20.700 ;
        RECT 434.310 20.640 434.630 20.700 ;
        RECT 430.630 20.500 434.630 20.640 ;
        RECT 430.630 20.440 430.950 20.500 ;
        RECT 434.310 20.440 434.630 20.500 ;
      LAYER via ;
        RECT 434.340 207.440 434.600 207.700 ;
        RECT 570.500 207.440 570.760 207.700 ;
        RECT 430.660 20.440 430.920 20.700 ;
        RECT 434.340 20.440 434.600 20.700 ;
      LAYER met2 ;
        RECT 572.380 220.730 572.660 224.000 ;
        RECT 570.560 220.590 572.660 220.730 ;
        RECT 570.560 207.730 570.700 220.590 ;
        RECT 572.380 220.000 572.660 220.590 ;
        RECT 434.340 207.410 434.600 207.730 ;
        RECT 570.500 207.410 570.760 207.730 ;
        RECT 434.400 20.730 434.540 207.410 ;
        RECT 430.660 20.410 430.920 20.730 ;
        RECT 434.340 20.410 434.600 20.730 ;
        RECT 430.720 2.400 430.860 20.410 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 455.010 211.040 455.330 211.100 ;
        RECT 587.030 211.040 587.350 211.100 ;
        RECT 455.010 210.900 587.350 211.040 ;
        RECT 455.010 210.840 455.330 210.900 ;
        RECT 587.030 210.840 587.350 210.900 ;
        RECT 448.570 17.920 448.890 17.980 ;
        RECT 455.010 17.920 455.330 17.980 ;
        RECT 448.570 17.780 455.330 17.920 ;
        RECT 448.570 17.720 448.890 17.780 ;
        RECT 455.010 17.720 455.330 17.780 ;
      LAYER via ;
        RECT 455.040 210.840 455.300 211.100 ;
        RECT 587.060 210.840 587.320 211.100 ;
        RECT 448.600 17.720 448.860 17.980 ;
        RECT 455.040 17.720 455.300 17.980 ;
      LAYER met2 ;
        RECT 587.100 220.000 587.380 224.000 ;
        RECT 587.120 211.130 587.260 220.000 ;
        RECT 455.040 210.810 455.300 211.130 ;
        RECT 587.060 210.810 587.320 211.130 ;
        RECT 455.100 18.010 455.240 210.810 ;
        RECT 448.600 17.690 448.860 18.010 ;
        RECT 455.040 17.690 455.300 18.010 ;
        RECT 448.660 2.400 448.800 17.690 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 468.810 211.380 469.130 211.440 ;
        RECT 601.750 211.380 602.070 211.440 ;
        RECT 468.810 211.240 602.070 211.380 ;
        RECT 468.810 211.180 469.130 211.240 ;
        RECT 601.750 211.180 602.070 211.240 ;
        RECT 466.510 20.640 466.830 20.700 ;
        RECT 468.810 20.640 469.130 20.700 ;
        RECT 466.510 20.500 469.130 20.640 ;
        RECT 466.510 20.440 466.830 20.500 ;
        RECT 468.810 20.440 469.130 20.500 ;
      LAYER via ;
        RECT 468.840 211.180 469.100 211.440 ;
        RECT 601.780 211.180 602.040 211.440 ;
        RECT 466.540 20.440 466.800 20.700 ;
        RECT 468.840 20.440 469.100 20.700 ;
      LAYER met2 ;
        RECT 601.820 220.000 602.100 224.000 ;
        RECT 601.840 211.470 601.980 220.000 ;
        RECT 468.840 211.150 469.100 211.470 ;
        RECT 601.780 211.150 602.040 211.470 ;
        RECT 468.900 20.730 469.040 211.150 ;
        RECT 466.540 20.410 466.800 20.730 ;
        RECT 468.840 20.410 469.100 20.730 ;
        RECT 466.600 2.400 466.740 20.410 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 489.510 211.720 489.830 211.780 ;
        RECT 616.470 211.720 616.790 211.780 ;
        RECT 489.510 211.580 616.790 211.720 ;
        RECT 489.510 211.520 489.830 211.580 ;
        RECT 616.470 211.520 616.790 211.580 ;
        RECT 484.450 20.640 484.770 20.700 ;
        RECT 489.510 20.640 489.830 20.700 ;
        RECT 484.450 20.500 489.830 20.640 ;
        RECT 484.450 20.440 484.770 20.500 ;
        RECT 489.510 20.440 489.830 20.500 ;
      LAYER via ;
        RECT 489.540 211.520 489.800 211.780 ;
        RECT 616.500 211.520 616.760 211.780 ;
        RECT 484.480 20.440 484.740 20.700 ;
        RECT 489.540 20.440 489.800 20.700 ;
      LAYER met2 ;
        RECT 616.540 220.000 616.820 224.000 ;
        RECT 616.560 211.810 616.700 220.000 ;
        RECT 489.540 211.490 489.800 211.810 ;
        RECT 616.500 211.490 616.760 211.810 ;
        RECT 489.600 20.730 489.740 211.490 ;
        RECT 484.480 20.410 484.740 20.730 ;
        RECT 489.540 20.410 489.800 20.730 ;
        RECT 484.540 2.400 484.680 20.410 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 502.465 2.805 502.635 48.195 ;
      LAYER mcon ;
        RECT 502.465 48.025 502.635 48.195 ;
      LAYER met1 ;
        RECT 503.310 97.620 503.630 97.880 ;
        RECT 503.400 97.200 503.540 97.620 ;
        RECT 503.310 96.940 503.630 97.200 ;
        RECT 502.405 48.180 502.695 48.225 ;
        RECT 503.310 48.180 503.630 48.240 ;
        RECT 502.405 48.040 503.630 48.180 ;
        RECT 502.405 47.995 502.695 48.040 ;
        RECT 503.310 47.980 503.630 48.040 ;
        RECT 502.390 2.960 502.710 3.020 ;
        RECT 502.195 2.820 502.710 2.960 ;
        RECT 502.390 2.760 502.710 2.820 ;
      LAYER via ;
        RECT 503.340 97.620 503.600 97.880 ;
        RECT 503.340 96.940 503.600 97.200 ;
        RECT 503.340 47.980 503.600 48.240 ;
        RECT 502.420 2.760 502.680 3.020 ;
      LAYER met2 ;
        RECT 631.260 220.000 631.540 224.000 ;
        RECT 631.280 210.645 631.420 220.000 ;
        RECT 503.330 210.275 503.610 210.645 ;
        RECT 631.210 210.275 631.490 210.645 ;
        RECT 503.400 97.910 503.540 210.275 ;
        RECT 503.340 97.590 503.600 97.910 ;
        RECT 503.340 96.910 503.600 97.230 ;
        RECT 503.400 48.270 503.540 96.910 ;
        RECT 503.340 47.950 503.600 48.270 ;
        RECT 502.420 2.730 502.680 3.050 ;
        RECT 502.480 2.400 502.620 2.730 ;
        RECT 502.270 -4.800 502.830 2.400 ;
      LAYER via2 ;
        RECT 503.330 210.320 503.610 210.600 ;
        RECT 631.210 210.320 631.490 210.600 ;
      LAYER met3 ;
        RECT 503.305 210.610 503.635 210.625 ;
        RECT 631.185 210.610 631.515 210.625 ;
        RECT 503.305 210.310 631.515 210.610 ;
        RECT 503.305 210.295 503.635 210.310 ;
        RECT 631.185 210.295 631.515 210.310 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 524.010 209.680 524.330 209.740 ;
        RECT 645.910 209.680 646.230 209.740 ;
        RECT 524.010 209.540 646.230 209.680 ;
        RECT 524.010 209.480 524.330 209.540 ;
        RECT 645.910 209.480 646.230 209.540 ;
        RECT 519.870 15.880 520.190 15.940 ;
        RECT 524.010 15.880 524.330 15.940 ;
        RECT 519.870 15.740 524.330 15.880 ;
        RECT 519.870 15.680 520.190 15.740 ;
        RECT 524.010 15.680 524.330 15.740 ;
      LAYER via ;
        RECT 524.040 209.480 524.300 209.740 ;
        RECT 645.940 209.480 646.200 209.740 ;
        RECT 519.900 15.680 520.160 15.940 ;
        RECT 524.040 15.680 524.300 15.940 ;
      LAYER met2 ;
        RECT 645.980 220.000 646.260 224.000 ;
        RECT 646.000 209.770 646.140 220.000 ;
        RECT 524.040 209.450 524.300 209.770 ;
        RECT 645.940 209.450 646.200 209.770 ;
        RECT 524.100 15.970 524.240 209.450 ;
        RECT 519.900 15.650 520.160 15.970 ;
        RECT 524.040 15.650 524.300 15.970 ;
        RECT 519.960 2.400 520.100 15.650 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 646.920 214.300 648.440 214.440 ;
        RECT 537.810 213.760 538.130 213.820 ;
        RECT 646.920 213.760 647.060 214.300 ;
        RECT 537.810 213.620 647.060 213.760 ;
        RECT 648.300 213.760 648.440 214.300 ;
        RECT 656.030 213.760 656.350 213.820 ;
        RECT 648.300 213.620 656.350 213.760 ;
        RECT 537.810 213.560 538.130 213.620 ;
        RECT 656.030 213.560 656.350 213.620 ;
      LAYER via ;
        RECT 537.840 213.560 538.100 213.820 ;
        RECT 656.060 213.560 656.320 213.820 ;
      LAYER met2 ;
        RECT 660.700 220.730 660.980 224.000 ;
        RECT 656.120 220.590 660.980 220.730 ;
        RECT 656.120 213.850 656.260 220.590 ;
        RECT 660.700 220.000 660.980 220.590 ;
        RECT 537.840 213.530 538.100 213.850 ;
        RECT 656.060 213.530 656.320 213.850 ;
        RECT 537.900 2.400 538.040 213.530 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 638.165 208.165 638.335 209.355 ;
      LAYER mcon ;
        RECT 638.165 209.185 638.335 209.355 ;
      LAYER met1 ;
        RECT 638.105 209.340 638.395 209.385 ;
        RECT 675.350 209.340 675.670 209.400 ;
        RECT 638.105 209.200 675.670 209.340 ;
        RECT 638.105 209.155 638.395 209.200 ;
        RECT 675.350 209.140 675.670 209.200 ;
        RECT 558.510 208.320 558.830 208.380 ;
        RECT 638.105 208.320 638.395 208.365 ;
        RECT 558.510 208.180 638.395 208.320 ;
        RECT 558.510 208.120 558.830 208.180 ;
        RECT 638.105 208.135 638.395 208.180 ;
        RECT 555.750 20.640 556.070 20.700 ;
        RECT 558.510 20.640 558.830 20.700 ;
        RECT 555.750 20.500 558.830 20.640 ;
        RECT 555.750 20.440 556.070 20.500 ;
        RECT 558.510 20.440 558.830 20.500 ;
      LAYER via ;
        RECT 675.380 209.140 675.640 209.400 ;
        RECT 558.540 208.120 558.800 208.380 ;
        RECT 555.780 20.440 556.040 20.700 ;
        RECT 558.540 20.440 558.800 20.700 ;
      LAYER met2 ;
        RECT 675.420 220.000 675.700 224.000 ;
        RECT 675.440 209.430 675.580 220.000 ;
        RECT 675.380 209.110 675.640 209.430 ;
        RECT 558.540 208.090 558.800 208.410 ;
        RECT 558.600 20.730 558.740 208.090 ;
        RECT 555.780 20.410 556.040 20.730 ;
        RECT 558.540 20.410 558.800 20.730 ;
        RECT 555.840 2.400 555.980 20.410 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 579.210 208.660 579.530 208.720 ;
        RECT 690.070 208.660 690.390 208.720 ;
        RECT 579.210 208.520 690.390 208.660 ;
        RECT 579.210 208.460 579.530 208.520 ;
        RECT 690.070 208.460 690.390 208.520 ;
        RECT 573.690 17.580 574.010 17.640 ;
        RECT 579.210 17.580 579.530 17.640 ;
        RECT 573.690 17.440 579.530 17.580 ;
        RECT 573.690 17.380 574.010 17.440 ;
        RECT 579.210 17.380 579.530 17.440 ;
      LAYER via ;
        RECT 579.240 208.460 579.500 208.720 ;
        RECT 690.100 208.460 690.360 208.720 ;
        RECT 573.720 17.380 573.980 17.640 ;
        RECT 579.240 17.380 579.500 17.640 ;
      LAYER met2 ;
        RECT 690.140 220.000 690.420 224.000 ;
        RECT 690.160 208.750 690.300 220.000 ;
        RECT 579.240 208.430 579.500 208.750 ;
        RECT 690.100 208.430 690.360 208.750 ;
        RECT 579.300 17.670 579.440 208.430 ;
        RECT 573.720 17.350 573.980 17.670 ;
        RECT 579.240 17.350 579.500 17.670 ;
        RECT 573.780 2.400 573.920 17.350 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 626.665 210.545 628.215 210.715 ;
      LAYER mcon ;
        RECT 628.045 210.545 628.215 210.715 ;
      LAYER met1 ;
        RECT 593.010 210.700 593.330 210.760 ;
        RECT 626.605 210.700 626.895 210.745 ;
        RECT 593.010 210.560 626.895 210.700 ;
        RECT 593.010 210.500 593.330 210.560 ;
        RECT 626.605 210.515 626.895 210.560 ;
        RECT 627.985 210.700 628.275 210.745 ;
        RECT 704.790 210.700 705.110 210.760 ;
        RECT 627.985 210.560 705.110 210.700 ;
        RECT 627.985 210.515 628.275 210.560 ;
        RECT 704.790 210.500 705.110 210.560 ;
        RECT 591.170 14.180 591.490 14.240 ;
        RECT 593.010 14.180 593.330 14.240 ;
        RECT 591.170 14.040 593.330 14.180 ;
        RECT 591.170 13.980 591.490 14.040 ;
        RECT 593.010 13.980 593.330 14.040 ;
      LAYER via ;
        RECT 593.040 210.500 593.300 210.760 ;
        RECT 704.820 210.500 705.080 210.760 ;
        RECT 591.200 13.980 591.460 14.240 ;
        RECT 593.040 13.980 593.300 14.240 ;
      LAYER met2 ;
        RECT 704.860 220.000 705.140 224.000 ;
        RECT 704.880 210.790 705.020 220.000 ;
        RECT 593.040 210.470 593.300 210.790 ;
        RECT 704.820 210.470 705.080 210.790 ;
        RECT 593.100 14.270 593.240 210.470 ;
        RECT 591.200 13.950 591.460 14.270 ;
        RECT 593.040 13.950 593.300 14.270 ;
        RECT 591.260 2.400 591.400 13.950 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 103.110 212.740 103.430 212.800 ;
        RECT 298.150 212.740 298.470 212.800 ;
        RECT 103.110 212.600 298.470 212.740 ;
        RECT 103.110 212.540 103.430 212.600 ;
        RECT 298.150 212.540 298.470 212.600 ;
        RECT 97.590 20.640 97.910 20.700 ;
        RECT 103.110 20.640 103.430 20.700 ;
        RECT 97.590 20.500 103.430 20.640 ;
        RECT 97.590 20.440 97.910 20.500 ;
        RECT 103.110 20.440 103.430 20.500 ;
      LAYER via ;
        RECT 103.140 212.540 103.400 212.800 ;
        RECT 298.180 212.540 298.440 212.800 ;
        RECT 97.620 20.440 97.880 20.700 ;
        RECT 103.140 20.440 103.400 20.700 ;
      LAYER met2 ;
        RECT 298.220 220.000 298.500 224.000 ;
        RECT 298.240 212.830 298.380 220.000 ;
        RECT 103.140 212.510 103.400 212.830 ;
        RECT 298.180 212.510 298.440 212.830 ;
        RECT 103.200 20.730 103.340 212.510 ;
        RECT 97.620 20.410 97.880 20.730 ;
        RECT 103.140 20.410 103.400 20.730 ;
        RECT 97.680 2.400 97.820 20.410 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 613.710 211.380 614.030 211.440 ;
        RECT 719.050 211.380 719.370 211.440 ;
        RECT 613.710 211.240 719.370 211.380 ;
        RECT 613.710 211.180 614.030 211.240 ;
        RECT 719.050 211.180 719.370 211.240 ;
        RECT 609.110 18.600 609.430 18.660 ;
        RECT 613.710 18.600 614.030 18.660 ;
        RECT 609.110 18.460 614.030 18.600 ;
        RECT 609.110 18.400 609.430 18.460 ;
        RECT 613.710 18.400 614.030 18.460 ;
      LAYER via ;
        RECT 613.740 211.180 614.000 211.440 ;
        RECT 719.080 211.180 719.340 211.440 ;
        RECT 609.140 18.400 609.400 18.660 ;
        RECT 613.740 18.400 614.000 18.660 ;
      LAYER met2 ;
        RECT 719.120 220.000 719.400 224.000 ;
        RECT 719.140 211.470 719.280 220.000 ;
        RECT 613.740 211.150 614.000 211.470 ;
        RECT 719.080 211.150 719.340 211.470 ;
        RECT 613.800 18.690 613.940 211.150 ;
        RECT 609.140 18.370 609.400 18.690 ;
        RECT 613.740 18.370 614.000 18.690 ;
        RECT 609.200 2.400 609.340 18.370 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 628.430 211.040 628.750 211.100 ;
        RECT 733.770 211.040 734.090 211.100 ;
        RECT 628.430 210.900 734.090 211.040 ;
        RECT 628.430 210.840 628.750 210.900 ;
        RECT 733.770 210.840 734.090 210.900 ;
        RECT 626.590 62.120 626.910 62.180 ;
        RECT 627.510 62.120 627.830 62.180 ;
        RECT 626.590 61.980 627.830 62.120 ;
        RECT 626.590 61.920 626.910 61.980 ;
        RECT 627.510 61.920 627.830 61.980 ;
      LAYER via ;
        RECT 628.460 210.840 628.720 211.100 ;
        RECT 733.800 210.840 734.060 211.100 ;
        RECT 626.620 61.920 626.880 62.180 ;
        RECT 627.540 61.920 627.800 62.180 ;
      LAYER met2 ;
        RECT 733.840 220.000 734.120 224.000 ;
        RECT 733.860 211.130 734.000 220.000 ;
        RECT 628.460 210.810 628.720 211.130 ;
        RECT 733.800 210.810 734.060 211.130 ;
        RECT 628.520 210.530 628.660 210.810 ;
        RECT 627.600 210.390 628.660 210.530 ;
        RECT 627.600 62.210 627.740 210.390 ;
        RECT 626.620 61.890 626.880 62.210 ;
        RECT 627.540 61.890 627.800 62.210 ;
        RECT 626.680 15.370 626.820 61.890 ;
        RECT 626.680 15.230 627.280 15.370 ;
        RECT 627.140 2.400 627.280 15.230 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 299.990 207.300 300.310 207.360 ;
        RECT 317.470 207.300 317.790 207.360 ;
        RECT 299.990 207.160 317.790 207.300 ;
        RECT 299.990 207.100 300.310 207.160 ;
        RECT 317.470 207.100 317.790 207.160 ;
        RECT 121.510 19.620 121.830 19.680 ;
        RECT 299.530 19.620 299.850 19.680 ;
        RECT 121.510 19.480 299.850 19.620 ;
        RECT 121.510 19.420 121.830 19.480 ;
        RECT 299.530 19.420 299.850 19.480 ;
      LAYER via ;
        RECT 300.020 207.100 300.280 207.360 ;
        RECT 317.500 207.100 317.760 207.360 ;
        RECT 121.540 19.420 121.800 19.680 ;
        RECT 299.560 19.420 299.820 19.680 ;
      LAYER met2 ;
        RECT 317.540 220.000 317.820 224.000 ;
        RECT 317.560 207.390 317.700 220.000 ;
        RECT 300.020 207.070 300.280 207.390 ;
        RECT 317.500 207.070 317.760 207.390 ;
        RECT 300.080 21.490 300.220 207.070 ;
        RECT 299.620 21.350 300.220 21.490 ;
        RECT 299.620 19.710 299.760 21.350 ;
        RECT 121.540 19.390 121.800 19.710 ;
        RECT 299.560 19.390 299.820 19.710 ;
        RECT 121.600 2.400 121.740 19.390 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 303.285 213.095 303.455 213.775 ;
        RECT 299.605 207.145 299.775 213.095 ;
        RECT 302.825 212.925 303.455 213.095 ;
      LAYER mcon ;
        RECT 303.285 213.605 303.455 213.775 ;
        RECT 299.605 212.925 299.775 213.095 ;
      LAYER met1 ;
        RECT 303.225 213.760 303.515 213.805 ;
        RECT 337.250 213.760 337.570 213.820 ;
        RECT 303.225 213.620 337.570 213.760 ;
        RECT 303.225 213.575 303.515 213.620 ;
        RECT 337.250 213.560 337.570 213.620 ;
        RECT 299.545 213.080 299.835 213.125 ;
        RECT 302.765 213.080 303.055 213.125 ;
        RECT 299.545 212.940 303.055 213.080 ;
        RECT 299.545 212.895 299.835 212.940 ;
        RECT 302.765 212.895 303.055 212.940 ;
        RECT 196.490 207.300 196.810 207.360 ;
        RECT 299.545 207.300 299.835 207.345 ;
        RECT 196.490 207.160 299.835 207.300 ;
        RECT 196.490 207.100 196.810 207.160 ;
        RECT 299.545 207.115 299.835 207.160 ;
        RECT 145.430 20.300 145.750 20.360 ;
        RECT 196.490 20.300 196.810 20.360 ;
        RECT 145.430 20.160 196.810 20.300 ;
        RECT 145.430 20.100 145.750 20.160 ;
        RECT 196.490 20.100 196.810 20.160 ;
      LAYER via ;
        RECT 337.280 213.560 337.540 213.820 ;
        RECT 196.520 207.100 196.780 207.360 ;
        RECT 145.460 20.100 145.720 20.360 ;
        RECT 196.520 20.100 196.780 20.360 ;
      LAYER met2 ;
        RECT 337.320 220.000 337.600 224.000 ;
        RECT 337.340 213.850 337.480 220.000 ;
        RECT 337.280 213.530 337.540 213.850 ;
        RECT 196.520 207.070 196.780 207.390 ;
        RECT 196.580 20.390 196.720 207.070 ;
        RECT 145.460 20.070 145.720 20.390 ;
        RECT 196.520 20.070 196.780 20.390 ;
        RECT 145.520 2.400 145.660 20.070 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 163.370 18.600 163.690 18.660 ;
        RECT 351.970 18.600 352.290 18.660 ;
        RECT 163.370 18.460 352.290 18.600 ;
        RECT 163.370 18.400 163.690 18.460 ;
        RECT 351.970 18.400 352.290 18.460 ;
      LAYER via ;
        RECT 163.400 18.400 163.660 18.660 ;
        RECT 352.000 18.400 352.260 18.660 ;
      LAYER met2 ;
        RECT 352.040 220.000 352.320 224.000 ;
        RECT 352.060 18.690 352.200 220.000 ;
        RECT 163.400 18.370 163.660 18.690 ;
        RECT 352.000 18.370 352.260 18.690 ;
        RECT 163.460 2.400 163.600 18.370 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 341.390 207.980 341.710 208.040 ;
        RECT 366.690 207.980 367.010 208.040 ;
        RECT 341.390 207.840 367.010 207.980 ;
        RECT 341.390 207.780 341.710 207.840 ;
        RECT 366.690 207.780 367.010 207.840 ;
        RECT 180.850 20.640 181.170 20.700 ;
        RECT 180.850 20.500 197.180 20.640 ;
        RECT 180.850 20.440 181.170 20.500 ;
        RECT 197.040 20.300 197.180 20.500 ;
        RECT 341.390 20.300 341.710 20.360 ;
        RECT 197.040 20.160 341.710 20.300 ;
        RECT 341.390 20.100 341.710 20.160 ;
      LAYER via ;
        RECT 341.420 207.780 341.680 208.040 ;
        RECT 366.720 207.780 366.980 208.040 ;
        RECT 180.880 20.440 181.140 20.700 ;
        RECT 341.420 20.100 341.680 20.360 ;
      LAYER met2 ;
        RECT 366.760 220.000 367.040 224.000 ;
        RECT 366.780 208.070 366.920 220.000 ;
        RECT 341.420 207.750 341.680 208.070 ;
        RECT 366.720 207.750 366.980 208.070 ;
        RECT 180.880 20.410 181.140 20.730 ;
        RECT 180.940 2.400 181.080 20.410 ;
        RECT 341.480 20.390 341.620 207.750 ;
        RECT 341.420 20.070 341.680 20.390 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 198.790 18.940 199.110 19.000 ;
        RECT 380.490 18.940 380.810 19.000 ;
        RECT 198.790 18.800 380.810 18.940 ;
        RECT 198.790 18.740 199.110 18.800 ;
        RECT 380.490 18.740 380.810 18.800 ;
      LAYER via ;
        RECT 198.820 18.740 199.080 19.000 ;
        RECT 380.520 18.740 380.780 19.000 ;
      LAYER met2 ;
        RECT 381.480 220.730 381.760 224.000 ;
        RECT 380.580 220.590 381.760 220.730 ;
        RECT 380.580 19.030 380.720 220.590 ;
        RECT 381.480 220.000 381.760 220.590 ;
        RECT 198.820 18.710 199.080 19.030 ;
        RECT 380.520 18.710 380.780 19.030 ;
        RECT 198.880 2.400 199.020 18.710 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 216.730 17.580 217.050 17.640 ;
        RECT 220.410 17.580 220.730 17.640 ;
        RECT 216.730 17.440 220.730 17.580 ;
        RECT 216.730 17.380 217.050 17.440 ;
        RECT 220.410 17.380 220.730 17.440 ;
      LAYER via ;
        RECT 216.760 17.380 217.020 17.640 ;
        RECT 220.440 17.380 220.700 17.640 ;
      LAYER met2 ;
        RECT 396.200 220.000 396.480 224.000 ;
        RECT 396.220 210.645 396.360 220.000 ;
        RECT 220.430 210.275 220.710 210.645 ;
        RECT 396.150 210.275 396.430 210.645 ;
        RECT 220.500 17.670 220.640 210.275 ;
        RECT 216.760 17.350 217.020 17.670 ;
        RECT 220.440 17.350 220.700 17.670 ;
        RECT 216.820 2.400 216.960 17.350 ;
        RECT 216.610 -4.800 217.170 2.400 ;
      LAYER via2 ;
        RECT 220.430 210.320 220.710 210.600 ;
        RECT 396.150 210.320 396.430 210.600 ;
      LAYER met3 ;
        RECT 220.405 210.610 220.735 210.625 ;
        RECT 396.125 210.610 396.455 210.625 ;
        RECT 220.405 210.310 396.455 210.610 ;
        RECT 220.405 210.295 220.735 210.310 ;
        RECT 396.125 210.295 396.455 210.310 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 375.965 17.765 376.135 20.655 ;
      LAYER mcon ;
        RECT 375.965 20.485 376.135 20.655 ;
      LAYER met1 ;
        RECT 403.490 207.640 403.810 207.700 ;
        RECT 410.850 207.640 411.170 207.700 ;
        RECT 403.490 207.500 411.170 207.640 ;
        RECT 403.490 207.440 403.810 207.500 ;
        RECT 410.850 207.440 411.170 207.500 ;
        RECT 375.905 20.640 376.195 20.685 ;
        RECT 403.490 20.640 403.810 20.700 ;
        RECT 375.905 20.500 403.810 20.640 ;
        RECT 375.905 20.455 376.195 20.500 ;
        RECT 403.490 20.440 403.810 20.500 ;
        RECT 234.670 17.920 234.990 17.980 ;
        RECT 375.905 17.920 376.195 17.965 ;
        RECT 234.670 17.780 376.195 17.920 ;
        RECT 234.670 17.720 234.990 17.780 ;
        RECT 375.905 17.735 376.195 17.780 ;
      LAYER via ;
        RECT 403.520 207.440 403.780 207.700 ;
        RECT 410.880 207.440 411.140 207.700 ;
        RECT 403.520 20.440 403.780 20.700 ;
        RECT 234.700 17.720 234.960 17.980 ;
      LAYER met2 ;
        RECT 410.920 220.000 411.200 224.000 ;
        RECT 410.940 207.730 411.080 220.000 ;
        RECT 403.520 207.410 403.780 207.730 ;
        RECT 410.880 207.410 411.140 207.730 ;
        RECT 403.580 20.730 403.720 207.410 ;
        RECT 403.520 20.410 403.780 20.730 ;
        RECT 234.700 17.690 234.960 18.010 ;
        RECT 234.760 2.400 234.900 17.690 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 61.710 211.380 62.030 211.440 ;
        RECT 263.650 211.380 263.970 211.440 ;
        RECT 61.710 211.240 263.970 211.380 ;
        RECT 61.710 211.180 62.030 211.240 ;
        RECT 263.650 211.180 263.970 211.240 ;
        RECT 56.190 16.900 56.510 16.960 ;
        RECT 61.710 16.900 62.030 16.960 ;
        RECT 56.190 16.760 62.030 16.900 ;
        RECT 56.190 16.700 56.510 16.760 ;
        RECT 61.710 16.700 62.030 16.760 ;
      LAYER via ;
        RECT 61.740 211.180 62.000 211.440 ;
        RECT 263.680 211.180 263.940 211.440 ;
        RECT 56.220 16.700 56.480 16.960 ;
        RECT 61.740 16.700 62.000 16.960 ;
      LAYER met2 ;
        RECT 263.720 220.000 264.000 224.000 ;
        RECT 263.740 211.470 263.880 220.000 ;
        RECT 61.740 211.150 62.000 211.470 ;
        RECT 263.680 211.150 263.940 211.470 ;
        RECT 61.800 16.990 61.940 211.150 ;
        RECT 56.220 16.670 56.480 16.990 ;
        RECT 61.740 16.670 62.000 16.990 ;
        RECT 56.280 2.400 56.420 16.670 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 82.410 211.720 82.730 211.780 ;
        RECT 283.430 211.720 283.750 211.780 ;
        RECT 82.410 211.580 283.750 211.720 ;
        RECT 82.410 211.520 82.730 211.580 ;
        RECT 283.430 211.520 283.750 211.580 ;
        RECT 80.110 20.640 80.430 20.700 ;
        RECT 82.410 20.640 82.730 20.700 ;
        RECT 80.110 20.500 82.730 20.640 ;
        RECT 80.110 20.440 80.430 20.500 ;
        RECT 82.410 20.440 82.730 20.500 ;
      LAYER via ;
        RECT 82.440 211.520 82.700 211.780 ;
        RECT 283.460 211.520 283.720 211.780 ;
        RECT 80.140 20.440 80.400 20.700 ;
        RECT 82.440 20.440 82.700 20.700 ;
      LAYER met2 ;
        RECT 283.500 220.000 283.780 224.000 ;
        RECT 283.520 211.810 283.660 220.000 ;
        RECT 82.440 211.490 82.700 211.810 ;
        RECT 283.460 211.490 283.720 211.810 ;
        RECT 82.500 20.730 82.640 211.490 ;
        RECT 80.140 20.410 80.400 20.730 ;
        RECT 82.440 20.410 82.700 20.730 ;
        RECT 80.200 2.400 80.340 20.410 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 213.760 109.870 213.820 ;
        RECT 302.750 213.760 303.070 213.820 ;
        RECT 109.550 213.620 303.070 213.760 ;
        RECT 109.550 213.560 109.870 213.620 ;
        RECT 302.750 213.560 303.070 213.620 ;
        RECT 103.570 20.640 103.890 20.700 ;
        RECT 109.550 20.640 109.870 20.700 ;
        RECT 103.570 20.500 109.870 20.640 ;
        RECT 103.570 20.440 103.890 20.500 ;
        RECT 109.550 20.440 109.870 20.500 ;
      LAYER via ;
        RECT 109.580 213.560 109.840 213.820 ;
        RECT 302.780 213.560 303.040 213.820 ;
        RECT 103.600 20.440 103.860 20.700 ;
        RECT 109.580 20.440 109.840 20.700 ;
      LAYER met2 ;
        RECT 302.820 220.000 303.100 224.000 ;
        RECT 302.840 213.850 302.980 220.000 ;
        RECT 109.580 213.530 109.840 213.850 ;
        RECT 302.780 213.530 303.040 213.850 ;
        RECT 109.640 20.730 109.780 213.530 ;
        RECT 103.600 20.410 103.860 20.730 ;
        RECT 109.580 20.410 109.840 20.730 ;
        RECT 103.660 2.400 103.800 20.410 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 286.190 207.640 286.510 207.700 ;
        RECT 322.530 207.640 322.850 207.700 ;
        RECT 286.190 207.500 322.850 207.640 ;
        RECT 286.190 207.440 286.510 207.500 ;
        RECT 322.530 207.440 322.850 207.500 ;
        RECT 127.490 19.960 127.810 20.020 ;
        RECT 286.190 19.960 286.510 20.020 ;
        RECT 127.490 19.820 286.510 19.960 ;
        RECT 127.490 19.760 127.810 19.820 ;
        RECT 286.190 19.760 286.510 19.820 ;
      LAYER via ;
        RECT 286.220 207.440 286.480 207.700 ;
        RECT 322.560 207.440 322.820 207.700 ;
        RECT 127.520 19.760 127.780 20.020 ;
        RECT 286.220 19.760 286.480 20.020 ;
      LAYER met2 ;
        RECT 322.600 220.000 322.880 224.000 ;
        RECT 322.620 207.730 322.760 220.000 ;
        RECT 286.220 207.410 286.480 207.730 ;
        RECT 322.560 207.410 322.820 207.730 ;
        RECT 286.280 20.050 286.420 207.410 ;
        RECT 127.520 19.730 127.780 20.050 ;
        RECT 286.220 19.730 286.480 20.050 ;
        RECT 127.580 2.400 127.720 19.730 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 27.210 210.360 27.530 210.420 ;
        RECT 239.270 210.360 239.590 210.420 ;
        RECT 27.210 210.220 239.590 210.360 ;
        RECT 27.210 210.160 27.530 210.220 ;
        RECT 239.270 210.160 239.590 210.220 ;
      LAYER via ;
        RECT 27.240 210.160 27.500 210.420 ;
        RECT 239.300 210.160 239.560 210.420 ;
      LAYER met2 ;
        RECT 239.340 220.000 239.620 224.000 ;
        RECT 239.360 210.450 239.500 220.000 ;
        RECT 27.240 210.130 27.500 210.450 ;
        RECT 239.300 210.130 239.560 210.450 ;
        RECT 27.300 24.210 27.440 210.130 ;
        RECT 26.380 24.070 27.440 24.210 ;
        RECT 26.380 2.400 26.520 24.070 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 203.005 17.425 203.175 18.275 ;
      LAYER mcon ;
        RECT 203.005 18.105 203.175 18.275 ;
      LAYER met1 ;
        RECT 230.990 207.640 231.310 207.700 ;
        RECT 244.330 207.640 244.650 207.700 ;
        RECT 230.990 207.500 244.650 207.640 ;
        RECT 230.990 207.440 231.310 207.500 ;
        RECT 244.330 207.440 244.650 207.500 ;
        RECT 82.500 18.800 135.080 18.940 ;
        RECT 32.270 18.260 32.590 18.320 ;
        RECT 82.500 18.260 82.640 18.800 ;
        RECT 32.270 18.120 82.640 18.260 ;
        RECT 134.940 18.260 135.080 18.800 ;
        RECT 202.945 18.260 203.235 18.305 ;
        RECT 134.940 18.120 203.235 18.260 ;
        RECT 32.270 18.060 32.590 18.120 ;
        RECT 202.945 18.075 203.235 18.120 ;
        RECT 230.990 17.920 231.310 17.980 ;
        RECT 203.940 17.780 231.310 17.920 ;
        RECT 202.945 17.580 203.235 17.625 ;
        RECT 203.940 17.580 204.080 17.780 ;
        RECT 230.990 17.720 231.310 17.780 ;
        RECT 202.945 17.440 204.080 17.580 ;
        RECT 202.945 17.395 203.235 17.440 ;
      LAYER via ;
        RECT 231.020 207.440 231.280 207.700 ;
        RECT 244.360 207.440 244.620 207.700 ;
        RECT 32.300 18.060 32.560 18.320 ;
        RECT 231.020 17.720 231.280 17.980 ;
      LAYER met2 ;
        RECT 244.400 220.000 244.680 224.000 ;
        RECT 244.420 207.730 244.560 220.000 ;
        RECT 231.020 207.410 231.280 207.730 ;
        RECT 244.360 207.410 244.620 207.730 ;
        RECT 32.300 18.030 32.560 18.350 ;
        RECT 32.360 2.400 32.500 18.030 ;
        RECT 231.080 18.010 231.220 207.410 ;
        RECT 231.020 17.690 231.280 18.010 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 -9.220 367.020 3528.900 ;
        RECT 544.020 -9.220 547.020 3528.900 ;
        RECT 724.020 -9.220 727.020 3528.900 ;
        RECT 904.020 -9.220 907.020 3528.900 ;
        RECT 1084.020 -9.220 1087.020 3528.900 ;
        RECT 1264.020 -9.220 1267.020 3528.900 ;
        RECT 1444.020 -9.220 1447.020 3528.900 ;
        RECT 1624.020 -9.220 1627.020 3528.900 ;
        RECT 1804.020 -9.220 1807.020 3528.900 ;
        RECT 1984.020 -9.220 1987.020 3528.900 ;
        RECT 2164.020 -9.220 2167.020 3528.900 ;
        RECT 2344.020 -9.220 2347.020 3528.900 ;
        RECT 2524.020 -9.220 2527.020 3528.900 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 -9.220 457.020 3528.900 ;
        RECT 634.020 -9.220 637.020 3528.900 ;
        RECT 814.020 -9.220 817.020 3528.900 ;
        RECT 994.020 -9.220 997.020 3528.900 ;
        RECT 1174.020 -9.220 1177.020 3528.900 ;
        RECT 1354.020 -9.220 1357.020 3528.900 ;
        RECT 1534.020 -9.220 1537.020 3528.900 ;
        RECT 1714.020 -9.220 1717.020 3528.900 ;
        RECT 1894.020 -9.220 1897.020 3528.900 ;
        RECT 2074.020 -9.220 2077.020 3528.900 ;
        RECT 2254.020 -9.220 2257.020 3528.900 ;
        RECT 2434.020 -9.220 2437.020 3528.900 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 -18.420 385.020 3538.100 ;
        RECT 562.020 -18.420 565.020 3538.100 ;
        RECT 742.020 -18.420 745.020 3538.100 ;
        RECT 922.020 -18.420 925.020 3538.100 ;
        RECT 1102.020 -18.420 1105.020 3538.100 ;
        RECT 1282.020 -18.420 1285.020 3538.100 ;
        RECT 1462.020 -18.420 1465.020 3538.100 ;
        RECT 1642.020 -18.420 1645.020 3538.100 ;
        RECT 1822.020 -18.420 1825.020 3538.100 ;
        RECT 2002.020 -18.420 2005.020 3538.100 ;
        RECT 2182.020 -18.420 2185.020 3538.100 ;
        RECT 2362.020 -18.420 2365.020 3538.100 ;
        RECT 2542.020 -18.420 2545.020 3538.100 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1282.930 2009.090 1284.110 2010.270 ;
        RECT 1282.930 2007.490 1284.110 2008.670 ;
        RECT 1282.930 1829.090 1284.110 1830.270 ;
        RECT 1282.930 1827.490 1284.110 1828.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 1282.020 2010.380 1285.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 1282.020 2007.370 1285.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 1282.020 1830.380 1285.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 1282.020 1827.370 1285.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 -18.420 475.020 3538.100 ;
        RECT 652.020 -18.420 655.020 3538.100 ;
        RECT 832.020 -18.420 835.020 3538.100 ;
        RECT 1012.020 -18.420 1015.020 3538.100 ;
        RECT 1192.020 -18.420 1195.020 3538.100 ;
        RECT 1372.020 -18.420 1375.020 3538.100 ;
        RECT 1552.020 -18.420 1555.020 3538.100 ;
        RECT 1732.020 -18.420 1735.020 3538.100 ;
        RECT 1912.020 -18.420 1915.020 3538.100 ;
        RECT 2092.020 -18.420 2095.020 3538.100 ;
        RECT 2272.020 -18.420 2275.020 3538.100 ;
        RECT 2452.020 -18.420 2455.020 3538.100 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 -27.620 403.020 3547.300 ;
        RECT 580.020 -27.620 583.020 3547.300 ;
        RECT 760.020 -27.620 763.020 3547.300 ;
        RECT 940.020 -27.620 943.020 3547.300 ;
        RECT 1120.020 -27.620 1123.020 3547.300 ;
        RECT 1300.020 -27.620 1303.020 3547.300 ;
        RECT 1480.020 -27.620 1483.020 3547.300 ;
        RECT 1660.020 -27.620 1663.020 3547.300 ;
        RECT 1840.020 -27.620 1843.020 3547.300 ;
        RECT 2020.020 -27.620 2023.020 3547.300 ;
        RECT 2200.020 -27.620 2203.020 3547.300 ;
        RECT 2380.020 -27.620 2383.020 3547.300 ;
        RECT 2560.020 -27.620 2563.020 3547.300 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1300.930 2027.090 1302.110 2028.270 ;
        RECT 1300.930 2025.490 1302.110 2026.670 ;
        RECT 1300.930 1847.090 1302.110 1848.270 ;
        RECT 1300.930 1845.490 1302.110 1846.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 1300.020 2028.380 1303.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 1300.020 2025.370 1303.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 1300.020 1848.380 1303.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 1300.020 1845.370 1303.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 -27.620 313.020 3547.300 ;
        RECT 490.020 -27.620 493.020 3547.300 ;
        RECT 670.020 -27.620 673.020 3547.300 ;
        RECT 850.020 -27.620 853.020 3547.300 ;
        RECT 1030.020 -27.620 1033.020 3547.300 ;
        RECT 1210.020 -27.620 1213.020 3547.300 ;
        RECT 1390.020 -27.620 1393.020 3547.300 ;
        RECT 1570.020 -27.620 1573.020 3547.300 ;
        RECT 1750.020 -27.620 1753.020 3547.300 ;
        RECT 1930.020 -27.620 1933.020 3547.300 ;
        RECT 2110.020 -27.620 2113.020 3547.300 ;
        RECT 2290.020 -27.620 2293.020 3547.300 ;
        RECT 2470.020 -27.620 2473.020 3547.300 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 1930.930 1757.090 1932.110 1758.270 ;
        RECT 1930.930 1755.490 1932.110 1756.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 1930.020 1758.380 1933.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 1930.020 1755.370 1933.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 -36.820 421.020 3556.500 ;
        RECT 598.020 -36.820 601.020 3556.500 ;
        RECT 778.020 -36.820 781.020 3556.500 ;
        RECT 958.020 -36.820 961.020 3556.500 ;
        RECT 1138.020 -36.820 1141.020 3556.500 ;
        RECT 1318.020 -36.820 1321.020 3556.500 ;
        RECT 1498.020 -36.820 1501.020 3556.500 ;
        RECT 1678.020 -36.820 1681.020 3556.500 ;
        RECT 1858.020 -36.820 1861.020 3556.500 ;
        RECT 2038.020 -36.820 2041.020 3556.500 ;
        RECT 2218.020 -36.820 2221.020 3556.500 ;
        RECT 2398.020 -36.820 2401.020 3556.500 ;
        RECT 2578.020 -36.820 2581.020 3556.500 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1318.930 2045.090 1320.110 2046.270 ;
        RECT 1318.930 2043.490 1320.110 2044.670 ;
        RECT 1318.930 1865.090 1320.110 1866.270 ;
        RECT 1318.930 1863.490 1320.110 1864.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 1318.020 2046.380 1321.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 1318.020 2043.370 1321.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 1318.020 1866.380 1321.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 1318.020 1863.370 1321.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 -36.820 331.020 3556.500 ;
        RECT 508.020 -36.820 511.020 3556.500 ;
        RECT 688.020 -36.820 691.020 3556.500 ;
        RECT 868.020 -36.820 871.020 3556.500 ;
        RECT 1048.020 -36.820 1051.020 3556.500 ;
        RECT 1228.020 -36.820 1231.020 3556.500 ;
        RECT 1408.020 -36.820 1411.020 3556.500 ;
        RECT 1588.020 -36.820 1591.020 3556.500 ;
        RECT 1768.020 -36.820 1771.020 3556.500 ;
        RECT 1948.020 -36.820 1951.020 3556.500 ;
        RECT 2128.020 -36.820 2131.020 3556.500 ;
        RECT 2308.020 -36.820 2311.020 3556.500 ;
        RECT 2488.020 -36.820 2491.020 3556.500 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 1948.930 1775.090 1950.110 1776.270 ;
        RECT 1948.930 1773.490 1950.110 1774.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 1948.020 1776.380 1951.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 1948.020 1773.370 1951.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 223.150 230.795 2611.930 3206.645 ;
      LAYER met1 ;
        RECT 220.000 224.460 2611.930 3208.220 ;
      LAYER met2 ;
        RECT 220.030 3215.720 227.560 3216.000 ;
        RECT 228.400 3215.720 248.260 3216.000 ;
        RECT 249.100 3215.720 269.420 3216.000 ;
        RECT 270.260 3215.720 290.580 3216.000 ;
        RECT 291.420 3215.720 311.740 3216.000 ;
        RECT 312.580 3215.720 332.440 3216.000 ;
        RECT 333.280 3215.720 353.600 3216.000 ;
        RECT 354.440 3215.720 374.760 3216.000 ;
        RECT 375.600 3215.720 395.920 3216.000 ;
        RECT 396.760 3215.720 416.620 3216.000 ;
        RECT 417.460 3215.720 437.780 3216.000 ;
        RECT 438.620 3215.720 458.940 3216.000 ;
        RECT 459.780 3215.720 480.100 3216.000 ;
        RECT 480.940 3215.720 500.800 3216.000 ;
        RECT 501.640 3215.720 521.960 3216.000 ;
        RECT 522.800 3215.720 543.120 3216.000 ;
        RECT 543.960 3215.720 564.280 3216.000 ;
        RECT 565.120 3215.720 584.980 3216.000 ;
        RECT 585.820 3215.720 606.140 3216.000 ;
        RECT 606.980 3215.720 627.300 3216.000 ;
        RECT 628.140 3215.720 648.460 3216.000 ;
        RECT 649.300 3215.720 669.620 3216.000 ;
        RECT 670.460 3215.720 690.320 3216.000 ;
        RECT 691.160 3215.720 711.480 3216.000 ;
        RECT 712.320 3215.720 732.640 3216.000 ;
        RECT 733.480 3215.720 753.800 3216.000 ;
        RECT 754.640 3215.720 774.500 3216.000 ;
        RECT 775.340 3215.720 795.660 3216.000 ;
        RECT 796.500 3215.720 816.820 3216.000 ;
        RECT 817.660 3215.720 837.980 3216.000 ;
        RECT 838.820 3215.720 858.680 3216.000 ;
        RECT 859.520 3215.720 879.840 3216.000 ;
        RECT 880.680 3215.720 901.000 3216.000 ;
        RECT 901.840 3215.720 922.160 3216.000 ;
        RECT 923.000 3215.720 942.860 3216.000 ;
        RECT 943.700 3215.720 964.020 3216.000 ;
        RECT 964.860 3215.720 985.180 3216.000 ;
        RECT 986.020 3215.720 1006.340 3216.000 ;
        RECT 1007.180 3215.720 1027.500 3216.000 ;
        RECT 1028.340 3215.720 1048.200 3216.000 ;
        RECT 1049.040 3215.720 1069.360 3216.000 ;
        RECT 1070.200 3215.720 1090.520 3216.000 ;
        RECT 1091.360 3215.720 1111.680 3216.000 ;
        RECT 1112.520 3215.720 1132.380 3216.000 ;
        RECT 1133.220 3215.720 1153.540 3216.000 ;
        RECT 1154.380 3215.720 1174.700 3216.000 ;
        RECT 1175.540 3215.720 1195.860 3216.000 ;
        RECT 1196.700 3215.720 1216.560 3216.000 ;
        RECT 1217.400 3215.720 1237.720 3216.000 ;
        RECT 1238.560 3215.720 1258.880 3216.000 ;
        RECT 1259.720 3215.720 1280.040 3216.000 ;
        RECT 1280.880 3215.720 1300.740 3216.000 ;
        RECT 1301.580 3215.720 1321.900 3216.000 ;
        RECT 1322.740 3215.720 1343.060 3216.000 ;
        RECT 1343.900 3215.720 1364.220 3216.000 ;
        RECT 1365.060 3215.720 1384.920 3216.000 ;
        RECT 1385.760 3215.720 1406.080 3216.000 ;
        RECT 1406.920 3215.720 1427.240 3216.000 ;
        RECT 1428.080 3215.720 1448.400 3216.000 ;
        RECT 1449.240 3215.720 1469.560 3216.000 ;
        RECT 1470.400 3215.720 1490.260 3216.000 ;
        RECT 1491.100 3215.720 1511.420 3216.000 ;
        RECT 1512.260 3215.720 1532.580 3216.000 ;
        RECT 1533.420 3215.720 1553.740 3216.000 ;
        RECT 1554.580 3215.720 1574.440 3216.000 ;
        RECT 1575.280 3215.720 1595.600 3216.000 ;
        RECT 1596.440 3215.720 1616.760 3216.000 ;
        RECT 1617.600 3215.720 1637.920 3216.000 ;
        RECT 1638.760 3215.720 1658.620 3216.000 ;
        RECT 1659.460 3215.720 1679.780 3216.000 ;
        RECT 1680.620 3215.720 1700.940 3216.000 ;
        RECT 1701.780 3215.720 1722.100 3216.000 ;
        RECT 1722.940 3215.720 1742.800 3216.000 ;
        RECT 1743.640 3215.720 1763.960 3216.000 ;
        RECT 1764.800 3215.720 1785.120 3216.000 ;
        RECT 1785.960 3215.720 1806.280 3216.000 ;
        RECT 1807.120 3215.720 1827.440 3216.000 ;
        RECT 1828.280 3215.720 1848.140 3216.000 ;
        RECT 1848.980 3215.720 1869.300 3216.000 ;
        RECT 1870.140 3215.720 1890.460 3216.000 ;
        RECT 1891.300 3215.720 1911.620 3216.000 ;
        RECT 1912.460 3215.720 1932.320 3216.000 ;
        RECT 1933.160 3215.720 1953.480 3216.000 ;
        RECT 1954.320 3215.720 1974.640 3216.000 ;
        RECT 1975.480 3215.720 1995.800 3216.000 ;
        RECT 1996.640 3215.720 2016.500 3216.000 ;
        RECT 2017.340 3215.720 2037.660 3216.000 ;
        RECT 2038.500 3215.720 2058.820 3216.000 ;
        RECT 2059.660 3215.720 2079.980 3216.000 ;
        RECT 2080.820 3215.720 2100.680 3216.000 ;
        RECT 2101.520 3215.720 2121.840 3216.000 ;
        RECT 2122.680 3215.720 2143.000 3216.000 ;
        RECT 2143.840 3215.720 2164.160 3216.000 ;
        RECT 2165.000 3215.720 2184.860 3216.000 ;
        RECT 2185.700 3215.720 2206.020 3216.000 ;
        RECT 2206.860 3215.720 2227.180 3216.000 ;
        RECT 2228.020 3215.720 2248.340 3216.000 ;
        RECT 2249.180 3215.720 2269.500 3216.000 ;
        RECT 2270.340 3215.720 2290.200 3216.000 ;
        RECT 2291.040 3215.720 2311.360 3216.000 ;
        RECT 2312.200 3215.720 2332.520 3216.000 ;
        RECT 2333.360 3215.720 2353.680 3216.000 ;
        RECT 2354.520 3215.720 2374.380 3216.000 ;
        RECT 2375.220 3215.720 2395.540 3216.000 ;
        RECT 2396.380 3215.720 2416.700 3216.000 ;
        RECT 2417.540 3215.720 2437.860 3216.000 ;
        RECT 2438.700 3215.720 2458.560 3216.000 ;
        RECT 2459.400 3215.720 2479.720 3216.000 ;
        RECT 2480.560 3215.720 2500.880 3216.000 ;
        RECT 2501.720 3215.720 2522.040 3216.000 ;
        RECT 2522.880 3215.720 2542.740 3216.000 ;
        RECT 2543.580 3215.720 2563.900 3216.000 ;
        RECT 2564.740 3215.720 2585.060 3216.000 ;
        RECT 2585.900 3215.720 2606.220 3216.000 ;
        RECT 2607.060 3215.720 2609.990 3216.000 ;
        RECT 220.030 224.280 2609.990 3215.720 ;
        RECT 220.580 224.000 224.340 224.280 ;
        RECT 225.180 224.000 229.400 224.280 ;
        RECT 230.240 224.000 234.000 224.280 ;
        RECT 234.840 224.000 239.060 224.280 ;
        RECT 239.900 224.000 244.120 224.280 ;
        RECT 244.960 224.000 248.720 224.280 ;
        RECT 249.560 224.000 253.780 224.280 ;
        RECT 254.620 224.000 258.840 224.280 ;
        RECT 259.680 224.000 263.440 224.280 ;
        RECT 264.280 224.000 268.500 224.280 ;
        RECT 269.340 224.000 273.560 224.280 ;
        RECT 274.400 224.000 278.160 224.280 ;
        RECT 279.000 224.000 283.220 224.280 ;
        RECT 284.060 224.000 288.280 224.280 ;
        RECT 289.120 224.000 292.880 224.280 ;
        RECT 293.720 224.000 297.940 224.280 ;
        RECT 298.780 224.000 302.540 224.280 ;
        RECT 303.380 224.000 307.600 224.280 ;
        RECT 308.440 224.000 312.660 224.280 ;
        RECT 313.500 224.000 317.260 224.280 ;
        RECT 318.100 224.000 322.320 224.280 ;
        RECT 323.160 224.000 327.380 224.280 ;
        RECT 328.220 224.000 331.980 224.280 ;
        RECT 332.820 224.000 337.040 224.280 ;
        RECT 337.880 224.000 342.100 224.280 ;
        RECT 342.940 224.000 346.700 224.280 ;
        RECT 347.540 224.000 351.760 224.280 ;
        RECT 352.600 224.000 356.820 224.280 ;
        RECT 357.660 224.000 361.420 224.280 ;
        RECT 362.260 224.000 366.480 224.280 ;
        RECT 367.320 224.000 371.540 224.280 ;
        RECT 372.380 224.000 376.140 224.280 ;
        RECT 376.980 224.000 381.200 224.280 ;
        RECT 382.040 224.000 385.800 224.280 ;
        RECT 386.640 224.000 390.860 224.280 ;
        RECT 391.700 224.000 395.920 224.280 ;
        RECT 396.760 224.000 400.520 224.280 ;
        RECT 401.360 224.000 405.580 224.280 ;
        RECT 406.420 224.000 410.640 224.280 ;
        RECT 411.480 224.000 415.240 224.280 ;
        RECT 416.080 224.000 420.300 224.280 ;
        RECT 421.140 224.000 425.360 224.280 ;
        RECT 426.200 224.000 429.960 224.280 ;
        RECT 430.800 224.000 435.020 224.280 ;
        RECT 435.860 224.000 440.080 224.280 ;
        RECT 440.920 224.000 444.680 224.280 ;
        RECT 445.520 224.000 449.740 224.280 ;
        RECT 450.580 224.000 454.800 224.280 ;
        RECT 455.640 224.000 459.400 224.280 ;
        RECT 460.240 224.000 464.460 224.280 ;
        RECT 465.300 224.000 469.060 224.280 ;
        RECT 469.900 224.000 474.120 224.280 ;
        RECT 474.960 224.000 479.180 224.280 ;
        RECT 480.020 224.000 483.780 224.280 ;
        RECT 484.620 224.000 488.840 224.280 ;
        RECT 489.680 224.000 493.900 224.280 ;
        RECT 494.740 224.000 498.500 224.280 ;
        RECT 499.340 224.000 503.560 224.280 ;
        RECT 504.400 224.000 508.620 224.280 ;
        RECT 509.460 224.000 513.220 224.280 ;
        RECT 514.060 224.000 518.280 224.280 ;
        RECT 519.120 224.000 523.340 224.280 ;
        RECT 524.180 224.000 527.940 224.280 ;
        RECT 528.780 224.000 533.000 224.280 ;
        RECT 533.840 224.000 538.060 224.280 ;
        RECT 538.900 224.000 542.660 224.280 ;
        RECT 543.500 224.000 547.720 224.280 ;
        RECT 548.560 224.000 552.320 224.280 ;
        RECT 553.160 224.000 557.380 224.280 ;
        RECT 558.220 224.000 562.440 224.280 ;
        RECT 563.280 224.000 567.040 224.280 ;
        RECT 567.880 224.000 572.100 224.280 ;
        RECT 572.940 224.000 577.160 224.280 ;
        RECT 578.000 224.000 581.760 224.280 ;
        RECT 582.600 224.000 586.820 224.280 ;
        RECT 587.660 224.000 591.880 224.280 ;
        RECT 592.720 224.000 596.480 224.280 ;
        RECT 597.320 224.000 601.540 224.280 ;
        RECT 602.380 224.000 606.600 224.280 ;
        RECT 607.440 224.000 611.200 224.280 ;
        RECT 612.040 224.000 616.260 224.280 ;
        RECT 617.100 224.000 621.320 224.280 ;
        RECT 622.160 224.000 625.920 224.280 ;
        RECT 626.760 224.000 630.980 224.280 ;
        RECT 631.820 224.000 635.580 224.280 ;
        RECT 636.420 224.000 640.640 224.280 ;
        RECT 641.480 224.000 645.700 224.280 ;
        RECT 646.540 224.000 650.300 224.280 ;
        RECT 651.140 224.000 655.360 224.280 ;
        RECT 656.200 224.000 660.420 224.280 ;
        RECT 661.260 224.000 665.020 224.280 ;
        RECT 665.860 224.000 670.080 224.280 ;
        RECT 670.920 224.000 675.140 224.280 ;
        RECT 675.980 224.000 679.740 224.280 ;
        RECT 680.580 224.000 684.800 224.280 ;
        RECT 685.640 224.000 689.860 224.280 ;
        RECT 690.700 224.000 694.460 224.280 ;
        RECT 695.300 224.000 699.520 224.280 ;
        RECT 700.360 224.000 704.580 224.280 ;
        RECT 705.420 224.000 709.180 224.280 ;
        RECT 710.020 224.000 714.240 224.280 ;
        RECT 715.080 224.000 718.840 224.280 ;
        RECT 719.680 224.000 723.900 224.280 ;
        RECT 724.740 224.000 728.960 224.280 ;
        RECT 729.800 224.000 733.560 224.280 ;
        RECT 734.400 224.000 738.620 224.280 ;
        RECT 739.460 224.000 743.680 224.280 ;
        RECT 744.520 224.000 748.280 224.280 ;
        RECT 749.120 224.000 753.340 224.280 ;
        RECT 754.180 224.000 758.400 224.280 ;
        RECT 759.240 224.000 763.000 224.280 ;
        RECT 763.840 224.000 768.060 224.280 ;
        RECT 768.900 224.000 773.120 224.280 ;
        RECT 773.960 224.000 777.720 224.280 ;
        RECT 778.560 224.000 782.780 224.280 ;
        RECT 783.620 224.000 787.840 224.280 ;
        RECT 788.680 224.000 792.440 224.280 ;
        RECT 793.280 224.000 797.500 224.280 ;
        RECT 798.340 224.000 802.100 224.280 ;
        RECT 802.940 224.000 807.160 224.280 ;
        RECT 808.000 224.000 812.220 224.280 ;
        RECT 813.060 224.000 816.820 224.280 ;
        RECT 817.660 224.000 821.880 224.280 ;
        RECT 822.720 224.000 826.940 224.280 ;
        RECT 827.780 224.000 831.540 224.280 ;
        RECT 832.380 224.000 836.600 224.280 ;
        RECT 837.440 224.000 841.660 224.280 ;
        RECT 842.500 224.000 846.260 224.280 ;
        RECT 847.100 224.000 851.320 224.280 ;
        RECT 852.160 224.000 856.380 224.280 ;
        RECT 857.220 224.000 860.980 224.280 ;
        RECT 861.820 224.000 866.040 224.280 ;
        RECT 866.880 224.000 871.100 224.280 ;
        RECT 871.940 224.000 875.700 224.280 ;
        RECT 876.540 224.000 880.760 224.280 ;
        RECT 881.600 224.000 885.360 224.280 ;
        RECT 886.200 224.000 890.420 224.280 ;
        RECT 891.260 224.000 895.480 224.280 ;
        RECT 896.320 224.000 900.080 224.280 ;
        RECT 900.920 224.000 905.140 224.280 ;
        RECT 905.980 224.000 910.200 224.280 ;
        RECT 911.040 224.000 914.800 224.280 ;
        RECT 915.640 224.000 919.860 224.280 ;
        RECT 920.700 224.000 924.920 224.280 ;
        RECT 925.760 224.000 929.520 224.280 ;
        RECT 930.360 224.000 934.580 224.280 ;
        RECT 935.420 224.000 939.640 224.280 ;
        RECT 940.480 224.000 944.240 224.280 ;
        RECT 945.080 224.000 949.300 224.280 ;
        RECT 950.140 224.000 954.360 224.280 ;
        RECT 955.200 224.000 958.960 224.280 ;
        RECT 959.800 224.000 964.020 224.280 ;
        RECT 964.860 224.000 968.620 224.280 ;
        RECT 969.460 224.000 973.680 224.280 ;
        RECT 974.520 224.000 978.740 224.280 ;
        RECT 979.580 224.000 983.340 224.280 ;
        RECT 984.180 224.000 988.400 224.280 ;
        RECT 989.240 224.000 993.460 224.280 ;
        RECT 994.300 224.000 998.060 224.280 ;
        RECT 998.900 224.000 1003.120 224.280 ;
        RECT 1003.960 224.000 1008.180 224.280 ;
        RECT 1009.020 224.000 1012.780 224.280 ;
        RECT 1013.620 224.000 1017.840 224.280 ;
        RECT 1018.680 224.000 1022.900 224.280 ;
        RECT 1023.740 224.000 1027.500 224.280 ;
        RECT 1028.340 224.000 1032.560 224.280 ;
        RECT 1033.400 224.000 1037.620 224.280 ;
        RECT 1038.460 224.000 1042.220 224.280 ;
        RECT 1043.060 224.000 1047.280 224.280 ;
        RECT 1048.120 224.000 1051.880 224.280 ;
        RECT 1052.720 224.000 1056.940 224.280 ;
        RECT 1057.780 224.000 1062.000 224.280 ;
        RECT 1062.840 224.000 1066.600 224.280 ;
        RECT 1067.440 224.000 1071.660 224.280 ;
        RECT 1072.500 224.000 1076.720 224.280 ;
        RECT 1077.560 224.000 1081.320 224.280 ;
        RECT 1082.160 224.000 1086.380 224.280 ;
        RECT 1087.220 224.000 1091.440 224.280 ;
        RECT 1092.280 224.000 1096.040 224.280 ;
        RECT 1096.880 224.000 1101.100 224.280 ;
        RECT 1101.940 224.000 1106.160 224.280 ;
        RECT 1107.000 224.000 1110.760 224.280 ;
        RECT 1111.600 224.000 1115.820 224.280 ;
        RECT 1116.660 224.000 1120.880 224.280 ;
        RECT 1121.720 224.000 1125.480 224.280 ;
        RECT 1126.320 224.000 1130.540 224.280 ;
        RECT 1131.380 224.000 1135.140 224.280 ;
        RECT 1135.980 224.000 1140.200 224.280 ;
        RECT 1141.040 224.000 1145.260 224.280 ;
        RECT 1146.100 224.000 1149.860 224.280 ;
        RECT 1150.700 224.000 1154.920 224.280 ;
        RECT 1155.760 224.000 1159.980 224.280 ;
        RECT 1160.820 224.000 1164.580 224.280 ;
        RECT 1165.420 224.000 1169.640 224.280 ;
        RECT 1170.480 224.000 1174.700 224.280 ;
        RECT 1175.540 224.000 1179.300 224.280 ;
        RECT 1180.140 224.000 1184.360 224.280 ;
        RECT 1185.200 224.000 1189.420 224.280 ;
        RECT 1190.260 224.000 1194.020 224.280 ;
        RECT 1194.860 224.000 1199.080 224.280 ;
        RECT 1199.920 224.000 1204.140 224.280 ;
        RECT 1204.980 224.000 1208.740 224.280 ;
        RECT 1209.580 224.000 1213.800 224.280 ;
        RECT 1214.640 224.000 1218.400 224.280 ;
        RECT 1219.240 224.000 1223.460 224.280 ;
        RECT 1224.300 224.000 1228.520 224.280 ;
        RECT 1229.360 224.000 1233.120 224.280 ;
        RECT 1233.960 224.000 1238.180 224.280 ;
        RECT 1239.020 224.000 1243.240 224.280 ;
        RECT 1244.080 224.000 1247.840 224.280 ;
        RECT 1248.680 224.000 1252.900 224.280 ;
        RECT 1253.740 224.000 1257.960 224.280 ;
        RECT 1258.800 224.000 1262.560 224.280 ;
        RECT 1263.400 224.000 1267.620 224.280 ;
        RECT 1268.460 224.000 1272.680 224.280 ;
        RECT 1273.520 224.000 1277.280 224.280 ;
        RECT 1278.120 224.000 1282.340 224.280 ;
        RECT 1283.180 224.000 1287.400 224.280 ;
        RECT 1288.240 224.000 1292.000 224.280 ;
        RECT 1292.840 224.000 1297.060 224.280 ;
        RECT 1297.900 224.000 1301.660 224.280 ;
        RECT 1302.500 224.000 1306.720 224.280 ;
        RECT 1307.560 224.000 1311.780 224.280 ;
        RECT 1312.620 224.000 1316.380 224.280 ;
        RECT 1317.220 224.000 1321.440 224.280 ;
        RECT 1322.280 224.000 1326.500 224.280 ;
        RECT 1327.340 224.000 1331.100 224.280 ;
        RECT 1331.940 224.000 1336.160 224.280 ;
        RECT 1337.000 224.000 1341.220 224.280 ;
        RECT 1342.060 224.000 1345.820 224.280 ;
        RECT 1346.660 224.000 1350.880 224.280 ;
        RECT 1351.720 224.000 1355.940 224.280 ;
        RECT 1356.780 224.000 1360.540 224.280 ;
        RECT 1361.380 224.000 1365.600 224.280 ;
        RECT 1366.440 224.000 1370.660 224.280 ;
        RECT 1371.500 224.000 1375.260 224.280 ;
        RECT 1376.100 224.000 1380.320 224.280 ;
        RECT 1381.160 224.000 1384.920 224.280 ;
        RECT 1385.760 224.000 1389.980 224.280 ;
        RECT 1390.820 224.000 1395.040 224.280 ;
        RECT 1395.880 224.000 1399.640 224.280 ;
        RECT 1400.480 224.000 1404.700 224.280 ;
        RECT 1405.540 224.000 1409.760 224.280 ;
        RECT 1410.600 224.000 1414.360 224.280 ;
        RECT 1415.200 224.000 1419.420 224.280 ;
        RECT 1420.260 224.000 1424.480 224.280 ;
        RECT 1425.320 224.000 1429.080 224.280 ;
        RECT 1429.920 224.000 1434.140 224.280 ;
        RECT 1434.980 224.000 1439.200 224.280 ;
        RECT 1440.040 224.000 1443.800 224.280 ;
        RECT 1444.640 224.000 1448.860 224.280 ;
        RECT 1449.700 224.000 1453.920 224.280 ;
        RECT 1454.760 224.000 1458.520 224.280 ;
        RECT 1459.360 224.000 1463.580 224.280 ;
        RECT 1464.420 224.000 1468.180 224.280 ;
        RECT 1469.020 224.000 1473.240 224.280 ;
        RECT 1474.080 224.000 1478.300 224.280 ;
        RECT 1479.140 224.000 1482.900 224.280 ;
        RECT 1483.740 224.000 1487.960 224.280 ;
        RECT 1488.800 224.000 1493.020 224.280 ;
        RECT 1493.860 224.000 1497.620 224.280 ;
        RECT 1498.460 224.000 1502.680 224.280 ;
        RECT 1503.520 224.000 1507.740 224.280 ;
        RECT 1508.580 224.000 1512.340 224.280 ;
        RECT 1513.180 224.000 1517.400 224.280 ;
        RECT 1518.240 224.000 1522.460 224.280 ;
        RECT 1523.300 224.000 1527.060 224.280 ;
        RECT 1527.900 224.000 1532.120 224.280 ;
        RECT 1532.960 224.000 1537.180 224.280 ;
        RECT 1538.020 224.000 1541.780 224.280 ;
        RECT 1542.620 224.000 1546.840 224.280 ;
        RECT 1547.680 224.000 1551.440 224.280 ;
        RECT 1552.280 224.000 1556.500 224.280 ;
        RECT 1557.340 224.000 1561.560 224.280 ;
        RECT 1562.400 224.000 1566.160 224.280 ;
        RECT 1567.000 224.000 1571.220 224.280 ;
        RECT 1572.060 224.000 1576.280 224.280 ;
        RECT 1577.120 224.000 1580.880 224.280 ;
        RECT 1581.720 224.000 1585.940 224.280 ;
        RECT 1586.780 224.000 1591.000 224.280 ;
        RECT 1591.840 224.000 1595.600 224.280 ;
        RECT 1596.440 224.000 1600.660 224.280 ;
        RECT 1601.500 224.000 1605.720 224.280 ;
        RECT 1606.560 224.000 1610.320 224.280 ;
        RECT 1611.160 224.000 1615.380 224.280 ;
        RECT 1616.220 224.000 1620.440 224.280 ;
        RECT 1621.280 224.000 1625.040 224.280 ;
        RECT 1625.880 224.000 1630.100 224.280 ;
        RECT 1630.940 224.000 1634.700 224.280 ;
        RECT 1635.540 224.000 1639.760 224.280 ;
        RECT 1640.600 224.000 1644.820 224.280 ;
        RECT 1645.660 224.000 1649.420 224.280 ;
        RECT 1650.260 224.000 1654.480 224.280 ;
        RECT 1655.320 224.000 1659.540 224.280 ;
        RECT 1660.380 224.000 1664.140 224.280 ;
        RECT 1664.980 224.000 1669.200 224.280 ;
        RECT 1670.040 224.000 1674.260 224.280 ;
        RECT 1675.100 224.000 1678.860 224.280 ;
        RECT 1679.700 224.000 1683.920 224.280 ;
        RECT 1684.760 224.000 1688.980 224.280 ;
        RECT 1689.820 224.000 1693.580 224.280 ;
        RECT 1694.420 224.000 1698.640 224.280 ;
        RECT 1699.480 224.000 1703.700 224.280 ;
        RECT 1704.540 224.000 1708.300 224.280 ;
        RECT 1709.140 224.000 1713.360 224.280 ;
        RECT 1714.200 224.000 1717.960 224.280 ;
        RECT 1718.800 224.000 1723.020 224.280 ;
        RECT 1723.860 224.000 1728.080 224.280 ;
        RECT 1728.920 224.000 1732.680 224.280 ;
        RECT 1733.520 224.000 1737.740 224.280 ;
        RECT 1738.580 224.000 1742.800 224.280 ;
        RECT 1743.640 224.000 1747.400 224.280 ;
        RECT 1748.240 224.000 1752.460 224.280 ;
        RECT 1753.300 224.000 1757.520 224.280 ;
        RECT 1758.360 224.000 1762.120 224.280 ;
        RECT 1762.960 224.000 1767.180 224.280 ;
        RECT 1768.020 224.000 1772.240 224.280 ;
        RECT 1773.080 224.000 1776.840 224.280 ;
        RECT 1777.680 224.000 1781.900 224.280 ;
        RECT 1782.740 224.000 1786.960 224.280 ;
        RECT 1787.800 224.000 1791.560 224.280 ;
        RECT 1792.400 224.000 1796.620 224.280 ;
        RECT 1797.460 224.000 1801.220 224.280 ;
        RECT 1802.060 224.000 1806.280 224.280 ;
        RECT 1807.120 224.000 1811.340 224.280 ;
        RECT 1812.180 224.000 1815.940 224.280 ;
        RECT 1816.780 224.000 1821.000 224.280 ;
        RECT 1821.840 224.000 1826.060 224.280 ;
        RECT 1826.900 224.000 1830.660 224.280 ;
        RECT 1831.500 224.000 1835.720 224.280 ;
        RECT 1836.560 224.000 1840.780 224.280 ;
        RECT 1841.620 224.000 1845.380 224.280 ;
        RECT 1846.220 224.000 1850.440 224.280 ;
        RECT 1851.280 224.000 1855.500 224.280 ;
        RECT 1856.340 224.000 1860.100 224.280 ;
        RECT 1860.940 224.000 1865.160 224.280 ;
        RECT 1866.000 224.000 1870.220 224.280 ;
        RECT 1871.060 224.000 1874.820 224.280 ;
        RECT 1875.660 224.000 1879.880 224.280 ;
        RECT 1880.720 224.000 1884.480 224.280 ;
        RECT 1885.320 224.000 1889.540 224.280 ;
        RECT 1890.380 224.000 1894.600 224.280 ;
        RECT 1895.440 224.000 1899.200 224.280 ;
        RECT 1900.040 224.000 1904.260 224.280 ;
        RECT 1905.100 224.000 1909.320 224.280 ;
        RECT 1910.160 224.000 1913.920 224.280 ;
        RECT 1914.760 224.000 1918.980 224.280 ;
        RECT 1919.820 224.000 1924.040 224.280 ;
        RECT 1924.880 224.000 1928.640 224.280 ;
        RECT 1929.480 224.000 1933.700 224.280 ;
        RECT 1934.540 224.000 1938.760 224.280 ;
        RECT 1939.600 224.000 1943.360 224.280 ;
        RECT 1944.200 224.000 1948.420 224.280 ;
        RECT 1949.260 224.000 1953.480 224.280 ;
        RECT 1954.320 224.000 1958.080 224.280 ;
        RECT 1958.920 224.000 1963.140 224.280 ;
        RECT 1963.980 224.000 1967.740 224.280 ;
        RECT 1968.580 224.000 1972.800 224.280 ;
        RECT 1973.640 224.000 1977.860 224.280 ;
        RECT 1978.700 224.000 1982.460 224.280 ;
        RECT 1983.300 224.000 1987.520 224.280 ;
        RECT 1988.360 224.000 1992.580 224.280 ;
        RECT 1993.420 224.000 1997.180 224.280 ;
        RECT 1998.020 224.000 2002.240 224.280 ;
        RECT 2003.080 224.000 2007.300 224.280 ;
        RECT 2008.140 224.000 2011.900 224.280 ;
        RECT 2012.740 224.000 2016.960 224.280 ;
        RECT 2017.800 224.000 2022.020 224.280 ;
        RECT 2022.860 224.000 2026.620 224.280 ;
        RECT 2027.460 224.000 2031.680 224.280 ;
        RECT 2032.520 224.000 2036.740 224.280 ;
        RECT 2037.580 224.000 2041.340 224.280 ;
        RECT 2042.180 224.000 2046.400 224.280 ;
        RECT 2047.240 224.000 2051.000 224.280 ;
        RECT 2051.840 224.000 2056.060 224.280 ;
        RECT 2056.900 224.000 2061.120 224.280 ;
        RECT 2061.960 224.000 2065.720 224.280 ;
        RECT 2066.560 224.000 2070.780 224.280 ;
        RECT 2071.620 224.000 2075.840 224.280 ;
        RECT 2076.680 224.000 2080.440 224.280 ;
        RECT 2081.280 224.000 2085.500 224.280 ;
        RECT 2086.340 224.000 2090.560 224.280 ;
        RECT 2091.400 224.000 2095.160 224.280 ;
        RECT 2096.000 224.000 2100.220 224.280 ;
        RECT 2101.060 224.000 2105.280 224.280 ;
        RECT 2106.120 224.000 2109.880 224.280 ;
        RECT 2110.720 224.000 2114.940 224.280 ;
        RECT 2115.780 224.000 2120.000 224.280 ;
        RECT 2120.840 224.000 2124.600 224.280 ;
        RECT 2125.440 224.000 2129.660 224.280 ;
        RECT 2130.500 224.000 2134.260 224.280 ;
        RECT 2135.100 224.000 2139.320 224.280 ;
        RECT 2140.160 224.000 2144.380 224.280 ;
        RECT 2145.220 224.000 2148.980 224.280 ;
        RECT 2149.820 224.000 2154.040 224.280 ;
        RECT 2154.880 224.000 2159.100 224.280 ;
        RECT 2159.940 224.000 2163.700 224.280 ;
        RECT 2164.540 224.000 2168.760 224.280 ;
        RECT 2169.600 224.000 2173.820 224.280 ;
        RECT 2174.660 224.000 2178.420 224.280 ;
        RECT 2179.260 224.000 2183.480 224.280 ;
        RECT 2184.320 224.000 2188.540 224.280 ;
        RECT 2189.380 224.000 2193.140 224.280 ;
        RECT 2193.980 224.000 2198.200 224.280 ;
        RECT 2199.040 224.000 2203.260 224.280 ;
        RECT 2204.100 224.000 2207.860 224.280 ;
        RECT 2208.700 224.000 2212.920 224.280 ;
        RECT 2213.760 224.000 2217.520 224.280 ;
        RECT 2218.360 224.000 2222.580 224.280 ;
        RECT 2223.420 224.000 2227.640 224.280 ;
        RECT 2228.480 224.000 2232.240 224.280 ;
        RECT 2233.080 224.000 2237.300 224.280 ;
        RECT 2238.140 224.000 2242.360 224.280 ;
        RECT 2243.200 224.000 2246.960 224.280 ;
        RECT 2247.800 224.000 2252.020 224.280 ;
        RECT 2252.860 224.000 2257.080 224.280 ;
        RECT 2257.920 224.000 2261.680 224.280 ;
        RECT 2262.520 224.000 2266.740 224.280 ;
        RECT 2267.580 224.000 2271.800 224.280 ;
        RECT 2272.640 224.000 2276.400 224.280 ;
        RECT 2277.240 224.000 2281.460 224.280 ;
        RECT 2282.300 224.000 2286.520 224.280 ;
        RECT 2287.360 224.000 2291.120 224.280 ;
        RECT 2291.960 224.000 2296.180 224.280 ;
        RECT 2297.020 224.000 2300.780 224.280 ;
        RECT 2301.620 224.000 2305.840 224.280 ;
        RECT 2306.680 224.000 2310.900 224.280 ;
        RECT 2311.740 224.000 2315.500 224.280 ;
        RECT 2316.340 224.000 2320.560 224.280 ;
        RECT 2321.400 224.000 2325.620 224.280 ;
        RECT 2326.460 224.000 2330.220 224.280 ;
        RECT 2331.060 224.000 2335.280 224.280 ;
        RECT 2336.120 224.000 2340.340 224.280 ;
        RECT 2341.180 224.000 2344.940 224.280 ;
        RECT 2345.780 224.000 2350.000 224.280 ;
        RECT 2350.840 224.000 2355.060 224.280 ;
        RECT 2355.900 224.000 2359.660 224.280 ;
        RECT 2360.500 224.000 2364.720 224.280 ;
        RECT 2365.560 224.000 2369.780 224.280 ;
        RECT 2370.620 224.000 2374.380 224.280 ;
        RECT 2375.220 224.000 2379.440 224.280 ;
        RECT 2380.280 224.000 2384.040 224.280 ;
        RECT 2384.880 224.000 2389.100 224.280 ;
        RECT 2389.940 224.000 2394.160 224.280 ;
        RECT 2395.000 224.000 2398.760 224.280 ;
        RECT 2399.600 224.000 2403.820 224.280 ;
        RECT 2404.660 224.000 2408.880 224.280 ;
        RECT 2409.720 224.000 2413.480 224.280 ;
        RECT 2414.320 224.000 2418.540 224.280 ;
        RECT 2419.380 224.000 2423.600 224.280 ;
        RECT 2424.440 224.000 2428.200 224.280 ;
        RECT 2429.040 224.000 2433.260 224.280 ;
        RECT 2434.100 224.000 2438.320 224.280 ;
        RECT 2439.160 224.000 2442.920 224.280 ;
        RECT 2443.760 224.000 2447.980 224.280 ;
        RECT 2448.820 224.000 2453.040 224.280 ;
        RECT 2453.880 224.000 2457.640 224.280 ;
        RECT 2458.480 224.000 2462.700 224.280 ;
        RECT 2463.540 224.000 2467.300 224.280 ;
        RECT 2468.140 224.000 2472.360 224.280 ;
        RECT 2473.200 224.000 2477.420 224.280 ;
        RECT 2478.260 224.000 2482.020 224.280 ;
        RECT 2482.860 224.000 2487.080 224.280 ;
        RECT 2487.920 224.000 2492.140 224.280 ;
        RECT 2492.980 224.000 2496.740 224.280 ;
        RECT 2497.580 224.000 2501.800 224.280 ;
        RECT 2502.640 224.000 2506.860 224.280 ;
        RECT 2507.700 224.000 2511.460 224.280 ;
        RECT 2512.300 224.000 2516.520 224.280 ;
        RECT 2517.360 224.000 2521.580 224.280 ;
        RECT 2522.420 224.000 2526.180 224.280 ;
        RECT 2527.020 224.000 2531.240 224.280 ;
        RECT 2532.080 224.000 2536.300 224.280 ;
        RECT 2537.140 224.000 2540.900 224.280 ;
        RECT 2541.740 224.000 2545.960 224.280 ;
        RECT 2546.800 224.000 2550.560 224.280 ;
        RECT 2551.400 224.000 2555.620 224.280 ;
        RECT 2556.460 224.000 2560.680 224.280 ;
        RECT 2561.520 224.000 2565.280 224.280 ;
        RECT 2566.120 224.000 2570.340 224.280 ;
        RECT 2571.180 224.000 2575.400 224.280 ;
        RECT 2576.240 224.000 2580.000 224.280 ;
        RECT 2580.840 224.000 2585.060 224.280 ;
        RECT 2585.900 224.000 2590.120 224.280 ;
        RECT 2590.960 224.000 2594.720 224.280 ;
        RECT 2595.560 224.000 2599.780 224.280 ;
        RECT 2600.620 224.000 2604.840 224.280 ;
        RECT 2605.680 224.000 2609.440 224.280 ;
      LAYER met3 ;
        RECT 228.275 224.255 2606.345 3207.745 ;
      LAYER met4 ;
        RECT 243.685 230.640 274.020 3206.800 ;
        RECT 277.020 230.640 292.020 3206.800 ;
        RECT 295.020 230.640 310.020 3206.800 ;
        RECT 313.020 230.640 315.070 3206.800 ;
      LAYER met4 ;
        RECT 315.470 230.640 317.070 3206.800 ;
      LAYER met4 ;
        RECT 317.470 230.640 328.020 3206.800 ;
        RECT 331.020 230.640 364.020 3206.800 ;
        RECT 367.020 230.640 382.020 3206.800 ;
        RECT 385.020 230.640 400.020 3206.800 ;
        RECT 403.020 230.640 418.020 3206.800 ;
        RECT 421.020 230.640 454.020 3206.800 ;
        RECT 457.020 230.640 472.020 3206.800 ;
        RECT 475.020 230.640 490.020 3206.800 ;
        RECT 493.020 230.640 508.020 3206.800 ;
        RECT 511.020 230.640 544.020 3206.800 ;
        RECT 547.020 230.640 562.020 3206.800 ;
        RECT 565.020 230.640 580.020 3206.800 ;
        RECT 583.020 230.640 598.020 3206.800 ;
        RECT 601.020 230.640 634.020 3206.800 ;
        RECT 637.020 230.640 652.020 3206.800 ;
        RECT 655.020 230.640 670.020 3206.800 ;
        RECT 673.020 230.640 688.020 3206.800 ;
        RECT 691.020 230.640 724.020 3206.800 ;
        RECT 727.020 230.640 742.020 3206.800 ;
        RECT 745.020 230.640 760.020 3206.800 ;
        RECT 763.020 230.640 778.020 3206.800 ;
        RECT 781.020 230.640 814.020 3206.800 ;
        RECT 817.020 230.640 832.020 3206.800 ;
        RECT 835.020 230.640 850.020 3206.800 ;
        RECT 853.020 230.640 868.020 3206.800 ;
        RECT 871.020 230.640 904.020 3206.800 ;
        RECT 907.020 230.640 922.020 3206.800 ;
        RECT 925.020 230.640 940.020 3206.800 ;
        RECT 943.020 230.640 958.020 3206.800 ;
        RECT 961.020 230.640 994.020 3206.800 ;
        RECT 997.020 230.640 1012.020 3206.800 ;
        RECT 1015.020 230.640 1030.020 3206.800 ;
        RECT 1033.020 230.640 1048.020 3206.800 ;
        RECT 1051.020 230.640 1084.020 3206.800 ;
        RECT 1087.020 230.640 1102.020 3206.800 ;
        RECT 1105.020 230.640 1120.020 3206.800 ;
        RECT 1123.020 230.640 1138.020 3206.800 ;
        RECT 1141.020 230.640 1174.020 3206.800 ;
        RECT 1177.020 230.640 1192.020 3206.800 ;
        RECT 1195.020 230.640 1210.020 3206.800 ;
        RECT 1213.020 230.640 1228.020 3206.800 ;
        RECT 1231.020 230.640 1264.020 3206.800 ;
        RECT 1267.020 230.640 1282.020 3206.800 ;
        RECT 1285.020 230.640 1300.020 3206.800 ;
        RECT 1303.020 230.640 1318.020 3206.800 ;
        RECT 1321.020 230.640 1354.020 3206.800 ;
        RECT 1357.020 230.640 1372.020 3206.800 ;
        RECT 1375.020 230.640 1390.020 3206.800 ;
        RECT 1393.020 230.640 1408.020 3206.800 ;
        RECT 1411.020 230.640 1444.020 3206.800 ;
        RECT 1447.020 230.640 1462.020 3206.800 ;
        RECT 1465.020 230.640 1480.020 3206.800 ;
        RECT 1483.020 230.640 1498.020 3206.800 ;
        RECT 1501.020 230.640 1534.020 3206.800 ;
        RECT 1537.020 230.640 1552.020 3206.800 ;
        RECT 1555.020 230.640 1570.020 3206.800 ;
        RECT 1573.020 230.640 1588.020 3206.800 ;
        RECT 1591.020 230.640 1624.020 3206.800 ;
        RECT 1627.020 230.640 1642.020 3206.800 ;
        RECT 1645.020 230.640 1660.020 3206.800 ;
        RECT 1663.020 230.640 1678.020 3206.800 ;
        RECT 1681.020 230.640 1714.020 3206.800 ;
        RECT 1717.020 230.640 1732.020 3206.800 ;
        RECT 1735.020 230.640 1750.020 3206.800 ;
        RECT 1753.020 230.640 1768.020 3206.800 ;
        RECT 1771.020 230.640 1804.020 3206.800 ;
        RECT 1807.020 230.640 1822.020 3206.800 ;
        RECT 1825.020 230.640 1840.020 3206.800 ;
        RECT 1843.020 230.640 1858.020 3206.800 ;
        RECT 1861.020 230.640 1894.020 3206.800 ;
        RECT 1897.020 230.640 1912.020 3206.800 ;
        RECT 1915.020 230.640 1930.020 3206.800 ;
        RECT 1933.020 230.640 1948.020 3206.800 ;
        RECT 1951.020 230.640 1984.020 3206.800 ;
        RECT 1987.020 230.640 2002.020 3206.800 ;
        RECT 2005.020 230.640 2020.020 3206.800 ;
        RECT 2023.020 230.640 2038.020 3206.800 ;
        RECT 2041.020 230.640 2074.020 3206.800 ;
        RECT 2077.020 230.640 2092.020 3206.800 ;
        RECT 2095.020 230.640 2110.020 3206.800 ;
        RECT 2113.020 230.640 2128.020 3206.800 ;
        RECT 2131.020 230.640 2164.020 3206.800 ;
        RECT 2167.020 230.640 2182.020 3206.800 ;
        RECT 2185.020 230.640 2200.020 3206.800 ;
        RECT 2203.020 230.640 2218.020 3206.800 ;
        RECT 2221.020 230.640 2254.020 3206.800 ;
        RECT 2257.020 230.640 2272.020 3206.800 ;
        RECT 2275.020 230.640 2290.020 3206.800 ;
        RECT 2293.020 230.640 2308.020 3206.800 ;
        RECT 2311.020 230.640 2344.020 3206.800 ;
        RECT 2347.020 230.640 2362.020 3206.800 ;
        RECT 2365.020 230.640 2380.020 3206.800 ;
        RECT 2383.020 230.640 2398.020 3206.800 ;
        RECT 2401.020 230.640 2434.020 3206.800 ;
        RECT 2437.020 230.640 2452.020 3206.800 ;
        RECT 2455.020 230.640 2470.020 3206.800 ;
        RECT 2473.020 230.640 2488.020 3206.800 ;
        RECT 2491.020 230.640 2524.020 3206.800 ;
        RECT 2527.020 230.640 2542.020 3206.800 ;
        RECT 2545.020 230.640 2560.020 3206.800 ;
        RECT 2563.020 230.640 2574.375 3206.800 ;
  END
END user_project_wrapper
END LIBRARY

