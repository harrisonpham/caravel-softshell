magic
tech sky130A
magscale 1 2
timestamp 1608291739
<< metal1 >>
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 325694 700992 325700 701004
rect 154172 700964 325700 700992
rect 154172 700952 154178 700964
rect 325694 700952 325700 700964
rect 325752 700952 325758 701004
rect 137830 700884 137836 700936
rect 137888 700924 137894 700936
rect 321554 700924 321560 700936
rect 137888 700896 321560 700924
rect 137888 700884 137894 700896
rect 321554 700884 321560 700896
rect 321612 700884 321618 700936
rect 256602 700816 256608 700868
rect 256660 700856 256666 700868
rect 462314 700856 462320 700868
rect 256660 700828 462320 700856
rect 256660 700816 256666 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 262122 700748 262128 700800
rect 262180 700788 262186 700800
rect 478506 700788 478512 700800
rect 262180 700760 478512 700788
rect 262180 700748 262186 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 339494 700720 339500 700732
rect 89220 700692 339500 700720
rect 89220 700680 89226 700692
rect 339494 700680 339500 700692
rect 339552 700680 339558 700732
rect 72970 700612 72976 700664
rect 73028 700652 73034 700664
rect 335354 700652 335360 700664
rect 73028 700624 335360 700652
rect 73028 700612 73034 700624
rect 335354 700612 335360 700624
rect 335412 700612 335418 700664
rect 244182 700544 244188 700596
rect 244240 700584 244246 700596
rect 527174 700584 527180 700596
rect 244240 700556 527180 700584
rect 244240 700544 244246 700556
rect 527174 700544 527180 700556
rect 527232 700544 527238 700596
rect 248322 700476 248328 700528
rect 248380 700516 248386 700528
rect 543458 700516 543464 700528
rect 248380 700488 543464 700516
rect 248380 700476 248386 700488
rect 543458 700476 543464 700488
rect 543516 700476 543522 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 343634 700448 343640 700460
rect 40552 700420 343640 700448
rect 40552 700408 40558 700420
rect 343634 700408 343640 700420
rect 343692 700408 343698 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 351914 700380 351920 700392
rect 24360 700352 351920 700380
rect 24360 700340 24366 700352
rect 351914 700340 351920 700352
rect 351972 700340 351978 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 347774 700312 347780 700324
rect 8168 700284 347780 700312
rect 8168 700272 8174 700284
rect 347774 700272 347780 700284
rect 347832 700272 347838 700324
rect 274542 700204 274548 700256
rect 274600 700244 274606 700256
rect 413646 700244 413652 700256
rect 274600 700216 413652 700244
rect 274600 700204 274606 700216
rect 413646 700204 413652 700216
rect 413704 700204 413710 700256
rect 270402 700136 270408 700188
rect 270460 700176 270466 700188
rect 397454 700176 397460 700188
rect 270460 700148 397460 700176
rect 270460 700136 270466 700148
rect 397454 700136 397460 700148
rect 397512 700136 397518 700188
rect 202782 700068 202788 700120
rect 202840 700108 202846 700120
rect 309134 700108 309140 700120
rect 202840 700080 309140 700108
rect 202840 700068 202846 700080
rect 309134 700068 309140 700080
rect 309192 700068 309198 700120
rect 218974 700000 218980 700052
rect 219032 700040 219038 700052
rect 313274 700040 313280 700052
rect 219032 700012 313280 700040
rect 219032 700000 219038 700012
rect 313274 700000 313280 700012
rect 313332 700000 313338 700052
rect 288342 699932 288348 699984
rect 288400 699972 288406 699984
rect 348786 699972 348792 699984
rect 288400 699944 348792 699972
rect 288400 699932 288406 699944
rect 348786 699932 348792 699944
rect 348844 699932 348850 699984
rect 284202 699864 284208 699916
rect 284260 699904 284266 699916
rect 332502 699904 332508 699916
rect 284260 699876 332508 699904
rect 284260 699864 284266 699876
rect 332502 699864 332508 699876
rect 332560 699864 332566 699916
rect 267642 699796 267648 699848
rect 267700 699836 267706 699848
rect 295334 699836 295340 699848
rect 267700 699808 295340 699836
rect 267700 699796 267706 699808
rect 295334 699796 295340 699808
rect 295392 699796 295398 699848
rect 283834 699728 283840 699780
rect 283892 699768 283898 699780
rect 299474 699768 299480 699780
rect 283892 699740 299480 699768
rect 283892 699728 283898 699740
rect 299474 699728 299480 699740
rect 299532 699728 299538 699780
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 230382 696940 230388 696992
rect 230440 696980 230446 696992
rect 580166 696980 580172 696992
rect 230440 696952 580172 696980
rect 230440 696940 230446 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 299566 692792 299572 692844
rect 299624 692832 299630 692844
rect 300210 692832 300216 692844
rect 299624 692804 300216 692832
rect 299624 692792 299630 692804
rect 300210 692792 300216 692804
rect 300268 692792 300274 692844
rect 364334 692792 364340 692844
rect 364392 692832 364398 692844
rect 365070 692832 365076 692844
rect 364392 692804 365076 692832
rect 364392 692792 364398 692804
rect 365070 692792 365076 692804
rect 365128 692792 365134 692844
rect 429194 692792 429200 692844
rect 429252 692832 429258 692844
rect 429930 692832 429936 692844
rect 429252 692804 429936 692832
rect 429252 692792 429258 692804
rect 429930 692792 429936 692804
rect 429988 692792 429994 692844
rect 494054 692792 494060 692844
rect 494112 692832 494118 692844
rect 494882 692832 494888 692844
rect 494112 692804 494888 692832
rect 494112 692792 494118 692804
rect 494882 692792 494888 692804
rect 494940 692792 494946 692844
rect 558914 692792 558920 692844
rect 558972 692832 558978 692844
rect 559742 692832 559748 692844
rect 558972 692804 559748 692832
rect 558972 692792 558978 692804
rect 559742 692792 559748 692804
rect 559800 692792 559806 692844
rect 229094 690684 229100 690736
rect 229152 690724 229158 690736
rect 230382 690724 230388 690736
rect 229152 690696 230388 690724
rect 229152 690684 229158 690696
rect 230382 690684 230388 690696
rect 230440 690684 230446 690736
rect 242894 690684 242900 690736
rect 242952 690724 242958 690736
rect 244182 690724 244188 690736
rect 242952 690696 244188 690724
rect 242952 690684 242958 690696
rect 244182 690684 244188 690696
rect 244240 690684 244246 690736
rect 247034 690684 247040 690736
rect 247092 690724 247098 690736
rect 248322 690724 248328 690736
rect 247092 690696 248328 690724
rect 247092 690684 247098 690696
rect 248322 690684 248328 690696
rect 248380 690684 248386 690736
rect 255314 690684 255320 690736
rect 255372 690724 255378 690736
rect 256602 690724 256608 690736
rect 255372 690696 256608 690724
rect 255372 690684 255378 690696
rect 256602 690684 256608 690696
rect 256660 690684 256666 690736
rect 260834 690684 260840 690736
rect 260892 690724 260898 690736
rect 262122 690724 262128 690736
rect 260892 690696 262128 690724
rect 260892 690684 260898 690696
rect 262122 690684 262128 690696
rect 262180 690684 262186 690736
rect 269114 690684 269120 690736
rect 269172 690724 269178 690736
rect 270402 690724 270408 690736
rect 269172 690696 270408 690724
rect 269172 690684 269178 690696
rect 270402 690684 270408 690696
rect 270460 690684 270466 690736
rect 273254 690684 273260 690736
rect 273312 690724 273318 690736
rect 274542 690724 274548 690736
rect 273312 690696 274548 690724
rect 273312 690684 273318 690696
rect 274542 690684 274548 690696
rect 274600 690684 274606 690736
rect 291930 688372 291936 688424
rect 291988 688412 291994 688424
rect 299566 688412 299572 688424
rect 291988 688384 299572 688412
rect 291988 688372 291994 688384
rect 299566 688372 299572 688384
rect 299624 688372 299630 688424
rect 235902 688304 235908 688356
rect 235960 688344 235966 688356
rect 304442 688344 304448 688356
rect 235960 688316 304448 688344
rect 235960 688304 235966 688316
rect 304442 688304 304448 688316
rect 304500 688304 304506 688356
rect 278682 688236 278688 688288
rect 278740 688276 278746 688288
rect 364334 688276 364340 688288
rect 278740 688248 364340 688276
rect 278740 688236 278746 688248
rect 364334 688236 364340 688248
rect 364392 688236 364398 688288
rect 171042 688168 171048 688220
rect 171100 688208 171106 688220
rect 317598 688208 317604 688220
rect 171100 688180 317604 688208
rect 171100 688168 171106 688180
rect 317598 688168 317604 688180
rect 317656 688168 317662 688220
rect 264974 688100 264980 688152
rect 265032 688140 265038 688152
rect 429194 688140 429200 688152
rect 265032 688112 429200 688140
rect 265032 688100 265038 688112
rect 429194 688100 429200 688112
rect 429252 688100 429258 688152
rect 106182 688072 106188 688084
rect 106141 688044 106188 688072
rect 106182 688032 106188 688044
rect 106240 688072 106246 688084
rect 330754 688072 330760 688084
rect 106240 688044 330760 688072
rect 106240 688032 106246 688044
rect 330754 688032 330760 688044
rect 330812 688032 330818 688084
rect 251174 687964 251180 688016
rect 251232 688004 251238 688016
rect 494054 688004 494060 688016
rect 251232 687976 494060 688004
rect 251232 687964 251238 687976
rect 494054 687964 494060 687976
rect 494112 687964 494118 688016
rect 238754 687896 238760 687948
rect 238812 687936 238818 687948
rect 558914 687936 558920 687948
rect 238812 687908 558920 687936
rect 238812 687896 238818 687908
rect 558914 687896 558920 687908
rect 558972 687896 558978 687948
rect 229002 687216 229008 687268
rect 229060 687256 229066 687268
rect 230014 687256 230020 687268
rect 229060 687228 230020 687256
rect 229060 687216 229066 687228
rect 230014 687216 230020 687228
rect 230072 687216 230078 687268
rect 283190 687216 283196 687268
rect 283248 687256 283254 687268
rect 284202 687256 284208 687268
rect 283248 687228 284208 687256
rect 283248 687216 283254 687228
rect 284202 687216 284208 687228
rect 284260 687216 284266 687268
rect 124214 687148 124220 687200
rect 124272 687188 124278 687200
rect 379422 687188 379428 687200
rect 124272 687160 379428 687188
rect 124272 687148 124278 687160
rect 379422 687148 379428 687160
rect 379480 687148 379486 687200
rect 111794 687080 111800 687132
rect 111852 687120 111858 687132
rect 365898 687120 365904 687132
rect 111852 687092 365904 687120
rect 111852 687080 111858 687092
rect 365898 687080 365904 687092
rect 365956 687080 365962 687132
rect 150434 687012 150440 687064
rect 150492 687052 150498 687064
rect 411162 687052 411168 687064
rect 150492 687024 411168 687052
rect 150492 687012 150498 687024
rect 411162 687012 411168 687024
rect 411220 687012 411226 687064
rect 63862 686944 63868 686996
rect 63920 686984 63926 686996
rect 229002 686984 229008 686996
rect 63920 686956 229008 686984
rect 63920 686944 63926 686956
rect 229002 686944 229008 686956
rect 229060 686944 229066 686996
rect 229094 686944 229100 686996
rect 229152 686984 229158 686996
rect 229922 686984 229928 686996
rect 229152 686956 229928 686984
rect 229152 686944 229158 686956
rect 229922 686944 229928 686956
rect 229980 686944 229986 686996
rect 230014 686944 230020 686996
rect 230072 686984 230078 686996
rect 233234 686984 233240 686996
rect 230072 686956 233240 686984
rect 230072 686944 230078 686956
rect 233234 686944 233240 686956
rect 233292 686944 233298 686996
rect 234614 686944 234620 686996
rect 234672 686984 234678 686996
rect 580166 686984 580172 686996
rect 234672 686956 580172 686984
rect 234672 686944 234678 686956
rect 580166 686944 580172 686956
rect 580224 686944 580230 686996
rect 168374 686876 168380 686928
rect 168432 686916 168438 686928
rect 539318 686916 539324 686928
rect 168432 686888 539324 686916
rect 168432 686876 168438 686888
rect 539318 686876 539324 686888
rect 539376 686876 539382 686928
rect 164234 686808 164240 686860
rect 164292 686848 164298 686860
rect 540330 686848 540336 686860
rect 164292 686820 540336 686848
rect 164292 686808 164298 686820
rect 540330 686808 540336 686820
rect 540388 686808 540394 686860
rect 154574 686740 154580 686792
rect 154632 686780 154638 686792
rect 541710 686780 541716 686792
rect 154632 686752 541716 686780
rect 154632 686740 154638 686752
rect 541710 686740 541716 686752
rect 541768 686740 541774 686792
rect 2866 686672 2872 686724
rect 2924 686712 2930 686724
rect 405734 686712 405740 686724
rect 2924 686684 405740 686712
rect 2924 686672 2930 686684
rect 405734 686672 405740 686684
rect 405792 686672 405798 686724
rect 128354 686604 128360 686656
rect 128412 686644 128418 686656
rect 539042 686644 539048 686656
rect 128412 686616 539048 686644
rect 128412 686604 128418 686616
rect 539042 686604 539048 686616
rect 539100 686604 539106 686656
rect 4982 686536 4988 686588
rect 5040 686576 5046 686588
rect 418522 686576 418528 686588
rect 5040 686548 418528 686576
rect 5040 686536 5046 686548
rect 418522 686536 418528 686548
rect 418580 686536 418586 686588
rect 115934 686468 115940 686520
rect 115992 686508 115998 686520
rect 538950 686508 538956 686520
rect 115992 686480 538956 686508
rect 115992 686468 115998 686480
rect 538950 686468 538956 686480
rect 539008 686468 539014 686520
rect 102134 686400 102140 686452
rect 102192 686440 102198 686452
rect 538858 686440 538864 686452
rect 102192 686412 538864 686440
rect 102192 686400 102198 686412
rect 538858 686400 538864 686412
rect 538916 686400 538922 686452
rect 7558 686332 7564 686384
rect 7616 686372 7622 686384
rect 444834 686372 444840 686384
rect 7616 686344 444840 686372
rect 7616 686332 7622 686344
rect 444834 686332 444840 686344
rect 444892 686332 444898 686384
rect 3050 686264 3056 686316
rect 3108 686304 3114 686316
rect 440418 686304 440424 686316
rect 3108 686276 440424 686304
rect 3108 686264 3114 686276
rect 440418 686264 440424 686276
rect 440476 686264 440482 686316
rect 132494 686196 132500 686248
rect 132552 686236 132558 686248
rect 577774 686236 577780 686248
rect 132552 686208 577780 686236
rect 132552 686196 132558 686208
rect 577774 686196 577780 686208
rect 577832 686196 577838 686248
rect 3234 686128 3240 686180
rect 3292 686168 3298 686180
rect 453574 686168 453580 686180
rect 3292 686140 453580 686168
rect 3292 686128 3298 686140
rect 453574 686128 453580 686140
rect 453632 686128 453638 686180
rect 3326 686060 3332 686112
rect 3384 686100 3390 686112
rect 471146 686100 471152 686112
rect 3384 686072 471152 686100
rect 3384 686060 3390 686072
rect 471146 686060 471152 686072
rect 471204 686060 471210 686112
rect 106274 685992 106280 686044
rect 106332 686032 106338 686044
rect 577682 686032 577688 686044
rect 106332 686004 577688 686032
rect 106332 685992 106338 686004
rect 577682 685992 577688 686004
rect 577740 685992 577746 686044
rect 4062 685924 4068 685976
rect 4120 685964 4126 685976
rect 484394 685964 484400 685976
rect 4120 685936 484400 685964
rect 4120 685924 4126 685936
rect 484394 685924 484400 685936
rect 484452 685924 484458 685976
rect 39850 685856 39856 685908
rect 39908 685896 39914 685908
rect 49694 685896 49700 685908
rect 39908 685868 49700 685896
rect 39908 685856 39914 685868
rect 49694 685856 49700 685868
rect 49752 685856 49758 685908
rect 93854 685856 93860 685908
rect 93912 685896 93918 685908
rect 577590 685896 577596 685908
rect 93912 685868 577596 685896
rect 93912 685856 93918 685868
rect 577590 685856 577596 685868
rect 577648 685856 577654 685908
rect 226150 685788 226156 685840
rect 226208 685828 226214 685840
rect 540882 685828 540888 685840
rect 226208 685800 540888 685828
rect 226208 685788 226214 685800
rect 540882 685788 540888 685800
rect 540940 685788 540946 685840
rect 212994 685720 213000 685772
rect 213052 685760 213058 685772
rect 540698 685760 540704 685772
rect 213052 685732 540704 685760
rect 213052 685720 213058 685732
rect 540698 685720 540704 685732
rect 540756 685720 540762 685772
rect 199838 685652 199844 685704
rect 199896 685692 199902 685704
rect 540514 685692 540520 685704
rect 199896 685664 540520 685692
rect 199896 685652 199902 685664
rect 540514 685652 540520 685664
rect 540572 685652 540578 685704
rect 5534 685584 5540 685636
rect 5592 685624 5598 685636
rect 357434 685624 357440 685636
rect 5592 685596 357440 685624
rect 5592 685584 5598 685596
rect 357434 685584 357440 685596
rect 357492 685584 357498 685636
rect 186682 685516 186688 685568
rect 186740 685556 186746 685568
rect 539502 685556 539508 685568
rect 186740 685528 539508 685556
rect 186740 685516 186746 685528
rect 539502 685516 539508 685528
rect 539560 685516 539566 685568
rect 217410 685448 217416 685500
rect 217468 685488 217474 685500
rect 578142 685488 578148 685500
rect 217468 685460 578148 685488
rect 217468 685448 217474 685460
rect 578142 685448 578148 685460
rect 578200 685448 578206 685500
rect 6730 685380 6736 685432
rect 6788 685420 6794 685432
rect 370222 685420 370228 685432
rect 6788 685392 370228 685420
rect 6788 685380 6794 685392
rect 370222 685380 370228 685392
rect 370280 685380 370286 685432
rect 173526 685312 173532 685364
rect 173584 685352 173590 685364
rect 539410 685352 539416 685364
rect 173584 685324 539416 685352
rect 173584 685312 173590 685324
rect 539410 685312 539416 685324
rect 539468 685312 539474 685364
rect 204162 685244 204168 685296
rect 204220 685284 204226 685296
rect 578050 685284 578056 685296
rect 204220 685256 578056 685284
rect 204220 685244 204226 685256
rect 578050 685244 578056 685256
rect 578108 685244 578114 685296
rect 6638 685176 6644 685228
rect 6696 685216 6702 685228
rect 383746 685216 383752 685228
rect 6696 685188 383752 685216
rect 6696 685176 6702 685188
rect 383746 685176 383752 685188
rect 383804 685176 383810 685228
rect 411162 685176 411168 685228
rect 411220 685216 411226 685228
rect 579982 685216 579988 685228
rect 411220 685188 579988 685216
rect 411220 685176 411226 685188
rect 579982 685176 579988 685188
rect 580040 685176 580046 685228
rect 191006 685108 191012 685160
rect 191064 685148 191070 685160
rect 577958 685148 577964 685160
rect 191064 685120 577964 685148
rect 191064 685108 191070 685120
rect 577958 685108 577964 685120
rect 578016 685108 578022 685160
rect 25590 685040 25596 685092
rect 25648 685080 25654 685092
rect 414106 685080 414112 685092
rect 25648 685052 414112 685080
rect 25648 685040 25654 685052
rect 414106 685040 414112 685052
rect 414164 685040 414170 685092
rect 6546 684972 6552 685024
rect 6604 685012 6610 685024
rect 396534 685012 396540 685024
rect 6604 684984 396540 685012
rect 6604 684972 6610 684984
rect 396534 684972 396540 684984
rect 396592 684972 396598 685024
rect 147214 684904 147220 684956
rect 147272 684944 147278 684956
rect 541618 684944 541624 684956
rect 147272 684916 541624 684944
rect 147272 684904 147278 684916
rect 541618 684904 541624 684916
rect 541676 684904 541682 684956
rect 177850 684836 177856 684888
rect 177908 684876 177914 684888
rect 579798 684876 579804 684888
rect 177908 684848 579804 684876
rect 177908 684836 177914 684848
rect 579798 684836 579804 684848
rect 579856 684836 579862 684888
rect 6454 684768 6460 684820
rect 6512 684808 6518 684820
rect 409874 684808 409880 684820
rect 6512 684780 409880 684808
rect 6512 684768 6518 684780
rect 409874 684768 409880 684780
rect 409932 684768 409938 684820
rect 6362 684700 6368 684752
rect 6420 684740 6426 684752
rect 422846 684740 422852 684752
rect 6420 684712 422852 684740
rect 6420 684700 6426 684712
rect 422846 684700 422852 684712
rect 422904 684700 422910 684752
rect 160370 684632 160376 684684
rect 160428 684672 160434 684684
rect 577866 684672 577872 684684
rect 160428 684644 577872 684672
rect 160428 684632 160434 684644
rect 577866 684632 577872 684644
rect 577924 684632 577930 684684
rect 25498 684564 25504 684616
rect 25556 684604 25562 684616
rect 449158 684604 449164 684616
rect 25556 684576 449164 684604
rect 25556 684564 25562 684576
rect 449158 684564 449164 684576
rect 449216 684564 449222 684616
rect 6270 684496 6276 684548
rect 6328 684536 6334 684548
rect 436094 684536 436100 684548
rect 6328 684508 436100 684536
rect 6328 684496 6334 684508
rect 436094 684496 436100 684508
rect 436152 684496 436158 684548
rect 221734 684428 221740 684480
rect 221792 684468 221798 684480
rect 543090 684468 543096 684480
rect 221792 684440 543096 684468
rect 221792 684428 221798 684440
rect 543090 684428 543096 684440
rect 543148 684428 543154 684480
rect 38102 684360 38108 684412
rect 38160 684400 38166 684412
rect 361574 684400 361580 684412
rect 38160 684372 361580 684400
rect 38160 684360 38166 684372
rect 361574 684360 361580 684372
rect 361632 684360 361638 684412
rect 398742 684360 398748 684412
rect 398800 684400 398806 684412
rect 405642 684400 405648 684412
rect 398800 684372 405648 684400
rect 398800 684360 398806 684372
rect 405642 684360 405648 684372
rect 405700 684360 405706 684412
rect 418062 684360 418068 684412
rect 418120 684400 418126 684412
rect 424962 684400 424968 684412
rect 418120 684372 424968 684400
rect 418120 684360 418126 684372
rect 424962 684360 424968 684372
rect 425020 684360 425026 684412
rect 437382 684360 437388 684412
rect 437440 684400 437446 684412
rect 444282 684400 444288 684412
rect 437440 684372 444288 684400
rect 437440 684360 437446 684372
rect 444282 684360 444288 684372
rect 444340 684360 444346 684412
rect 456702 684360 456708 684412
rect 456760 684400 456766 684412
rect 463602 684400 463608 684412
rect 456760 684372 463608 684400
rect 456760 684360 456766 684372
rect 463602 684360 463608 684372
rect 463660 684360 463666 684412
rect 33778 684292 33784 684344
rect 33836 684332 33842 684344
rect 365806 684332 365812 684344
rect 33836 684304 365812 684332
rect 33836 684292 33842 684304
rect 365806 684292 365812 684304
rect 365864 684292 365870 684344
rect 365898 684292 365904 684344
rect 365956 684332 365962 684344
rect 580902 684332 580908 684344
rect 365956 684304 580908 684332
rect 365956 684292 365962 684304
rect 580902 684292 580908 684304
rect 580960 684292 580966 684344
rect 208302 684224 208308 684276
rect 208360 684264 208366 684276
rect 542998 684264 543004 684276
rect 208360 684236 543004 684264
rect 208360 684224 208366 684236
rect 542998 684224 543004 684236
rect 543056 684224 543062 684276
rect 38010 684156 38016 684208
rect 38068 684196 38074 684208
rect 374638 684196 374644 684208
rect 38068 684168 374644 684196
rect 38068 684156 38074 684168
rect 374638 684156 374644 684168
rect 374696 684156 374702 684208
rect 379330 684156 379336 684208
rect 379388 684196 379394 684208
rect 386322 684196 386328 684208
rect 379388 684168 386328 684196
rect 379388 684156 379394 684168
rect 386322 684156 386328 684168
rect 386380 684156 386386 684208
rect 476022 684156 476028 684208
rect 476080 684196 476086 684208
rect 482922 684196 482928 684208
rect 476080 684168 482928 684196
rect 476080 684156 476086 684168
rect 482922 684156 482928 684168
rect 482980 684156 482986 684208
rect 195100 684088 195106 684140
rect 195158 684128 195164 684140
rect 541802 684128 541808 684140
rect 195158 684100 541808 684128
rect 195158 684088 195164 684100
rect 541802 684088 541808 684100
rect 541860 684088 541866 684140
rect 39482 684020 39488 684072
rect 39540 684060 39546 684072
rect 387794 684060 387800 684072
rect 39540 684032 387800 684060
rect 39540 684020 39546 684032
rect 387794 684020 387800 684032
rect 387852 684020 387858 684072
rect 495342 684020 495348 684072
rect 495400 684060 495406 684072
rect 497918 684060 497924 684072
rect 495400 684032 497924 684060
rect 495400 684020 495406 684032
rect 497918 684020 497924 684032
rect 497976 684020 497982 684072
rect 39574 683952 39580 684004
rect 39632 683992 39638 684004
rect 392210 683992 392216 684004
rect 39632 683964 392216 683992
rect 39632 683952 39638 683964
rect 392210 683952 392216 683964
rect 392268 683952 392274 684004
rect 37918 683884 37924 683936
rect 37976 683924 37982 683936
rect 400950 683924 400956 683936
rect 37976 683896 400956 683924
rect 37976 683884 37982 683896
rect 400950 683884 400956 683896
rect 401008 683884 401014 683936
rect 5074 683816 5080 683868
rect 5132 683856 5138 683868
rect 379054 683856 379060 683868
rect 5132 683828 379060 683856
rect 5132 683816 5138 683828
rect 379054 683816 379060 683828
rect 379112 683816 379118 683868
rect 379514 683816 379520 683868
rect 379572 683856 379578 683868
rect 580166 683856 580172 683868
rect 379572 683828 580172 683856
rect 379572 683816 379578 683828
rect 580166 683816 580172 683828
rect 580224 683816 580230 683868
rect 32398 683748 32404 683800
rect 32456 683788 32462 683800
rect 427262 683788 427268 683800
rect 32456 683760 427268 683788
rect 32456 683748 32462 683760
rect 427262 683748 427268 683760
rect 427320 683748 427326 683800
rect 142798 683680 142804 683732
rect 142856 683720 142862 683732
rect 539134 683720 539140 683732
rect 142856 683692 539140 683720
rect 142856 683680 142862 683692
rect 539134 683680 539140 683692
rect 539192 683680 539198 683732
rect 182082 683612 182088 683664
rect 182140 683652 182146 683664
rect 579890 683652 579896 683664
rect 182140 683624 579896 683652
rect 182140 683612 182146 683624
rect 579890 683612 579896 683624
rect 579948 683612 579954 683664
rect 138382 683544 138388 683596
rect 138440 683584 138446 683596
rect 539226 683584 539232 683596
rect 138440 683556 539232 683584
rect 138440 683544 138446 683556
rect 539226 683544 539232 683556
rect 539284 683544 539290 683596
rect 2958 683476 2964 683528
rect 3016 683516 3022 683528
rect 431862 683516 431868 683528
rect 3016 683488 431868 683516
rect 3016 683476 3022 683488
rect 431862 683476 431868 683488
rect 431920 683476 431926 683528
rect 29638 683408 29644 683460
rect 29696 683448 29702 683460
rect 466730 683448 466736 683460
rect 29696 683420 466736 683448
rect 29696 683408 29702 683420
rect 466730 683408 466736 683420
rect 466788 683408 466794 683460
rect 3142 683340 3148 683392
rect 3200 683380 3206 683392
rect 458174 683380 458180 683392
rect 3200 683352 458180 683380
rect 3200 683340 3206 683352
rect 458174 683340 458180 683352
rect 458232 683340 458238 683392
rect 4890 683272 4896 683324
rect 4948 683312 4954 683324
rect 475470 683312 475476 683324
rect 4948 683284 475476 683312
rect 4948 683272 4954 683284
rect 475470 683272 475476 683284
rect 475528 683272 475534 683324
rect 521654 683272 521660 683324
rect 521712 683312 521718 683324
rect 523770 683312 523776 683324
rect 521712 683284 523776 683312
rect 521712 683272 521718 683284
rect 523770 683272 523776 683284
rect 523828 683272 523834 683324
rect 89852 683204 89858 683256
rect 89910 683204 89916 683256
rect 98592 683204 98598 683256
rect 98650 683244 98656 683256
rect 580718 683244 580724 683256
rect 98650 683216 580724 683244
rect 98650 683204 98656 683216
rect 580718 683204 580724 683216
rect 580776 683204 580782 683256
rect 89870 683176 89898 683204
rect 580534 683176 580540 683188
rect 89870 683148 580540 683176
rect 580534 683136 580540 683148
rect 580592 683136 580598 683188
rect 2774 682252 2780 682304
rect 2832 682292 2838 682304
rect 5534 682292 5540 682304
rect 2832 682264 5540 682292
rect 2832 682252 2838 682264
rect 5534 682252 5540 682264
rect 5592 682252 5598 682304
rect 540882 674772 540888 674824
rect 540940 674812 540946 674824
rect 579706 674812 579712 674824
rect 540940 674784 579712 674812
rect 540940 674772 540946 674784
rect 579706 674772 579712 674784
rect 579764 674772 579770 674824
rect 2774 669264 2780 669316
rect 2832 669304 2838 669316
rect 33778 669304 33784 669316
rect 2832 669276 33784 669304
rect 2832 669264 2838 669276
rect 33778 669264 33784 669276
rect 33836 669264 33842 669316
rect 2774 654032 2780 654084
rect 2832 654072 2838 654084
rect 38102 654072 38108 654084
rect 2832 654044 38108 654072
rect 2832 654032 2838 654044
rect 38102 654032 38108 654044
rect 38160 654032 38166 654084
rect 578142 651312 578148 651364
rect 578200 651352 578206 651364
rect 579614 651352 579620 651364
rect 578200 651324 579620 651352
rect 578200 651312 578206 651324
rect 579614 651312 579620 651324
rect 579672 651312 579678 651364
rect 543090 640228 543096 640280
rect 543148 640268 543154 640280
rect 579706 640268 579712 640280
rect 543148 640240 579712 640268
rect 543148 640228 543154 640240
rect 579706 640228 579712 640240
rect 579764 640228 579770 640280
rect 540698 627852 540704 627904
rect 540756 627892 540762 627904
rect 579706 627892 579712 627904
rect 540756 627864 579712 627892
rect 540756 627852 540762 627864
rect 579706 627852 579712 627864
rect 579764 627852 579770 627904
rect 2774 624860 2780 624912
rect 2832 624900 2838 624912
rect 6730 624900 6736 624912
rect 2832 624872 6736 624900
rect 2832 624860 2838 624872
rect 6730 624860 6736 624872
rect 6788 624860 6794 624912
rect 2774 610444 2780 610496
rect 2832 610484 2838 610496
rect 5074 610484 5080 610496
rect 2832 610456 5080 610484
rect 2832 610444 2838 610456
rect 5074 610444 5080 610456
rect 5132 610444 5138 610496
rect 578050 604392 578056 604444
rect 578108 604432 578114 604444
rect 579614 604432 579620 604444
rect 578108 604404 579620 604432
rect 578108 604392 578114 604404
rect 579614 604392 579620 604404
rect 579672 604392 579678 604444
rect 2774 596096 2780 596148
rect 2832 596136 2838 596148
rect 38010 596136 38016 596148
rect 2832 596108 38016 596136
rect 2832 596096 2838 596108
rect 38010 596096 38016 596108
rect 38068 596096 38074 596148
rect 542998 593308 543004 593360
rect 543056 593348 543062 593360
rect 579706 593348 579712 593360
rect 543056 593320 579712 593348
rect 543056 593308 543062 593320
rect 579706 593308 579712 593320
rect 579764 593308 579770 593360
rect 540514 580932 540520 580984
rect 540572 580972 540578 580984
rect 579706 580972 579712 580984
rect 540572 580944 579712 580972
rect 540572 580932 540578 580944
rect 579706 580932 579712 580944
rect 579764 580932 579770 580984
rect 2774 567332 2780 567384
rect 2832 567372 2838 567384
rect 6638 567372 6644 567384
rect 2832 567344 6644 567372
rect 2832 567332 2838 567344
rect 6638 567332 6644 567344
rect 6696 567332 6702 567384
rect 577958 557336 577964 557388
rect 578016 557376 578022 557388
rect 579614 557376 579620 557388
rect 578016 557348 579620 557376
rect 578016 557336 578022 557348
rect 579614 557336 579620 557348
rect 579672 557336 579678 557388
rect 2774 553324 2780 553376
rect 2832 553364 2838 553376
rect 39574 553364 39580 553376
rect 2832 553336 39580 553364
rect 2832 553324 2838 553336
rect 39574 553324 39580 553336
rect 39632 553324 39638 553376
rect 541802 546388 541808 546440
rect 541860 546428 541866 546440
rect 579706 546428 579712 546440
rect 541860 546400 579712 546428
rect 541860 546388 541866 546400
rect 579706 546388 579712 546400
rect 579764 546388 579770 546440
rect 2774 539520 2780 539572
rect 2832 539560 2838 539572
rect 39482 539560 39488 539572
rect 2832 539532 39488 539560
rect 2832 539520 2838 539532
rect 39482 539520 39488 539532
rect 39540 539520 39546 539572
rect 539502 534012 539508 534064
rect 539560 534052 539566 534064
rect 579706 534052 579712 534064
rect 539560 534024 579712 534052
rect 539560 534012 539566 534024
rect 579706 534012 579712 534024
rect 579764 534012 579770 534064
rect 2774 509940 2780 509992
rect 2832 509980 2838 509992
rect 6546 509980 6552 509992
rect 2832 509952 6552 509980
rect 2832 509940 2838 509952
rect 6546 509940 6552 509952
rect 6604 509940 6610 509992
rect 539410 487092 539416 487144
rect 539468 487132 539474 487144
rect 579890 487132 579896 487144
rect 539468 487104 579896 487132
rect 539468 487092 539474 487104
rect 579890 487092 579896 487104
rect 579948 487092 579954 487144
rect 2866 481584 2872 481636
rect 2924 481624 2930 481636
rect 37918 481624 37924 481636
rect 2924 481596 37924 481624
rect 2924 481584 2930 481596
rect 37918 481584 37924 481596
rect 37976 481584 37982 481636
rect 540330 463632 540336 463684
rect 540388 463672 540394 463684
rect 579890 463672 579896 463684
rect 540388 463644 579896 463672
rect 540388 463632 540394 463644
rect 579890 463632 579896 463644
rect 579948 463632 579954 463684
rect 539318 452548 539324 452600
rect 539376 452588 539382 452600
rect 579890 452588 579896 452600
rect 539376 452560 579896 452588
rect 539376 452548 539382 452560
rect 579890 452548 579896 452560
rect 579948 452548 579954 452600
rect 2866 452412 2872 452464
rect 2924 452452 2930 452464
rect 6454 452452 6460 452464
rect 2924 452424 6460 452452
rect 2924 452412 2930 452424
rect 6454 452412 6460 452424
rect 6512 452412 6518 452464
rect 577866 440172 577872 440224
rect 577924 440212 577930 440224
rect 579890 440212 579896 440224
rect 577924 440184 579896 440212
rect 577924 440172 577930 440184
rect 579890 440172 579896 440184
rect 579948 440172 579954 440224
rect 2774 438676 2780 438728
rect 2832 438716 2838 438728
rect 4982 438716 4988 438728
rect 2832 438688 4988 438716
rect 2832 438676 2838 438688
rect 4982 438676 4988 438688
rect 5040 438676 5046 438728
rect 2866 425008 2872 425060
rect 2924 425048 2930 425060
rect 25590 425048 25596 425060
rect 2924 425020 25596 425048
rect 2924 425008 2930 425020
rect 25590 425008 25596 425020
rect 25648 425008 25654 425060
rect 541710 405628 541716 405680
rect 541768 405668 541774 405680
rect 579982 405668 579988 405680
rect 541768 405640 579988 405668
rect 541768 405628 541774 405640
rect 579982 405628 579988 405640
rect 580040 405628 580046 405680
rect 2866 395020 2872 395072
rect 2924 395060 2930 395072
rect 6362 395060 6368 395072
rect 2924 395032 6368 395060
rect 2924 395020 2930 395032
rect 6362 395020 6368 395032
rect 6420 395020 6426 395072
rect 541618 393252 541624 393304
rect 541676 393292 541682 393304
rect 579982 393292 579988 393304
rect 541676 393264 579988 393292
rect 541676 393252 541682 393264
rect 579982 393252 579988 393264
rect 580040 393252 580046 393304
rect 539226 369792 539232 369844
rect 539284 369832 539290 369844
rect 579982 369832 579988 369844
rect 539284 369804 579988 369832
rect 539284 369792 539290 369804
rect 579982 369792 579988 369804
rect 580040 369792 580046 369844
rect 2958 367004 2964 367056
rect 3016 367044 3022 367056
rect 32398 367044 32404 367056
rect 3016 367016 32404 367044
rect 3016 367004 3022 367016
rect 32398 367004 32404 367016
rect 32456 367004 32462 367056
rect 539134 358708 539140 358760
rect 539192 358748 539198 358760
rect 579982 358748 579988 358760
rect 539192 358720 579988 358748
rect 539192 358708 539198 358720
rect 579982 358708 579988 358720
rect 580040 358708 580046 358760
rect 577774 346332 577780 346384
rect 577832 346372 577838 346384
rect 579890 346372 579896 346384
rect 577832 346344 579896 346372
rect 577832 346332 577838 346344
rect 579890 346332 579896 346344
rect 579948 346332 579954 346384
rect 2958 337560 2964 337612
rect 3016 337600 3022 337612
rect 6270 337600 6276 337612
rect 3016 337572 6276 337600
rect 3016 337560 3022 337572
rect 6270 337560 6276 337572
rect 6328 337560 6334 337612
rect 2958 323076 2964 323128
rect 3016 323116 3022 323128
rect 7558 323116 7564 323128
rect 3016 323088 7564 323116
rect 3016 323076 3022 323088
rect 7558 323076 7564 323088
rect 7616 323076 7622 323128
rect 539042 311788 539048 311840
rect 539100 311828 539106 311840
rect 580166 311828 580172 311840
rect 539100 311800 580172 311828
rect 539100 311788 539106 311800
rect 580166 311788 580172 311800
rect 580224 311788 580230 311840
rect 540790 299412 540796 299464
rect 540848 299452 540854 299464
rect 580166 299452 580172 299464
rect 540848 299424 580172 299452
rect 540848 299412 540854 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 3050 295264 3056 295316
rect 3108 295304 3114 295316
rect 25498 295304 25504 295316
rect 3108 295276 25504 295304
rect 3108 295264 3114 295276
rect 25498 295264 25504 295276
rect 25556 295264 25562 295316
rect 538950 264868 538956 264920
rect 539008 264908 539014 264920
rect 580166 264908 580172 264920
rect 539008 264880 580172 264908
rect 539008 264868 539014 264880
rect 580166 264868 580172 264880
rect 580224 264868 580230 264920
rect 577682 252492 577688 252544
rect 577740 252532 577746 252544
rect 579982 252532 579988 252544
rect 577740 252504 579988 252532
rect 577740 252492 577746 252504
rect 579982 252492 579988 252504
rect 580040 252492 580046 252544
rect 3142 251268 3148 251320
rect 3200 251308 3206 251320
rect 6178 251308 6184 251320
rect 3200 251280 6184 251308
rect 3200 251268 3206 251280
rect 6178 251268 6184 251280
rect 6236 251268 6242 251320
rect 3326 223524 3332 223576
rect 3384 223564 3390 223576
rect 29638 223564 29644 223576
rect 3384 223536 29644 223564
rect 3384 223524 3390 223536
rect 29638 223524 29644 223536
rect 29696 223524 29702 223576
rect 538858 217948 538864 218000
rect 538916 217988 538922 218000
rect 580166 217988 580172 218000
rect 538916 217960 580172 217988
rect 538916 217948 538922 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 2774 208156 2780 208208
rect 2832 208196 2838 208208
rect 4890 208196 4896 208208
rect 2832 208168 4896 208196
rect 2832 208156 2838 208168
rect 4890 208156 4896 208168
rect 4948 208156 4954 208208
rect 577590 205572 577596 205624
rect 577648 205612 577654 205624
rect 580718 205612 580724 205624
rect 577648 205584 580724 205612
rect 577648 205572 577654 205584
rect 580718 205572 580724 205584
rect 580776 205572 580782 205624
rect 2774 179460 2780 179512
rect 2832 179500 2838 179512
rect 4798 179500 4804 179512
rect 2832 179472 4804 179500
rect 2832 179460 2838 179472
rect 4798 179460 4804 179472
rect 4856 179460 4862 179512
rect 3142 165520 3148 165572
rect 3200 165560 3206 165572
rect 39390 165560 39396 165572
rect 3200 165532 39396 165560
rect 3200 165520 3206 165532
rect 39390 165520 39396 165532
rect 39448 165520 39454 165572
rect 540606 158652 540612 158704
rect 540664 158692 540670 158704
rect 580166 158692 580172 158704
rect 540664 158664 580172 158692
rect 540664 158652 540670 158664
rect 580166 158652 580172 158664
rect 580224 158652 580230 158704
rect 3326 136552 3332 136604
rect 3384 136592 3390 136604
rect 22738 136592 22744 136604
rect 3384 136564 22744 136592
rect 3384 136552 3390 136564
rect 22738 136552 22744 136564
rect 22796 136552 22802 136604
rect 3326 122748 3332 122800
rect 3384 122788 3390 122800
rect 24118 122788 24124 122800
rect 3384 122760 24124 122788
rect 3384 122748 3390 122760
rect 24118 122748 24124 122760
rect 24176 122748 24182 122800
rect 540422 111732 540428 111784
rect 540480 111772 540486 111784
rect 580166 111772 580172 111784
rect 540480 111744 580172 111772
rect 540480 111732 540486 111744
rect 580166 111732 580172 111744
rect 580224 111732 580230 111784
rect 3326 79976 3332 80028
rect 3384 80016 3390 80028
rect 39298 80016 39304 80028
rect 3384 79988 39304 80016
rect 3384 79976 3390 79988
rect 39298 79976 39304 79988
rect 39356 79976 39362 80028
rect 540238 64812 540244 64864
rect 540296 64852 540302 64864
rect 580166 64852 580172 64864
rect 540296 64824 580172 64852
rect 540296 64812 540302 64824
rect 580166 64812 580172 64824
rect 580224 64812 580230 64864
rect 26142 62024 26148 62076
rect 26200 62064 26206 62076
rect 61010 62064 61016 62076
rect 26200 62036 61016 62064
rect 26200 62024 26206 62036
rect 61010 62024 61016 62036
rect 61068 62024 61074 62076
rect 64782 62024 64788 62076
rect 64840 62064 64846 62076
rect 93854 62064 93860 62076
rect 64840 62036 93860 62064
rect 64840 62024 64846 62036
rect 93854 62024 93860 62036
rect 93912 62024 93918 62076
rect 107470 62024 107476 62076
rect 107528 62064 107534 62076
rect 131482 62064 131488 62076
rect 107528 62036 131488 62064
rect 107528 62024 107534 62036
rect 131482 62024 131488 62036
rect 131540 62024 131546 62076
rect 132402 62024 132408 62076
rect 132460 62064 132466 62076
rect 151906 62064 151912 62076
rect 132460 62036 151912 62064
rect 132460 62024 132466 62036
rect 151906 62024 151912 62036
rect 151964 62024 151970 62076
rect 153102 62024 153108 62076
rect 153160 62064 153166 62076
rect 170214 62064 170220 62076
rect 153160 62036 170220 62064
rect 153160 62024 153166 62036
rect 170214 62024 170220 62036
rect 170272 62024 170278 62076
rect 171042 62024 171048 62076
rect 171100 62064 171106 62076
rect 185578 62064 185584 62076
rect 171100 62036 185584 62064
rect 171100 62024 171106 62036
rect 185578 62024 185584 62036
rect 185636 62024 185642 62076
rect 198642 62024 198648 62076
rect 198700 62064 198706 62076
rect 209038 62064 209044 62076
rect 198700 62036 209044 62064
rect 198700 62024 198706 62036
rect 209038 62024 209044 62036
rect 209096 62024 209102 62076
rect 517790 62024 517796 62076
rect 517848 62064 517854 62076
rect 518802 62064 518808 62076
rect 517848 62036 518808 62064
rect 517848 62024 517854 62036
rect 518802 62024 518808 62036
rect 518860 62024 518866 62076
rect 521930 62024 521936 62076
rect 521988 62064 521994 62076
rect 522850 62064 522856 62076
rect 521988 62036 522856 62064
rect 521988 62024 521994 62036
rect 522850 62024 522856 62036
rect 522908 62024 522914 62076
rect 24762 61956 24768 62008
rect 24820 61996 24826 62008
rect 59998 61996 60004 62008
rect 24820 61968 60004 61996
rect 24820 61956 24826 61968
rect 59998 61956 60004 61968
rect 60056 61956 60062 62008
rect 60642 61956 60648 62008
rect 60700 61996 60706 62008
rect 90634 61996 90640 62008
rect 60700 61968 90640 61996
rect 60700 61956 60706 61968
rect 90634 61956 90640 61968
rect 90692 61956 90698 62008
rect 96522 61956 96528 62008
rect 96580 61996 96586 62008
rect 121454 61996 121460 62008
rect 96580 61968 121460 61996
rect 96580 61956 96586 61968
rect 121454 61956 121460 61968
rect 121512 61956 121518 62008
rect 124122 61956 124128 62008
rect 124180 61996 124186 62008
rect 144914 61996 144920 62008
rect 124180 61968 144920 61996
rect 124180 61956 124186 61968
rect 144914 61956 144920 61968
rect 144972 61956 144978 62008
rect 146202 61956 146208 62008
rect 146260 61996 146266 62008
rect 164234 61996 164240 62008
rect 146260 61968 164240 61996
rect 146260 61956 146266 61968
rect 164234 61956 164240 61968
rect 164292 61956 164298 62008
rect 168282 61956 168288 62008
rect 168340 61996 168346 62008
rect 183554 61996 183560 62008
rect 168340 61968 183560 61996
rect 168340 61956 168346 61968
rect 183554 61956 183560 61968
rect 183612 61956 183618 62008
rect 186222 61956 186228 62008
rect 186280 61996 186286 62008
rect 198826 61996 198832 62008
rect 186280 61968 198832 61996
rect 186280 61956 186286 61968
rect 198826 61956 198832 61968
rect 198884 61956 198890 62008
rect 202690 61956 202696 62008
rect 202748 61996 202754 62008
rect 212074 61996 212080 62008
rect 202748 61968 212080 61996
rect 202748 61956 202754 61968
rect 212074 61956 212080 61968
rect 212132 61956 212138 62008
rect 216582 61956 216588 62008
rect 216640 61996 216646 62008
rect 224310 61996 224316 62008
rect 216640 61968 224316 61996
rect 216640 61956 216646 61968
rect 224310 61956 224316 61968
rect 224368 61956 224374 62008
rect 475010 61956 475016 62008
rect 475068 61996 475074 62008
rect 496078 61996 496084 62008
rect 475068 61968 496084 61996
rect 475068 61956 475074 61968
rect 496078 61956 496084 61968
rect 496136 61956 496142 62008
rect 516778 61956 516784 62008
rect 516836 61996 516842 62008
rect 519538 61996 519544 62008
rect 516836 61968 519544 61996
rect 516836 61956 516842 61968
rect 519538 61956 519544 61968
rect 519596 61956 519602 62008
rect 524966 61956 524972 62008
rect 525024 61996 525030 62008
rect 531958 61996 531964 62008
rect 525024 61968 531964 61996
rect 525024 61956 525030 61968
rect 531958 61956 531964 61968
rect 532016 61956 532022 62008
rect 19242 61888 19248 61940
rect 19300 61928 19306 61940
rect 55306 61928 55312 61940
rect 19300 61900 55312 61928
rect 19300 61888 19306 61900
rect 55306 61888 55312 61900
rect 55364 61888 55370 61940
rect 59906 61888 59912 61940
rect 59964 61928 59970 61940
rect 67174 61928 67180 61940
rect 59964 61900 67180 61928
rect 59964 61888 59970 61900
rect 67174 61888 67180 61900
rect 67232 61888 67238 61940
rect 68922 61888 68928 61940
rect 68980 61928 68986 61940
rect 97994 61928 98000 61940
rect 68980 61900 98000 61928
rect 68980 61888 68986 61900
rect 97994 61888 98000 61900
rect 98052 61888 98058 61940
rect 99282 61888 99288 61940
rect 99340 61928 99346 61940
rect 124306 61928 124312 61940
rect 99340 61900 124312 61928
rect 99340 61888 99346 61900
rect 124306 61888 124312 61900
rect 124364 61888 124370 61940
rect 133782 61888 133788 61940
rect 133840 61928 133846 61940
rect 153930 61928 153936 61940
rect 133840 61900 153936 61928
rect 133840 61888 133846 61900
rect 153930 61888 153936 61900
rect 153988 61888 153994 61940
rect 158622 61888 158628 61940
rect 158680 61928 158686 61940
rect 174354 61928 174360 61940
rect 158680 61900 174360 61928
rect 158680 61888 158686 61900
rect 174354 61888 174360 61900
rect 174412 61888 174418 61940
rect 175182 61888 175188 61940
rect 175240 61928 175246 61940
rect 188614 61928 188620 61940
rect 175240 61900 188620 61928
rect 175240 61888 175246 61900
rect 188614 61888 188620 61900
rect 188672 61888 188678 61940
rect 197262 61888 197268 61940
rect 197320 61928 197326 61940
rect 208394 61928 208400 61940
rect 197320 61900 208400 61928
rect 197320 61888 197326 61900
rect 208394 61888 208400 61900
rect 208452 61888 208458 61940
rect 209682 61888 209688 61940
rect 209740 61928 209746 61940
rect 218238 61928 218244 61940
rect 209740 61900 218244 61928
rect 209740 61888 209746 61900
rect 218238 61888 218244 61900
rect 218296 61888 218302 61940
rect 229002 61888 229008 61940
rect 229060 61928 229066 61940
rect 235534 61928 235540 61940
rect 229060 61900 235540 61928
rect 229060 61888 229066 61900
rect 235534 61888 235540 61900
rect 235592 61888 235598 61940
rect 423950 61888 423956 61940
rect 424008 61928 424014 61940
rect 447134 61928 447140 61940
rect 424008 61900 447140 61928
rect 424008 61888 424014 61900
rect 447134 61888 447140 61900
rect 447192 61888 447198 61940
rect 484118 61888 484124 61940
rect 484176 61928 484182 61940
rect 512638 61928 512644 61940
rect 484176 61900 512644 61928
rect 484176 61888 484182 61900
rect 512638 61888 512644 61900
rect 512696 61888 512702 61940
rect 515766 61888 515772 61940
rect 515824 61928 515830 61940
rect 522298 61928 522304 61940
rect 515824 61900 522304 61928
rect 515824 61888 515830 61900
rect 522298 61888 522304 61900
rect 522356 61888 522362 61940
rect 23382 61820 23388 61872
rect 23440 61860 23446 61872
rect 59354 61860 59360 61872
rect 23440 61832 59360 61860
rect 23440 61820 23446 61832
rect 59354 61820 59360 61832
rect 59412 61820 59418 61872
rect 62022 61820 62028 61872
rect 62080 61860 62086 61872
rect 91646 61860 91652 61872
rect 62080 61832 91652 61860
rect 62080 61820 62086 61832
rect 91646 61820 91652 61832
rect 91704 61820 91710 61872
rect 92382 61820 92388 61872
rect 92440 61860 92446 61872
rect 118234 61860 118240 61872
rect 92440 61832 118240 61860
rect 92440 61820 92446 61832
rect 118234 61820 118240 61832
rect 118292 61820 118298 61872
rect 122742 61820 122748 61872
rect 122800 61860 122806 61872
rect 143718 61860 143724 61872
rect 122800 61832 143724 61860
rect 122800 61820 122806 61832
rect 143718 61820 143724 61832
rect 143776 61820 143782 61872
rect 144822 61820 144828 61872
rect 144880 61860 144886 61872
rect 163130 61860 163136 61872
rect 144880 61832 163136 61860
rect 144880 61820 144886 61832
rect 163130 61820 163136 61832
rect 163188 61820 163194 61872
rect 165522 61820 165528 61872
rect 165580 61860 165586 61872
rect 180794 61860 180800 61872
rect 165580 61832 180800 61860
rect 165580 61820 165586 61832
rect 180794 61820 180800 61832
rect 180852 61820 180858 61872
rect 184842 61820 184848 61872
rect 184900 61860 184906 61872
rect 197814 61860 197820 61872
rect 184900 61832 197820 61860
rect 184900 61820 184906 61832
rect 197814 61820 197820 61832
rect 197872 61820 197878 61872
rect 200022 61820 200028 61872
rect 200080 61860 200086 61872
rect 210050 61860 210056 61872
rect 200080 61832 210056 61860
rect 200080 61820 200086 61832
rect 210050 61820 210056 61832
rect 210108 61820 210114 61872
rect 217962 61820 217968 61872
rect 218020 61860 218026 61872
rect 225322 61860 225328 61872
rect 218020 61832 225328 61860
rect 218020 61820 218026 61832
rect 225322 61820 225328 61832
rect 225380 61820 225386 61872
rect 226242 61820 226248 61872
rect 226300 61860 226306 61872
rect 232498 61860 232504 61872
rect 226300 61832 232504 61860
rect 226300 61820 226306 61832
rect 232498 61820 232504 61832
rect 232556 61820 232562 61872
rect 439222 61820 439228 61872
rect 439280 61860 439286 61872
rect 465166 61860 465172 61872
rect 439280 61832 465172 61860
rect 439280 61820 439286 61832
rect 465166 61820 465172 61832
rect 465224 61820 465230 61872
rect 487062 61820 487068 61872
rect 487120 61860 487126 61872
rect 516870 61860 516876 61872
rect 487120 61832 516876 61860
rect 487120 61820 487126 61832
rect 516870 61820 516876 61832
rect 516928 61820 516934 61872
rect 525702 61820 525708 61872
rect 525760 61860 525766 61872
rect 534718 61860 534724 61872
rect 525760 61832 534724 61860
rect 525760 61820 525766 61832
rect 534718 61820 534724 61832
rect 534776 61820 534782 61872
rect 538030 61820 538036 61872
rect 538088 61860 538094 61872
rect 541618 61860 541624 61872
rect 538088 61832 541624 61860
rect 538088 61820 538094 61832
rect 541618 61820 541624 61832
rect 541676 61820 541682 61872
rect 15102 61752 15108 61804
rect 15160 61792 15166 61804
rect 51902 61792 51908 61804
rect 15160 61764 51908 61792
rect 15160 61752 15166 61764
rect 51902 61752 51908 61764
rect 51960 61752 51966 61804
rect 56502 61752 56508 61804
rect 56560 61792 56566 61804
rect 87598 61792 87604 61804
rect 56560 61764 87604 61792
rect 56560 61752 56566 61764
rect 87598 61752 87604 61764
rect 87656 61752 87662 61804
rect 100662 61752 100668 61804
rect 100720 61792 100726 61804
rect 125686 61792 125692 61804
rect 100720 61764 125692 61792
rect 100720 61752 100726 61764
rect 125686 61752 125692 61764
rect 125744 61752 125750 61804
rect 133690 61752 133696 61804
rect 133748 61792 133754 61804
rect 153286 61792 153292 61804
rect 133748 61764 153292 61792
rect 133748 61752 133754 61764
rect 153286 61752 153292 61764
rect 153344 61752 153350 61804
rect 154482 61752 154488 61804
rect 154540 61792 154546 61804
rect 171318 61792 171324 61804
rect 154540 61764 171324 61792
rect 154540 61752 154546 61764
rect 171318 61752 171324 61764
rect 171376 61752 171382 61804
rect 173802 61752 173808 61804
rect 173860 61792 173866 61804
rect 187694 61792 187700 61804
rect 173860 61764 187700 61792
rect 173860 61752 173866 61764
rect 187694 61752 187700 61764
rect 187752 61752 187758 61804
rect 188982 61752 188988 61804
rect 189040 61792 189046 61804
rect 200850 61792 200856 61804
rect 189040 61764 200856 61792
rect 189040 61752 189046 61764
rect 200850 61752 200856 61764
rect 200908 61752 200914 61804
rect 201402 61752 201408 61804
rect 201460 61792 201466 61804
rect 211154 61792 211160 61804
rect 201460 61764 211160 61792
rect 201460 61752 201466 61764
rect 211154 61752 211160 61764
rect 211212 61752 211218 61804
rect 212442 61752 212448 61804
rect 212500 61792 212506 61804
rect 221274 61792 221280 61804
rect 212500 61764 221280 61792
rect 212500 61752 212506 61764
rect 221274 61752 221280 61764
rect 221332 61752 221338 61804
rect 222102 61752 222108 61804
rect 222160 61792 222166 61804
rect 229462 61792 229468 61804
rect 222160 61764 229468 61792
rect 222160 61752 222166 61764
rect 229462 61752 229468 61764
rect 229520 61752 229526 61804
rect 414750 61752 414756 61804
rect 414808 61792 414814 61804
rect 436186 61792 436192 61804
rect 414808 61764 436192 61792
rect 414808 61752 414814 61764
rect 436186 61752 436192 61764
rect 436244 61752 436250 61804
rect 442350 61752 442356 61804
rect 442408 61792 442414 61804
rect 467926 61792 467932 61804
rect 442408 61764 467932 61792
rect 442408 61752 442414 61764
rect 467926 61752 467932 61764
rect 467984 61752 467990 61804
rect 471882 61752 471888 61804
rect 471940 61792 471946 61804
rect 483658 61792 483664 61804
rect 471940 61764 483664 61792
rect 471940 61752 471946 61764
rect 483658 61752 483664 61764
rect 483716 61752 483722 61804
rect 490282 61752 490288 61804
rect 490340 61792 490346 61804
rect 520826 61792 520832 61804
rect 490340 61764 520832 61792
rect 490340 61752 490346 61764
rect 520826 61752 520832 61764
rect 520884 61752 520890 61804
rect 526990 61752 526996 61804
rect 527048 61792 527054 61804
rect 547230 61792 547236 61804
rect 527048 61764 547236 61792
rect 527048 61752 527054 61764
rect 547230 61752 547236 61764
rect 547288 61752 547294 61804
rect 10962 61684 10968 61736
rect 11020 61724 11026 61736
rect 47762 61724 47768 61736
rect 11020 61696 47768 61724
rect 11020 61684 11026 61696
rect 47762 61684 47768 61696
rect 47820 61684 47826 61736
rect 53742 61684 53748 61736
rect 53800 61724 53806 61736
rect 84562 61724 84568 61736
rect 53800 61696 84568 61724
rect 53800 61684 53806 61696
rect 84562 61684 84568 61696
rect 84620 61684 84626 61736
rect 85482 61684 85488 61736
rect 85540 61724 85546 61736
rect 112070 61724 112076 61736
rect 85540 61696 112076 61724
rect 85540 61684 85546 61696
rect 112070 61684 112076 61696
rect 112128 61684 112134 61736
rect 113082 61684 113088 61736
rect 113140 61724 113146 61736
rect 135530 61724 135536 61736
rect 113140 61696 135536 61724
rect 113140 61684 113146 61696
rect 135530 61684 135536 61696
rect 135588 61684 135594 61736
rect 136542 61684 136548 61736
rect 136600 61724 136606 61736
rect 155954 61724 155960 61736
rect 136600 61696 155960 61724
rect 136600 61684 136606 61696
rect 155954 61684 155960 61696
rect 156012 61684 156018 61736
rect 159910 61684 159916 61736
rect 159968 61724 159974 61736
rect 175366 61724 175372 61736
rect 159968 61696 175372 61724
rect 159968 61684 159974 61696
rect 175366 61684 175372 61696
rect 175424 61684 175430 61736
rect 176470 61684 176476 61736
rect 176528 61724 176534 61736
rect 189626 61724 189632 61736
rect 176528 61696 189632 61724
rect 176528 61684 176534 61696
rect 189626 61684 189632 61696
rect 189684 61684 189690 61736
rect 190362 61684 190368 61736
rect 190420 61724 190426 61736
rect 201862 61724 201868 61736
rect 190420 61696 201868 61724
rect 190420 61684 190426 61696
rect 201862 61684 201868 61696
rect 201920 61684 201926 61736
rect 211062 61684 211068 61736
rect 211120 61724 211126 61736
rect 219434 61724 219440 61736
rect 211120 61696 219440 61724
rect 211120 61684 211126 61696
rect 219434 61684 219440 61696
rect 219492 61684 219498 61736
rect 399478 61684 399484 61736
rect 399536 61724 399542 61736
rect 418246 61724 418252 61736
rect 399536 61696 418252 61724
rect 399536 61684 399542 61696
rect 418246 61684 418252 61696
rect 418304 61684 418310 61736
rect 420822 61684 420828 61736
rect 420880 61724 420886 61736
rect 443178 61724 443184 61736
rect 420880 61696 443184 61724
rect 420880 61684 420886 61696
rect 443178 61684 443184 61696
rect 443236 61684 443242 61736
rect 445386 61684 445392 61736
rect 445444 61724 445450 61736
rect 472066 61724 472072 61736
rect 445444 61696 472072 61724
rect 445444 61684 445450 61696
rect 472066 61684 472072 61696
rect 472124 61684 472130 61736
rect 478046 61684 478052 61736
rect 478104 61724 478110 61736
rect 508498 61724 508504 61736
rect 478104 61696 508504 61724
rect 478104 61684 478110 61696
rect 508498 61684 508504 61696
rect 508556 61684 508562 61736
rect 514662 61684 514668 61736
rect 514720 61724 514726 61736
rect 545758 61724 545764 61736
rect 514720 61696 545764 61724
rect 514720 61684 514726 61696
rect 545758 61684 545764 61696
rect 545816 61684 545822 61736
rect 16482 61616 16488 61668
rect 16540 61656 16546 61668
rect 52914 61656 52920 61668
rect 16540 61628 52920 61656
rect 16540 61616 16546 61628
rect 52914 61616 52920 61628
rect 52972 61616 52978 61668
rect 57882 61616 57888 61668
rect 57940 61656 57946 61668
rect 88610 61656 88616 61668
rect 57940 61628 88616 61656
rect 57940 61616 57946 61628
rect 88610 61616 88616 61628
rect 88668 61616 88674 61668
rect 91002 61616 91008 61668
rect 91060 61656 91066 61668
rect 116118 61656 116124 61668
rect 91060 61628 116124 61656
rect 91060 61616 91066 61628
rect 116118 61616 116124 61628
rect 116176 61616 116182 61668
rect 117222 61616 117228 61668
rect 117280 61656 117286 61668
rect 139670 61656 139676 61668
rect 117280 61628 139676 61656
rect 117280 61616 117286 61628
rect 139670 61616 139676 61628
rect 139728 61616 139734 61668
rect 142062 61616 142068 61668
rect 142120 61656 142126 61668
rect 160094 61656 160100 61668
rect 142120 61628 160100 61656
rect 142120 61616 142126 61628
rect 160094 61616 160100 61628
rect 160152 61616 160158 61668
rect 164142 61616 164148 61668
rect 164200 61656 164206 61668
rect 179414 61656 179420 61668
rect 164200 61628 179420 61656
rect 164200 61616 164206 61628
rect 179414 61616 179420 61628
rect 179472 61616 179478 61668
rect 182082 61616 182088 61668
rect 182140 61656 182146 61668
rect 194686 61656 194692 61668
rect 182140 61628 194692 61656
rect 182140 61616 182146 61628
rect 194686 61616 194692 61628
rect 194744 61616 194750 61668
rect 195882 61616 195888 61668
rect 195940 61656 195946 61668
rect 207014 61656 207020 61668
rect 195940 61628 207020 61656
rect 195940 61616 195946 61628
rect 207014 61616 207020 61628
rect 207072 61616 207078 61668
rect 208302 61616 208308 61668
rect 208360 61656 208366 61668
rect 217134 61656 217140 61668
rect 208360 61628 217140 61656
rect 208360 61616 208366 61628
rect 217134 61616 217140 61628
rect 217192 61616 217198 61668
rect 219250 61616 219256 61668
rect 219308 61656 219314 61668
rect 226334 61656 226340 61668
rect 219308 61628 226340 61656
rect 219308 61616 219314 61628
rect 226334 61616 226340 61628
rect 226392 61616 226398 61668
rect 227622 61616 227628 61668
rect 227680 61656 227686 61668
rect 233510 61656 233516 61668
rect 227680 61628 233516 61656
rect 227680 61616 227686 61628
rect 233510 61616 233516 61628
rect 233568 61616 233574 61668
rect 417786 61616 417792 61668
rect 417844 61656 417850 61668
rect 440326 61656 440332 61668
rect 417844 61628 440332 61656
rect 417844 61616 417850 61628
rect 440326 61616 440332 61628
rect 440384 61616 440390 61668
rect 454586 61616 454592 61668
rect 454644 61656 454650 61668
rect 483014 61656 483020 61668
rect 454644 61628 483020 61656
rect 454644 61616 454650 61628
rect 483014 61616 483020 61628
rect 483072 61616 483078 61668
rect 496446 61616 496452 61668
rect 496504 61656 496510 61668
rect 529198 61656 529204 61668
rect 496504 61628 529204 61656
rect 496504 61616 496510 61628
rect 529198 61616 529204 61628
rect 529256 61616 529262 61668
rect 533154 61616 533160 61668
rect 533212 61656 533218 61668
rect 547138 61656 547144 61668
rect 533212 61628 547144 61656
rect 533212 61616 533218 61628
rect 547138 61616 547144 61628
rect 547196 61616 547202 61668
rect 9582 61548 9588 61600
rect 9640 61588 9646 61600
rect 46934 61588 46940 61600
rect 9640 61560 46940 61588
rect 9640 61548 9646 61560
rect 46934 61548 46940 61560
rect 46992 61548 46998 61600
rect 49602 61548 49608 61600
rect 49660 61588 49666 61600
rect 81434 61588 81440 61600
rect 49660 61560 81440 61588
rect 49660 61548 49666 61560
rect 81434 61548 81440 61560
rect 81492 61548 81498 61600
rect 82630 61548 82636 61600
rect 82688 61588 82694 61600
rect 109126 61588 109132 61600
rect 82688 61560 109132 61588
rect 82688 61548 82694 61560
rect 109126 61548 109132 61560
rect 109184 61548 109190 61600
rect 110322 61548 110328 61600
rect 110380 61588 110386 61600
rect 133874 61588 133880 61600
rect 110380 61560 133880 61588
rect 110380 61548 110386 61560
rect 133874 61548 133880 61560
rect 133932 61548 133938 61600
rect 135162 61548 135168 61600
rect 135220 61588 135226 61600
rect 154942 61588 154948 61600
rect 135220 61560 154948 61588
rect 135220 61548 135226 61560
rect 154942 61548 154948 61560
rect 155000 61548 155006 61600
rect 155862 61548 155868 61600
rect 155920 61588 155926 61600
rect 172606 61588 172612 61600
rect 155920 61560 172612 61588
rect 155920 61548 155926 61560
rect 172606 61548 172612 61560
rect 172664 61548 172670 61600
rect 176562 61548 176568 61600
rect 176620 61588 176626 61600
rect 190730 61588 190736 61600
rect 176620 61560 190736 61588
rect 176620 61548 176626 61560
rect 190730 61548 190736 61560
rect 190788 61548 190794 61600
rect 191742 61548 191748 61600
rect 191800 61588 191806 61600
rect 202874 61588 202880 61600
rect 191800 61560 202880 61588
rect 191800 61548 191806 61560
rect 202874 61548 202880 61560
rect 202932 61548 202938 61600
rect 204162 61548 204168 61600
rect 204220 61588 204226 61600
rect 214098 61588 214104 61600
rect 204220 61560 214104 61588
rect 204220 61548 204226 61560
rect 214098 61548 214104 61560
rect 214156 61548 214162 61600
rect 215202 61548 215208 61600
rect 215260 61588 215266 61600
rect 223666 61588 223672 61600
rect 215260 61560 223672 61588
rect 215260 61548 215266 61560
rect 223666 61548 223672 61560
rect 223724 61548 223730 61600
rect 238662 61548 238668 61600
rect 238720 61588 238726 61600
rect 243722 61588 243728 61600
rect 238720 61560 243728 61588
rect 238720 61548 238726 61560
rect 243722 61548 243728 61560
rect 243780 61548 243786 61600
rect 402514 61548 402520 61600
rect 402572 61588 402578 61600
rect 422386 61588 422392 61600
rect 402572 61560 422392 61588
rect 402572 61548 402578 61560
rect 422386 61548 422392 61560
rect 422444 61548 422450 61600
rect 430114 61548 430120 61600
rect 430172 61588 430178 61600
rect 454218 61588 454224 61600
rect 430172 61560 454224 61588
rect 430172 61548 430178 61560
rect 454218 61548 454224 61560
rect 454276 61548 454282 61600
rect 457622 61548 457628 61600
rect 457680 61588 457686 61600
rect 485866 61588 485872 61600
rect 457680 61560 485872 61588
rect 457680 61548 457686 61560
rect 485866 61548 485872 61560
rect 485924 61548 485930 61600
rect 491202 61548 491208 61600
rect 491260 61588 491266 61600
rect 525794 61588 525800 61600
rect 491260 61560 525800 61588
rect 491260 61548 491266 61560
rect 525794 61548 525800 61560
rect 525852 61548 525858 61600
rect 537202 61548 537208 61600
rect 537260 61588 537266 61600
rect 567838 61588 567844 61600
rect 537260 61560 567844 61588
rect 537260 61548 537266 61560
rect 567838 61548 567844 61560
rect 567896 61548 567902 61600
rect 13630 61480 13636 61532
rect 13688 61520 13694 61532
rect 51074 61520 51080 61532
rect 13688 61492 51080 61520
rect 13688 61480 13694 61492
rect 51074 61480 51080 61492
rect 51132 61480 51138 61532
rect 55122 61480 55128 61532
rect 55180 61520 55186 61532
rect 85574 61520 85580 61532
rect 55180 61492 85580 61520
rect 55180 61480 55186 61492
rect 85574 61480 85580 61492
rect 85632 61480 85638 61532
rect 93762 61480 93768 61532
rect 93820 61520 93826 61532
rect 119246 61520 119252 61532
rect 93820 61492 119252 61520
rect 93820 61480 93826 61492
rect 119246 61480 119252 61492
rect 119304 61480 119310 61532
rect 125410 61480 125416 61532
rect 125468 61520 125474 61532
rect 146754 61520 146760 61532
rect 125468 61492 146760 61520
rect 125468 61480 125474 61492
rect 146754 61480 146760 61492
rect 146812 61480 146818 61532
rect 151630 61480 151636 61532
rect 151688 61520 151694 61532
rect 169202 61520 169208 61532
rect 151688 61492 169208 61520
rect 151688 61480 151694 61492
rect 169202 61480 169208 61492
rect 169260 61480 169266 61532
rect 169662 61480 169668 61532
rect 169720 61520 169726 61532
rect 184934 61520 184940 61532
rect 169720 61492 184940 61520
rect 169720 61480 169726 61492
rect 184934 61480 184940 61492
rect 184992 61480 184998 61532
rect 187602 61480 187608 61532
rect 187660 61520 187666 61532
rect 200206 61520 200212 61532
rect 187660 61492 200212 61520
rect 187660 61480 187666 61492
rect 200206 61480 200212 61492
rect 200264 61480 200270 61532
rect 202782 61480 202788 61532
rect 202840 61520 202846 61532
rect 213086 61520 213092 61532
rect 202840 61492 213092 61520
rect 202840 61480 202846 61492
rect 213086 61480 213092 61492
rect 213144 61480 213150 61532
rect 213822 61480 213828 61532
rect 213880 61520 213886 61532
rect 222286 61520 222292 61532
rect 213880 61492 222292 61520
rect 213880 61480 213886 61492
rect 222286 61480 222292 61492
rect 222344 61480 222350 61532
rect 224862 61480 224868 61532
rect 224920 61520 224926 61532
rect 231854 61520 231860 61532
rect 224920 61492 231860 61520
rect 224920 61480 224926 61492
rect 231854 61480 231860 61492
rect 231912 61480 231918 61532
rect 246942 61480 246948 61532
rect 247000 61520 247006 61532
rect 251266 61520 251272 61532
rect 247000 61492 251272 61520
rect 247000 61480 247006 61492
rect 251266 61480 251272 61492
rect 251324 61480 251330 61532
rect 411714 61480 411720 61532
rect 411772 61520 411778 61532
rect 433426 61520 433432 61532
rect 411772 61492 433432 61520
rect 411772 61480 411778 61492
rect 433426 61480 433432 61492
rect 433484 61480 433490 61532
rect 436002 61480 436008 61532
rect 436060 61520 436066 61532
rect 461026 61520 461032 61532
rect 436060 61492 461032 61520
rect 436060 61480 436066 61492
rect 461026 61480 461032 61492
rect 461084 61480 461090 61532
rect 466822 61480 466828 61532
rect 466880 61520 466886 61532
rect 496814 61520 496820 61532
rect 466880 61492 496820 61520
rect 466880 61480 466886 61492
rect 496814 61480 496820 61492
rect 496872 61480 496878 61532
rect 508682 61480 508688 61532
rect 508740 61520 508746 61532
rect 544378 61520 544384 61532
rect 508740 61492 544384 61520
rect 508740 61480 508746 61492
rect 544378 61480 544384 61492
rect 544436 61480 544442 61532
rect 6822 61412 6828 61464
rect 6880 61452 6886 61464
rect 44726 61452 44732 61464
rect 6880 61424 44732 61452
rect 6880 61412 6886 61424
rect 44726 61412 44732 61424
rect 44784 61412 44790 61464
rect 46842 61412 46848 61464
rect 46900 61452 46906 61464
rect 74534 61452 74540 61464
rect 46900 61424 74540 61452
rect 46900 61412 46906 61424
rect 74534 61412 74540 61424
rect 74592 61412 74598 61464
rect 76558 61412 76564 61464
rect 76616 61452 76622 61464
rect 79410 61452 79416 61464
rect 76616 61424 79416 61452
rect 76616 61412 76622 61424
rect 79410 61412 79416 61424
rect 79468 61412 79474 61464
rect 82722 61412 82728 61464
rect 82780 61452 82786 61464
rect 110414 61452 110420 61464
rect 82780 61424 110420 61452
rect 82780 61412 82786 61424
rect 110414 61412 110420 61424
rect 110472 61412 110478 61464
rect 111702 61412 111708 61464
rect 111760 61452 111766 61464
rect 134518 61452 134524 61464
rect 111760 61424 134524 61452
rect 111760 61412 111766 61424
rect 134518 61412 134524 61424
rect 134576 61412 134582 61464
rect 137922 61412 137928 61464
rect 137980 61452 137986 61464
rect 157334 61452 157340 61464
rect 137980 61424 157340 61452
rect 137980 61412 137986 61424
rect 157334 61412 157340 61424
rect 157392 61412 157398 61464
rect 160002 61412 160008 61464
rect 160060 61452 160066 61464
rect 176746 61452 176752 61464
rect 160060 61424 176752 61452
rect 160060 61412 160066 61424
rect 176746 61412 176752 61424
rect 176804 61412 176810 61464
rect 177942 61412 177948 61464
rect 178000 61452 178006 61464
rect 191834 61452 191840 61464
rect 178000 61424 191840 61452
rect 178000 61412 178006 61424
rect 191834 61412 191840 61424
rect 191892 61412 191898 61464
rect 193122 61412 193128 61464
rect 193180 61452 193186 61464
rect 204254 61452 204260 61464
rect 193180 61424 204260 61452
rect 193180 61412 193186 61424
rect 204254 61412 204260 61424
rect 204312 61412 204318 61464
rect 205542 61412 205548 61464
rect 205600 61452 205606 61464
rect 215294 61452 215300 61464
rect 205600 61424 215300 61452
rect 205600 61412 205606 61424
rect 215294 61412 215300 61424
rect 215352 61412 215358 61464
rect 219342 61412 219348 61464
rect 219400 61452 219406 61464
rect 227714 61452 227720 61464
rect 219400 61424 227720 61452
rect 219400 61412 219406 61424
rect 227714 61412 227720 61424
rect 227772 61412 227778 61464
rect 228910 61412 228916 61464
rect 228968 61452 228974 61464
rect 234614 61452 234620 61464
rect 228968 61424 234620 61452
rect 228968 61412 228974 61424
rect 234614 61412 234620 61424
rect 234672 61412 234678 61464
rect 237282 61412 237288 61464
rect 237340 61452 237346 61464
rect 241698 61452 241704 61464
rect 237340 61424 241704 61452
rect 237340 61412 237346 61424
rect 241698 61412 241704 61424
rect 241756 61412 241762 61464
rect 405550 61412 405556 61464
rect 405608 61452 405614 61464
rect 425146 61452 425152 61464
rect 405608 61424 425152 61452
rect 405608 61412 405614 61424
rect 425146 61412 425152 61424
rect 425204 61412 425210 61464
rect 426986 61412 426992 61464
rect 427044 61452 427050 61464
rect 451458 61452 451464 61464
rect 427044 61424 451464 61452
rect 427044 61412 427050 61424
rect 451458 61412 451464 61424
rect 451516 61412 451522 61464
rect 460658 61412 460664 61464
rect 460716 61452 460722 61464
rect 489914 61452 489920 61464
rect 460716 61424 489920 61452
rect 460716 61412 460722 61424
rect 489914 61412 489920 61424
rect 489972 61412 489978 61464
rect 505554 61412 505560 61464
rect 505612 61452 505618 61464
rect 542354 61452 542360 61464
rect 505612 61424 542360 61452
rect 505612 61412 505618 61424
rect 542354 61412 542360 61424
rect 542412 61412 542418 61464
rect 4062 61344 4068 61396
rect 4120 61384 4126 61396
rect 42794 61384 42800 61396
rect 4120 61356 42800 61384
rect 4120 61344 4126 61356
rect 42794 61344 42800 61356
rect 42852 61344 42858 61396
rect 43438 61344 43444 61396
rect 43496 61384 43502 61396
rect 48774 61384 48780 61396
rect 43496 61356 48780 61384
rect 43496 61344 43502 61356
rect 48774 61344 48780 61356
rect 48832 61344 48838 61396
rect 50982 61344 50988 61396
rect 51040 61384 51046 61396
rect 82814 61384 82820 61396
rect 51040 61356 82820 61384
rect 51040 61344 51046 61356
rect 82814 61344 82820 61356
rect 82872 61344 82878 61396
rect 86862 61344 86868 61396
rect 86920 61384 86926 61396
rect 113174 61384 113180 61396
rect 86920 61356 113180 61384
rect 86920 61344 86926 61356
rect 113174 61344 113180 61356
rect 113232 61344 113238 61396
rect 118602 61344 118608 61396
rect 118660 61384 118666 61396
rect 140774 61384 140780 61396
rect 118660 61356 140780 61384
rect 118660 61344 118666 61356
rect 140774 61344 140780 61356
rect 140832 61344 140838 61396
rect 141970 61344 141976 61396
rect 142028 61384 142034 61396
rect 161014 61384 161020 61396
rect 142028 61356 161020 61384
rect 142028 61344 142034 61356
rect 161014 61344 161020 61356
rect 161072 61344 161078 61396
rect 162762 61344 162768 61396
rect 162820 61384 162826 61396
rect 178402 61384 178408 61396
rect 162820 61356 178408 61384
rect 162820 61344 162826 61356
rect 178402 61344 178408 61356
rect 178460 61344 178466 61396
rect 180702 61344 180708 61396
rect 180760 61384 180766 61396
rect 193674 61384 193680 61396
rect 180760 61356 193680 61384
rect 180760 61344 180766 61356
rect 193674 61344 193680 61356
rect 193732 61344 193738 61396
rect 194410 61344 194416 61396
rect 194468 61384 194474 61396
rect 205910 61384 205916 61396
rect 194468 61356 205916 61384
rect 194468 61344 194474 61356
rect 205910 61344 205916 61356
rect 205968 61344 205974 61396
rect 210970 61344 210976 61396
rect 211028 61384 211034 61396
rect 220262 61384 220268 61396
rect 211028 61356 220268 61384
rect 211028 61344 211034 61356
rect 220262 61344 220268 61356
rect 220320 61344 220326 61396
rect 237190 61344 237196 61396
rect 237248 61384 237254 61396
rect 242894 61384 242900 61396
rect 237248 61356 242900 61384
rect 237248 61344 237254 61356
rect 242894 61344 242900 61356
rect 242952 61344 242958 61396
rect 408402 61344 408408 61396
rect 408460 61384 408466 61396
rect 429194 61384 429200 61396
rect 408460 61356 429200 61384
rect 408460 61344 408466 61356
rect 429194 61344 429200 61356
rect 429252 61344 429258 61396
rect 433150 61344 433156 61396
rect 433208 61384 433214 61396
rect 458358 61384 458364 61396
rect 433208 61356 458364 61384
rect 433208 61344 433214 61356
rect 458358 61344 458364 61356
rect 458416 61344 458422 61396
rect 463602 61344 463608 61396
rect 463660 61384 463666 61396
rect 494238 61384 494244 61396
rect 463660 61356 494244 61384
rect 463660 61344 463666 61356
rect 494238 61344 494244 61356
rect 494296 61344 494302 61396
rect 502242 61344 502248 61396
rect 502300 61384 502306 61396
rect 538306 61384 538312 61396
rect 502300 61356 538312 61384
rect 502300 61344 502306 61356
rect 538306 61344 538312 61356
rect 538364 61344 538370 61396
rect 539226 61344 539232 61396
rect 539284 61384 539290 61396
rect 548518 61384 548524 61396
rect 539284 61356 548524 61384
rect 539284 61344 539290 61356
rect 548518 61344 548524 61356
rect 548576 61344 548582 61396
rect 31662 61276 31668 61328
rect 31720 61316 31726 61328
rect 66254 61316 66260 61328
rect 31720 61288 66260 61316
rect 31720 61276 31726 61288
rect 66254 61276 66260 61288
rect 66312 61276 66318 61328
rect 67542 61276 67548 61328
rect 67600 61316 67606 61328
rect 96798 61316 96804 61328
rect 67600 61288 96804 61316
rect 67600 61276 67606 61288
rect 96798 61276 96804 61288
rect 96856 61276 96862 61328
rect 97902 61276 97908 61328
rect 97960 61316 97966 61328
rect 122282 61316 122288 61328
rect 97960 61288 122288 61316
rect 97960 61276 97966 61288
rect 122282 61276 122288 61288
rect 122340 61276 122346 61328
rect 125502 61276 125508 61328
rect 125560 61316 125566 61328
rect 145742 61316 145748 61328
rect 125560 61288 145748 61316
rect 125560 61276 125566 61288
rect 145742 61276 145748 61288
rect 145800 61276 145806 61328
rect 148962 61276 148968 61328
rect 149020 61316 149026 61328
rect 166166 61316 166172 61328
rect 149020 61288 166172 61316
rect 149020 61276 149026 61288
rect 166166 61276 166172 61288
rect 166224 61276 166230 61328
rect 168190 61276 168196 61328
rect 168248 61316 168254 61328
rect 182450 61316 182456 61328
rect 168248 61288 182456 61316
rect 168248 61276 168254 61288
rect 182450 61276 182456 61288
rect 182508 61276 182514 61328
rect 183462 61276 183468 61328
rect 183520 61316 183526 61328
rect 195974 61316 195980 61328
rect 183520 61288 195980 61316
rect 183520 61276 183526 61288
rect 195974 61276 195980 61288
rect 196032 61276 196038 61328
rect 206922 61276 206928 61328
rect 206980 61316 206986 61328
rect 216122 61316 216128 61328
rect 206980 61288 216128 61316
rect 206980 61276 206986 61288
rect 216122 61276 216128 61288
rect 216180 61276 216186 61328
rect 28902 61208 28908 61260
rect 28960 61248 28966 61260
rect 63494 61248 63500 61260
rect 28960 61220 63500 61248
rect 28960 61208 28966 61220
rect 63494 61208 63500 61220
rect 63552 61208 63558 61260
rect 64138 61208 64144 61260
rect 64196 61248 64202 61260
rect 70394 61248 70400 61260
rect 64196 61220 70400 61248
rect 64196 61208 64202 61220
rect 70394 61208 70400 61220
rect 70452 61208 70458 61260
rect 73062 61208 73068 61260
rect 73120 61248 73126 61260
rect 100846 61248 100852 61260
rect 73120 61220 100852 61248
rect 73120 61208 73126 61220
rect 100846 61208 100852 61220
rect 100904 61208 100910 61260
rect 104802 61208 104808 61260
rect 104860 61248 104866 61260
rect 128354 61248 128360 61260
rect 104860 61220 128360 61248
rect 104860 61208 104866 61220
rect 128354 61208 128360 61220
rect 128412 61208 128418 61260
rect 129642 61208 129648 61260
rect 129700 61248 129706 61260
rect 149790 61248 149796 61260
rect 129700 61220 149796 61248
rect 129700 61208 129706 61220
rect 149790 61208 149796 61220
rect 149848 61208 149854 61260
rect 150342 61208 150348 61260
rect 150400 61248 150406 61260
rect 167178 61248 167184 61260
rect 150400 61220 167184 61248
rect 150400 61208 150406 61220
rect 167178 61208 167184 61220
rect 167236 61208 167242 61260
rect 172422 61208 172428 61260
rect 172480 61248 172486 61260
rect 186590 61248 186596 61260
rect 172480 61220 186596 61248
rect 172480 61208 172486 61220
rect 186590 61208 186596 61220
rect 186648 61208 186654 61260
rect 194502 61208 194508 61260
rect 194560 61248 194566 61260
rect 204898 61248 204904 61260
rect 194560 61220 204904 61248
rect 194560 61208 194566 61220
rect 204898 61208 204904 61220
rect 204956 61208 204962 61260
rect 520918 61208 520924 61260
rect 520976 61248 520982 61260
rect 521562 61248 521568 61260
rect 520976 61220 521568 61248
rect 520976 61208 520982 61220
rect 521562 61208 521568 61220
rect 521620 61208 521626 61260
rect 33042 61140 33048 61192
rect 33100 61180 33106 61192
rect 59906 61180 59912 61192
rect 33100 61152 59912 61180
rect 33100 61140 33106 61152
rect 59906 61140 59912 61152
rect 59964 61140 59970 61192
rect 71590 61140 71596 61192
rect 71648 61180 71654 61192
rect 75362 61180 75368 61192
rect 71648 61152 75368 61180
rect 71648 61140 71654 61152
rect 75362 61140 75368 61152
rect 75420 61140 75426 61192
rect 75822 61140 75828 61192
rect 75880 61180 75886 61192
rect 103882 61180 103888 61192
rect 75880 61152 103888 61180
rect 75880 61140 75886 61152
rect 103882 61140 103888 61152
rect 103940 61140 103946 61192
rect 107562 61140 107568 61192
rect 107620 61180 107626 61192
rect 130470 61180 130476 61192
rect 107620 61152 130476 61180
rect 107620 61140 107626 61152
rect 130470 61140 130476 61152
rect 130528 61140 130534 61192
rect 139302 61140 139308 61192
rect 139360 61180 139366 61192
rect 157978 61180 157984 61192
rect 139360 61152 157984 61180
rect 139360 61140 139366 61152
rect 157978 61140 157984 61152
rect 158036 61140 158042 61192
rect 161382 61140 161388 61192
rect 161440 61180 161446 61192
rect 177390 61180 177396 61192
rect 161440 61152 177396 61180
rect 161440 61140 161446 61152
rect 177390 61140 177396 61152
rect 177448 61140 177454 61192
rect 179322 61140 179328 61192
rect 179380 61180 179386 61192
rect 192662 61180 192668 61192
rect 179380 61152 192668 61180
rect 179380 61140 179386 61152
rect 192662 61140 192668 61152
rect 192720 61140 192726 61192
rect 39942 61072 39948 61124
rect 40000 61112 40006 61124
rect 73338 61112 73344 61124
rect 40000 61084 73344 61112
rect 40000 61072 40006 61084
rect 73338 61072 73344 61084
rect 73396 61072 73402 61124
rect 75178 61072 75184 61124
rect 75236 61112 75242 61124
rect 76374 61112 76380 61124
rect 75236 61084 76380 61112
rect 75236 61072 75242 61084
rect 76374 61072 76380 61084
rect 76432 61072 76438 61124
rect 78582 61072 78588 61124
rect 78640 61112 78646 61124
rect 106274 61112 106280 61124
rect 78640 61084 106280 61112
rect 78640 61072 78646 61084
rect 106274 61072 106280 61084
rect 106332 61072 106338 61124
rect 114462 61072 114468 61124
rect 114520 61112 114526 61124
rect 136634 61112 136640 61124
rect 114520 61084 136640 61112
rect 114520 61072 114526 61084
rect 136634 61072 136640 61084
rect 136692 61072 136698 61124
rect 143442 61072 143448 61124
rect 143500 61112 143506 61124
rect 162118 61112 162124 61124
rect 143500 61084 162124 61112
rect 143500 61072 143506 61084
rect 162118 61072 162124 61084
rect 162176 61072 162182 61124
rect 166902 61072 166908 61124
rect 166960 61112 166966 61124
rect 181438 61112 181444 61124
rect 166960 61084 181444 61112
rect 166960 61072 166966 61084
rect 181438 61072 181444 61084
rect 181496 61072 181502 61124
rect 184750 61072 184756 61124
rect 184808 61112 184814 61124
rect 196802 61112 196808 61124
rect 184808 61084 196808 61112
rect 184808 61072 184814 61084
rect 196802 61072 196808 61084
rect 196860 61072 196866 61124
rect 233142 61072 233148 61124
rect 233200 61112 233206 61124
rect 238754 61112 238760 61124
rect 233200 61084 238760 61112
rect 233200 61072 233206 61084
rect 238754 61072 238760 61084
rect 238812 61072 238818 61124
rect 245470 61072 245476 61124
rect 245528 61112 245534 61124
rect 249794 61112 249800 61124
rect 245528 61084 249800 61112
rect 245528 61072 245534 61084
rect 249794 61072 249800 61084
rect 249852 61072 249858 61124
rect 256602 61072 256608 61124
rect 256660 61112 256666 61124
rect 258994 61112 259000 61124
rect 256660 61084 259000 61112
rect 256660 61072 256666 61084
rect 258994 61072 259000 61084
rect 259052 61072 259058 61124
rect 497458 61072 497464 61124
rect 497516 61112 497522 61124
rect 501598 61112 501604 61124
rect 497516 61084 501604 61112
rect 497516 61072 497522 61084
rect 501598 61072 501604 61084
rect 501656 61072 501662 61124
rect 38470 61004 38476 61056
rect 38528 61044 38534 61056
rect 72234 61044 72240 61056
rect 38528 61016 72240 61044
rect 38528 61004 38534 61016
rect 72234 61004 72240 61016
rect 72292 61004 72298 61056
rect 75270 61004 75276 61056
rect 75328 61044 75334 61056
rect 102870 61044 102876 61056
rect 75328 61016 102876 61044
rect 75328 61004 75334 61016
rect 102870 61004 102876 61016
rect 102928 61004 102934 61056
rect 103422 61004 103428 61056
rect 103480 61044 103486 61056
rect 127342 61044 127348 61056
rect 103480 61016 127348 61044
rect 103480 61004 103486 61016
rect 127342 61004 127348 61016
rect 127400 61004 127406 61056
rect 140682 61004 140688 61056
rect 140740 61044 140746 61056
rect 158990 61044 158996 61056
rect 140740 61016 158996 61044
rect 140740 61004 140746 61016
rect 158990 61004 158996 61016
rect 159048 61004 159054 61056
rect 223482 61004 223488 61056
rect 223540 61044 223546 61056
rect 230474 61044 230480 61056
rect 223540 61016 230480 61044
rect 223540 61004 223546 61016
rect 230474 61004 230480 61016
rect 230532 61004 230538 61056
rect 234522 61004 234528 61056
rect 234580 61044 234586 61056
rect 239674 61044 239680 61056
rect 234580 61016 239680 61044
rect 234580 61004 234586 61016
rect 239674 61004 239680 61016
rect 239732 61004 239738 61056
rect 241422 61004 241428 61056
rect 241480 61044 241486 61056
rect 245746 61044 245752 61056
rect 241480 61016 245752 61044
rect 241480 61004 241486 61016
rect 245746 61004 245752 61016
rect 245804 61004 245810 61056
rect 257982 61004 257988 61056
rect 258040 61044 258046 61056
rect 260006 61044 260012 61056
rect 258040 61016 260012 61044
rect 258040 61004 258046 61016
rect 260006 61004 260012 61016
rect 260064 61004 260070 61056
rect 535178 61004 535184 61056
rect 535236 61044 535242 61056
rect 540238 61044 540244 61056
rect 535236 61016 540244 61044
rect 535236 61004 535242 61016
rect 540238 61004 540244 61016
rect 540296 61004 540302 61056
rect 35802 60936 35808 60988
rect 35860 60976 35866 60988
rect 69198 60976 69204 60988
rect 35860 60948 69204 60976
rect 35860 60936 35866 60948
rect 69198 60936 69204 60948
rect 69256 60936 69262 60988
rect 71590 60976 71596 60988
rect 69676 60948 71596 60976
rect 42702 60868 42708 60920
rect 42760 60908 42766 60920
rect 69676 60908 69704 60948
rect 71590 60936 71596 60948
rect 71648 60936 71654 60988
rect 71682 60936 71688 60988
rect 71740 60976 71746 60988
rect 99834 60976 99840 60988
rect 71740 60948 99840 60976
rect 71740 60936 71746 60948
rect 99834 60936 99840 60948
rect 99892 60936 99898 60988
rect 117130 60936 117136 60988
rect 117188 60976 117194 60988
rect 138566 60976 138572 60988
rect 117188 60948 138572 60976
rect 117188 60936 117194 60948
rect 138566 60936 138572 60948
rect 138624 60936 138630 60988
rect 151722 60936 151728 60988
rect 151780 60976 151786 60988
rect 168374 60976 168380 60988
rect 151780 60948 168380 60976
rect 151780 60936 151786 60948
rect 168374 60936 168380 60948
rect 168432 60936 168438 60988
rect 235902 60936 235908 60988
rect 235960 60976 235966 60988
rect 240686 60976 240692 60988
rect 235960 60948 240692 60976
rect 235960 60936 235966 60948
rect 240686 60936 240692 60948
rect 240744 60936 240750 60988
rect 245562 60936 245568 60988
rect 245620 60976 245626 60988
rect 248782 60976 248788 60988
rect 245620 60948 248788 60976
rect 245620 60936 245626 60948
rect 248782 60936 248788 60948
rect 248840 60936 248846 60988
rect 251082 60936 251088 60988
rect 251140 60976 251146 60988
rect 253934 60976 253940 60988
rect 251140 60948 253940 60976
rect 251140 60936 251146 60948
rect 253934 60936 253940 60948
rect 253992 60936 253998 60988
rect 255222 60936 255228 60988
rect 255280 60976 255286 60988
rect 258166 60976 258172 60988
rect 255280 60948 258172 60976
rect 255280 60936 255286 60948
rect 258166 60936 258172 60948
rect 258224 60936 258230 60988
rect 42760 60880 69704 60908
rect 42760 60868 42766 60880
rect 74534 60868 74540 60920
rect 74592 60908 74598 60920
rect 78766 60908 78772 60920
rect 74592 60880 78772 60908
rect 74592 60868 74598 60880
rect 78766 60868 78772 60880
rect 78824 60868 78830 60920
rect 79962 60868 79968 60920
rect 80020 60908 80026 60920
rect 107010 60908 107016 60920
rect 80020 60880 107016 60908
rect 80020 60868 80026 60880
rect 107010 60868 107016 60880
rect 107068 60868 107074 60920
rect 115842 60868 115848 60920
rect 115900 60908 115906 60920
rect 137554 60908 137560 60920
rect 115900 60880 137560 60908
rect 115900 60868 115906 60880
rect 137554 60868 137560 60880
rect 137612 60868 137618 60920
rect 147582 60868 147588 60920
rect 147640 60908 147646 60920
rect 165154 60908 165160 60920
rect 147640 60880 165160 60908
rect 147640 60868 147646 60880
rect 165154 60868 165160 60880
rect 165212 60868 165218 60920
rect 242802 60868 242808 60920
rect 242860 60908 242866 60920
rect 247126 60908 247132 60920
rect 242860 60880 247132 60908
rect 242860 60868 242866 60880
rect 247126 60868 247132 60880
rect 247184 60868 247190 60920
rect 249702 60868 249708 60920
rect 249760 60908 249766 60920
rect 252922 60908 252928 60920
rect 249760 60880 252928 60908
rect 249760 60868 249766 60880
rect 252922 60868 252928 60880
rect 252980 60868 252986 60920
rect 253750 60868 253756 60920
rect 253808 60908 253814 60920
rect 256970 60908 256976 60920
rect 253808 60880 256976 60908
rect 253808 60868 253814 60880
rect 256970 60868 256976 60880
rect 257028 60868 257034 60920
rect 529014 60868 529020 60920
rect 529072 60908 529078 60920
rect 537478 60908 537484 60920
rect 529072 60880 537484 60908
rect 529072 60868 529078 60880
rect 537478 60868 537484 60880
rect 537536 60868 537542 60920
rect 40770 60800 40776 60852
rect 40828 60840 40834 60852
rect 55950 60840 55956 60852
rect 40828 60812 55956 60840
rect 40828 60800 40834 60812
rect 55950 60800 55956 60812
rect 56008 60800 56014 60852
rect 68278 60800 68284 60852
rect 68336 60840 68342 60852
rect 94682 60840 94688 60852
rect 68336 60812 94688 60840
rect 68336 60800 68342 60812
rect 94682 60800 94688 60812
rect 94740 60800 94746 60852
rect 119982 60800 119988 60852
rect 120040 60840 120046 60852
rect 141694 60840 141700 60852
rect 120040 60812 141700 60840
rect 120040 60800 120046 60812
rect 141694 60800 141700 60812
rect 141752 60800 141758 60852
rect 157242 60800 157248 60852
rect 157300 60840 157306 60852
rect 173342 60840 173348 60852
rect 157300 60812 173348 60840
rect 157300 60800 157306 60812
rect 173342 60800 173348 60812
rect 173400 60800 173406 60852
rect 231762 60800 231768 60852
rect 231820 60840 231826 60852
rect 237558 60840 237564 60852
rect 231820 60812 237564 60840
rect 231820 60800 231826 60812
rect 237558 60800 237564 60812
rect 237616 60800 237622 60852
rect 240042 60800 240048 60852
rect 240100 60840 240106 60852
rect 244734 60840 244740 60852
rect 240100 60812 244740 60840
rect 240100 60800 240106 60812
rect 244734 60800 244740 60812
rect 244792 60800 244798 60852
rect 252462 60800 252468 60852
rect 252520 60840 252526 60852
rect 255314 60840 255320 60852
rect 252520 60812 255320 60840
rect 252520 60800 252526 60812
rect 255314 60800 255320 60812
rect 255372 60800 255378 60852
rect 260742 60800 260748 60852
rect 260800 60840 260806 60852
rect 262214 60840 262220 60852
rect 260800 60812 262220 60840
rect 260800 60800 260806 60812
rect 262214 60800 262220 60812
rect 262272 60800 262278 60852
rect 264882 60800 264888 60852
rect 264940 60840 264946 60852
rect 266354 60840 266360 60852
rect 264940 60812 266360 60840
rect 264940 60800 264946 60812
rect 266354 60800 266360 60812
rect 266412 60800 266418 60852
rect 503530 60800 503536 60852
rect 503588 60840 503594 60852
rect 505738 60840 505744 60852
rect 503588 60812 505744 60840
rect 503588 60800 503594 60812
rect 505738 60800 505744 60812
rect 505796 60800 505802 60852
rect 512730 60800 512736 60852
rect 512788 60840 512794 60852
rect 515398 60840 515404 60852
rect 512788 60812 515404 60840
rect 512788 60800 512794 60812
rect 515398 60800 515404 60812
rect 515456 60800 515462 60852
rect 519906 60800 519912 60852
rect 519964 60840 519970 60852
rect 526438 60840 526444 60852
rect 519964 60812 526444 60840
rect 519964 60800 519970 60812
rect 526438 60800 526444 60812
rect 526496 60800 526502 60852
rect 531130 60800 531136 60852
rect 531188 60840 531194 60852
rect 533338 60840 533344 60852
rect 531188 60812 533344 60840
rect 531188 60800 531194 60812
rect 533338 60800 533344 60812
rect 533396 60800 533402 60852
rect 47578 60732 47584 60784
rect 47636 60772 47642 60784
rect 56962 60772 56968 60784
rect 47636 60744 56968 60772
rect 47636 60732 47642 60744
rect 56962 60732 56968 60744
rect 57020 60732 57026 60784
rect 59998 60732 60004 60784
rect 60056 60772 60062 60784
rect 64230 60772 64236 60784
rect 60056 60744 64236 60772
rect 60056 60732 60062 60744
rect 64230 60732 64236 60744
rect 64288 60732 64294 60784
rect 89622 60732 89628 60784
rect 89680 60772 89686 60784
rect 115106 60772 115112 60784
rect 89680 60744 115112 60772
rect 89680 60732 89686 60744
rect 115106 60732 115112 60744
rect 115164 60732 115170 60784
rect 121362 60732 121368 60784
rect 121420 60772 121426 60784
rect 142706 60772 142712 60784
rect 121420 60744 142712 60772
rect 121420 60732 121426 60744
rect 142706 60732 142712 60744
rect 142764 60732 142770 60784
rect 220722 60732 220728 60784
rect 220780 60772 220786 60784
rect 228358 60772 228364 60784
rect 220780 60744 228364 60772
rect 220780 60732 220786 60744
rect 228358 60732 228364 60744
rect 228416 60732 228422 60784
rect 230382 60732 230388 60784
rect 230440 60772 230446 60784
rect 236546 60772 236552 60784
rect 230440 60744 236552 60772
rect 230440 60732 230446 60744
rect 236546 60732 236552 60744
rect 236604 60732 236610 60784
rect 244182 60732 244188 60784
rect 244240 60772 244246 60784
rect 247770 60772 247776 60784
rect 244240 60744 247776 60772
rect 244240 60732 244246 60744
rect 247770 60732 247776 60744
rect 247828 60732 247834 60784
rect 249058 60732 249064 60784
rect 249116 60772 249122 60784
rect 251910 60772 251916 60784
rect 249116 60744 251916 60772
rect 249116 60732 249122 60744
rect 251910 60732 251916 60744
rect 251968 60732 251974 60784
rect 253842 60732 253848 60784
rect 253900 60772 253906 60784
rect 255958 60772 255964 60784
rect 253900 60744 255964 60772
rect 253900 60732 253906 60744
rect 255958 60732 255964 60744
rect 256016 60732 256022 60784
rect 259362 60732 259368 60784
rect 259420 60772 259426 60784
rect 261018 60772 261024 60784
rect 259420 60744 261024 60772
rect 259420 60732 259426 60744
rect 261018 60732 261024 60744
rect 261076 60732 261082 60784
rect 262122 60732 262128 60784
rect 262180 60772 262186 60784
rect 263134 60772 263140 60784
rect 262180 60744 263140 60772
rect 262180 60732 262186 60744
rect 263134 60732 263140 60744
rect 263192 60732 263198 60784
rect 263502 60732 263508 60784
rect 263560 60772 263566 60784
rect 265158 60772 265164 60784
rect 263560 60744 265164 60772
rect 263560 60732 263566 60744
rect 265158 60732 265164 60744
rect 265216 60732 265222 60784
rect 266262 60732 266268 60784
rect 266320 60772 266326 60784
rect 267182 60772 267188 60784
rect 266320 60744 267188 60772
rect 266320 60732 266326 60744
rect 267182 60732 267188 60744
rect 267240 60732 267246 60784
rect 286226 60732 286232 60784
rect 286284 60772 286290 60784
rect 286962 60772 286968 60784
rect 286284 60744 286968 60772
rect 286284 60732 286290 60744
rect 286962 60732 286968 60744
rect 287020 60732 287026 60784
rect 289262 60732 289268 60784
rect 289320 60772 289326 60784
rect 289998 60772 290004 60784
rect 289320 60744 290004 60772
rect 289320 60732 289326 60744
rect 289998 60732 290004 60744
rect 290056 60732 290062 60784
rect 290274 60732 290280 60784
rect 290332 60772 290338 60784
rect 291102 60772 291108 60784
rect 290332 60744 291108 60772
rect 290332 60732 290338 60744
rect 291102 60732 291108 60744
rect 291160 60732 291166 60784
rect 293310 60732 293316 60784
rect 293368 60772 293374 60784
rect 293862 60772 293868 60784
rect 293368 60744 293868 60772
rect 293368 60732 293374 60744
rect 293862 60732 293868 60744
rect 293920 60732 293926 60784
rect 294322 60732 294328 60784
rect 294380 60772 294386 60784
rect 295150 60772 295156 60784
rect 294380 60744 295156 60772
rect 294380 60732 294386 60744
rect 295150 60732 295156 60744
rect 295208 60732 295214 60784
rect 297450 60732 297456 60784
rect 297508 60772 297514 60784
rect 298002 60772 298008 60784
rect 297508 60744 298008 60772
rect 297508 60732 297514 60744
rect 298002 60732 298008 60744
rect 298060 60732 298066 60784
rect 298462 60732 298468 60784
rect 298520 60772 298526 60784
rect 299382 60772 299388 60784
rect 298520 60744 299388 60772
rect 298520 60732 298526 60744
rect 299382 60732 299388 60744
rect 299440 60732 299446 60784
rect 301498 60732 301504 60784
rect 301556 60772 301562 60784
rect 302142 60772 302148 60784
rect 301556 60744 302148 60772
rect 301556 60732 301562 60744
rect 302142 60732 302148 60744
rect 302200 60732 302206 60784
rect 302510 60732 302516 60784
rect 302568 60772 302574 60784
rect 303522 60772 303528 60784
rect 302568 60744 303528 60772
rect 302568 60732 302574 60744
rect 303522 60732 303528 60744
rect 303580 60732 303586 60784
rect 305546 60732 305552 60784
rect 305604 60772 305610 60784
rect 306282 60772 306288 60784
rect 305604 60744 306288 60772
rect 305604 60732 305610 60744
rect 306282 60732 306288 60744
rect 306340 60732 306346 60784
rect 309686 60732 309692 60784
rect 309744 60772 309750 60784
rect 310422 60772 310428 60784
rect 309744 60744 310428 60772
rect 309744 60732 309750 60744
rect 310422 60732 310428 60744
rect 310480 60732 310486 60784
rect 312722 60732 312728 60784
rect 312780 60772 312786 60784
rect 313182 60772 313188 60784
rect 312780 60744 313188 60772
rect 312780 60732 312786 60744
rect 313182 60732 313188 60744
rect 313240 60732 313246 60784
rect 313734 60732 313740 60784
rect 313792 60772 313798 60784
rect 314470 60772 314476 60784
rect 313792 60744 314476 60772
rect 313792 60732 313798 60744
rect 314470 60732 314476 60744
rect 314528 60732 314534 60784
rect 316770 60732 316776 60784
rect 316828 60772 316834 60784
rect 317322 60772 317328 60784
rect 316828 60744 317328 60772
rect 316828 60732 316834 60744
rect 317322 60732 317328 60744
rect 317380 60732 317386 60784
rect 317782 60732 317788 60784
rect 317840 60772 317846 60784
rect 318702 60772 318708 60784
rect 317840 60744 318708 60772
rect 317840 60732 317846 60744
rect 318702 60732 318708 60744
rect 318760 60732 318766 60784
rect 320910 60732 320916 60784
rect 320968 60772 320974 60784
rect 321462 60772 321468 60784
rect 320968 60744 321468 60772
rect 320968 60732 320974 60744
rect 321462 60732 321468 60744
rect 321520 60732 321526 60784
rect 321922 60732 321928 60784
rect 321980 60772 321986 60784
rect 322842 60772 322848 60784
rect 321980 60744 322848 60772
rect 321980 60732 321986 60744
rect 322842 60732 322848 60744
rect 322900 60732 322906 60784
rect 324958 60732 324964 60784
rect 325016 60772 325022 60784
rect 325602 60772 325608 60784
rect 325016 60744 325608 60772
rect 325016 60732 325022 60744
rect 325602 60732 325608 60744
rect 325660 60732 325666 60784
rect 325970 60732 325976 60784
rect 326028 60772 326034 60784
rect 326890 60772 326896 60784
rect 326028 60744 326896 60772
rect 326028 60732 326034 60744
rect 326890 60732 326896 60744
rect 326948 60732 326954 60784
rect 329006 60732 329012 60784
rect 329064 60772 329070 60784
rect 329742 60772 329748 60784
rect 329064 60744 329748 60772
rect 329064 60732 329070 60744
rect 329742 60732 329748 60744
rect 329800 60732 329806 60784
rect 330110 60732 330116 60784
rect 330168 60772 330174 60784
rect 331122 60772 331128 60784
rect 330168 60744 331128 60772
rect 330168 60732 330174 60744
rect 331122 60732 331128 60744
rect 331180 60732 331186 60784
rect 333146 60732 333152 60784
rect 333204 60772 333210 60784
rect 333882 60772 333888 60784
rect 333204 60744 333888 60772
rect 333204 60732 333210 60744
rect 333882 60732 333888 60744
rect 333940 60732 333946 60784
rect 336182 60732 336188 60784
rect 336240 60772 336246 60784
rect 336642 60772 336648 60784
rect 336240 60744 336648 60772
rect 336240 60732 336246 60744
rect 336642 60732 336648 60744
rect 336700 60732 336706 60784
rect 337194 60732 337200 60784
rect 337252 60772 337258 60784
rect 337930 60772 337936 60784
rect 337252 60744 337936 60772
rect 337252 60732 337258 60744
rect 337930 60732 337936 60744
rect 337988 60732 337994 60784
rect 340322 60732 340328 60784
rect 340380 60772 340386 60784
rect 340782 60772 340788 60784
rect 340380 60744 340788 60772
rect 340380 60732 340386 60744
rect 340782 60732 340788 60744
rect 340840 60732 340846 60784
rect 341334 60732 341340 60784
rect 341392 60772 341398 60784
rect 342070 60772 342076 60784
rect 341392 60744 342076 60772
rect 341392 60732 341398 60744
rect 342070 60732 342076 60744
rect 342128 60732 342134 60784
rect 344370 60732 344376 60784
rect 344428 60772 344434 60784
rect 344922 60772 344928 60784
rect 344428 60744 344928 60772
rect 344428 60732 344434 60744
rect 344922 60732 344928 60744
rect 344980 60732 344986 60784
rect 345382 60732 345388 60784
rect 345440 60772 345446 60784
rect 346302 60772 346308 60784
rect 345440 60744 346308 60772
rect 345440 60732 345446 60744
rect 346302 60732 346308 60744
rect 346360 60732 346366 60784
rect 348418 60732 348424 60784
rect 348476 60772 348482 60784
rect 349062 60772 349068 60784
rect 348476 60744 349068 60772
rect 348476 60732 348482 60744
rect 349062 60732 349068 60744
rect 349120 60732 349126 60784
rect 349430 60732 349436 60784
rect 349488 60772 349494 60784
rect 350350 60772 350356 60784
rect 349488 60744 350356 60772
rect 349488 60732 349494 60744
rect 350350 60732 350356 60744
rect 350408 60732 350414 60784
rect 352558 60732 352564 60784
rect 352616 60772 352622 60784
rect 353202 60772 353208 60784
rect 352616 60744 353208 60772
rect 352616 60732 352622 60744
rect 353202 60732 353208 60744
rect 353260 60732 353266 60784
rect 353570 60732 353576 60784
rect 353628 60772 353634 60784
rect 354582 60772 354588 60784
rect 353628 60744 354588 60772
rect 353628 60732 353634 60744
rect 354582 60732 354588 60744
rect 354640 60732 354646 60784
rect 356606 60732 356612 60784
rect 356664 60772 356670 60784
rect 357250 60772 357256 60784
rect 356664 60744 357256 60772
rect 356664 60732 356670 60744
rect 357250 60732 357256 60744
rect 357308 60732 357314 60784
rect 359642 60732 359648 60784
rect 359700 60772 359706 60784
rect 360102 60772 360108 60784
rect 359700 60744 360108 60772
rect 359700 60732 359706 60744
rect 360102 60732 360108 60744
rect 360160 60732 360166 60784
rect 360654 60732 360660 60784
rect 360712 60772 360718 60784
rect 361482 60772 361488 60784
rect 360712 60744 361488 60772
rect 360712 60732 360718 60744
rect 361482 60732 361488 60744
rect 361540 60732 361546 60784
rect 363782 60732 363788 60784
rect 363840 60772 363846 60784
rect 364242 60772 364248 60784
rect 363840 60744 364248 60772
rect 363840 60732 363846 60744
rect 364242 60732 364248 60744
rect 364300 60732 364306 60784
rect 364794 60732 364800 60784
rect 364852 60772 364858 60784
rect 365530 60772 365536 60784
rect 364852 60744 365536 60772
rect 364852 60732 364858 60744
rect 365530 60732 365536 60744
rect 365588 60732 365594 60784
rect 367830 60732 367836 60784
rect 367888 60772 367894 60784
rect 368382 60772 368388 60784
rect 367888 60744 368388 60772
rect 367888 60732 367894 60744
rect 368382 60732 368388 60744
rect 368440 60732 368446 60784
rect 368842 60732 368848 60784
rect 368900 60772 368906 60784
rect 369670 60772 369676 60784
rect 368900 60744 369676 60772
rect 368900 60732 368906 60744
rect 369670 60732 369676 60744
rect 369728 60732 369734 60784
rect 371878 60732 371884 60784
rect 371936 60772 371942 60784
rect 372522 60772 372528 60784
rect 371936 60744 372528 60772
rect 371936 60732 371942 60744
rect 372522 60732 372528 60744
rect 372580 60732 372586 60784
rect 372890 60732 372896 60784
rect 372948 60772 372954 60784
rect 373902 60772 373908 60784
rect 372948 60744 373908 60772
rect 372948 60732 372954 60744
rect 373902 60732 373908 60744
rect 373960 60732 373966 60784
rect 376018 60732 376024 60784
rect 376076 60772 376082 60784
rect 376662 60772 376668 60784
rect 376076 60744 376668 60772
rect 376076 60732 376082 60744
rect 376662 60732 376668 60744
rect 376720 60732 376726 60784
rect 377030 60732 377036 60784
rect 377088 60772 377094 60784
rect 377950 60772 377956 60784
rect 377088 60744 377956 60772
rect 377088 60732 377094 60744
rect 377950 60732 377956 60744
rect 378008 60732 378014 60784
rect 380066 60732 380072 60784
rect 380124 60772 380130 60784
rect 380802 60772 380808 60784
rect 380124 60744 380808 60772
rect 380124 60732 380130 60744
rect 380802 60732 380808 60744
rect 380860 60732 380866 60784
rect 383102 60732 383108 60784
rect 383160 60772 383166 60784
rect 383562 60772 383568 60784
rect 383160 60744 383568 60772
rect 383160 60732 383166 60744
rect 383562 60732 383568 60744
rect 383620 60732 383626 60784
rect 384114 60732 384120 60784
rect 384172 60772 384178 60784
rect 384850 60772 384856 60784
rect 384172 60744 384856 60772
rect 384172 60732 384178 60744
rect 384850 60732 384856 60744
rect 384908 60732 384914 60784
rect 387242 60732 387248 60784
rect 387300 60772 387306 60784
rect 387702 60772 387708 60784
rect 387300 60744 387708 60772
rect 387300 60732 387306 60744
rect 387702 60732 387708 60744
rect 387760 60732 387766 60784
rect 388254 60732 388260 60784
rect 388312 60772 388318 60784
rect 389082 60772 389088 60784
rect 388312 60744 389088 60772
rect 388312 60732 388318 60744
rect 389082 60732 389088 60744
rect 389140 60732 389146 60784
rect 391290 60732 391296 60784
rect 391348 60772 391354 60784
rect 391842 60772 391848 60784
rect 391348 60744 391848 60772
rect 391348 60732 391354 60744
rect 391842 60732 391848 60744
rect 391900 60732 391906 60784
rect 392302 60732 392308 60784
rect 392360 60772 392366 60784
rect 393222 60772 393228 60784
rect 392360 60744 393228 60772
rect 392360 60732 392366 60744
rect 393222 60732 393228 60744
rect 393280 60732 393286 60784
rect 395338 60732 395344 60784
rect 395396 60772 395402 60784
rect 395982 60772 395988 60784
rect 395396 60744 395988 60772
rect 395396 60732 395402 60744
rect 395982 60732 395988 60744
rect 396040 60732 396046 60784
rect 396442 60732 396448 60784
rect 396500 60772 396506 60784
rect 397270 60772 397276 60784
rect 396500 60744 397276 60772
rect 396500 60732 396506 60744
rect 397270 60732 397276 60744
rect 397328 60732 397334 60784
rect 400490 60732 400496 60784
rect 400548 60772 400554 60784
rect 401410 60772 401416 60784
rect 400548 60744 401416 60772
rect 400548 60732 400554 60744
rect 401410 60732 401416 60744
rect 401468 60732 401474 60784
rect 403526 60732 403532 60784
rect 403584 60772 403590 60784
rect 404262 60772 404268 60784
rect 403584 60744 404268 60772
rect 403584 60732 403590 60744
rect 404262 60732 404268 60744
rect 404320 60732 404326 60784
rect 406562 60732 406568 60784
rect 406620 60772 406626 60784
rect 407022 60772 407028 60784
rect 406620 60744 407028 60772
rect 406620 60732 406626 60744
rect 407022 60732 407028 60744
rect 407080 60732 407086 60784
rect 407666 60732 407672 60784
rect 407724 60772 407730 60784
rect 408402 60772 408408 60784
rect 407724 60744 408408 60772
rect 407724 60732 407730 60744
rect 408402 60732 408408 60744
rect 408460 60732 408466 60784
rect 410702 60732 410708 60784
rect 410760 60772 410766 60784
rect 411162 60772 411168 60784
rect 410760 60744 411168 60772
rect 410760 60732 410766 60744
rect 411162 60732 411168 60744
rect 411220 60732 411226 60784
rect 415762 60732 415768 60784
rect 415820 60772 415826 60784
rect 416682 60772 416688 60784
rect 415820 60744 416688 60772
rect 415820 60732 415826 60744
rect 416682 60732 416688 60744
rect 416740 60732 416746 60784
rect 418890 60732 418896 60784
rect 418948 60772 418954 60784
rect 419442 60772 419448 60784
rect 418948 60744 419448 60772
rect 418948 60732 418954 60744
rect 419442 60732 419448 60744
rect 419500 60732 419506 60784
rect 419902 60732 419908 60784
rect 419960 60772 419966 60784
rect 420822 60772 420828 60784
rect 419960 60744 420828 60772
rect 419960 60732 419966 60744
rect 420822 60732 420828 60744
rect 420880 60732 420886 60784
rect 422938 60732 422944 60784
rect 422996 60772 423002 60784
rect 423582 60772 423588 60784
rect 422996 60744 423588 60772
rect 422996 60732 423002 60744
rect 423582 60732 423588 60744
rect 423640 60732 423646 60784
rect 431126 60732 431132 60784
rect 431184 60772 431190 60784
rect 431862 60772 431868 60784
rect 431184 60744 431868 60772
rect 431184 60732 431190 60744
rect 431862 60732 431868 60744
rect 431920 60732 431926 60784
rect 434162 60732 434168 60784
rect 434220 60772 434226 60784
rect 434622 60772 434628 60784
rect 434220 60744 434628 60772
rect 434220 60732 434226 60744
rect 434622 60732 434628 60744
rect 434680 60732 434686 60784
rect 435174 60732 435180 60784
rect 435232 60772 435238 60784
rect 436002 60772 436008 60784
rect 435232 60744 436008 60772
rect 435232 60732 435238 60744
rect 436002 60732 436008 60744
rect 436060 60732 436066 60784
rect 438210 60732 438216 60784
rect 438268 60772 438274 60784
rect 438762 60772 438768 60784
rect 438268 60744 438768 60772
rect 438268 60732 438274 60744
rect 438762 60732 438768 60744
rect 438820 60732 438826 60784
rect 443362 60732 443368 60784
rect 443420 60772 443426 60784
rect 444282 60772 444288 60784
rect 443420 60744 444288 60772
rect 443420 60732 443426 60744
rect 444282 60732 444288 60744
rect 444340 60732 444346 60784
rect 446398 60732 446404 60784
rect 446456 60772 446462 60784
rect 447042 60772 447048 60784
rect 446456 60744 447048 60772
rect 446456 60732 446462 60744
rect 447042 60732 447048 60744
rect 447100 60732 447106 60784
rect 447410 60732 447416 60784
rect 447468 60772 447474 60784
rect 448422 60772 448428 60784
rect 447468 60744 448428 60772
rect 447468 60732 447474 60744
rect 448422 60732 448428 60744
rect 448480 60732 448486 60784
rect 450446 60732 450452 60784
rect 450504 60772 450510 60784
rect 451182 60772 451188 60784
rect 450504 60744 451188 60772
rect 450504 60732 450510 60744
rect 451182 60732 451188 60744
rect 451240 60732 451246 60784
rect 451550 60732 451556 60784
rect 451608 60772 451614 60784
rect 452470 60772 452476 60784
rect 451608 60744 452476 60772
rect 451608 60732 451614 60744
rect 452470 60732 452476 60744
rect 452528 60732 452534 60784
rect 458634 60732 458640 60784
rect 458692 60772 458698 60784
rect 459370 60772 459376 60784
rect 458692 60744 459376 60772
rect 458692 60732 458698 60744
rect 459370 60732 459376 60744
rect 459428 60732 459434 60784
rect 461670 60732 461676 60784
rect 461728 60772 461734 60784
rect 462222 60772 462228 60784
rect 461728 60744 462228 60772
rect 461728 60732 461734 60744
rect 462222 60732 462228 60744
rect 462280 60732 462286 60784
rect 462774 60732 462780 60784
rect 462832 60772 462838 60784
rect 463602 60772 463608 60784
rect 462832 60744 463608 60772
rect 462832 60732 462838 60744
rect 463602 60732 463608 60744
rect 463660 60732 463666 60784
rect 465810 60732 465816 60784
rect 465868 60772 465874 60784
rect 466362 60772 466368 60784
rect 465868 60744 466368 60772
rect 465868 60732 465874 60744
rect 466362 60732 466368 60744
rect 466420 60732 466426 60784
rect 469858 60732 469864 60784
rect 469916 60772 469922 60784
rect 470502 60772 470508 60784
rect 469916 60744 470508 60772
rect 469916 60732 469922 60744
rect 470502 60732 470508 60744
rect 470560 60732 470566 60784
rect 470870 60732 470876 60784
rect 470928 60772 470934 60784
rect 471882 60772 471888 60784
rect 470928 60744 471888 60772
rect 470928 60732 470934 60744
rect 471882 60732 471888 60744
rect 471940 60732 471946 60784
rect 473998 60732 474004 60784
rect 474056 60772 474062 60784
rect 474642 60772 474648 60784
rect 474056 60744 474648 60772
rect 474056 60732 474062 60744
rect 474642 60732 474648 60744
rect 474700 60732 474706 60784
rect 481082 60732 481088 60784
rect 481140 60772 481146 60784
rect 481542 60772 481548 60784
rect 481140 60744 481548 60772
rect 481140 60732 481146 60744
rect 481542 60732 481548 60744
rect 481600 60732 481606 60784
rect 482094 60732 482100 60784
rect 482152 60772 482158 60784
rect 482830 60772 482836 60784
rect 482152 60744 482836 60772
rect 482152 60732 482158 60744
rect 482830 60732 482836 60744
rect 482888 60732 482894 60784
rect 485222 60732 485228 60784
rect 485280 60772 485286 60784
rect 485682 60772 485688 60784
rect 485280 60744 485688 60772
rect 485280 60732 485286 60744
rect 485682 60732 485688 60744
rect 485740 60732 485746 60784
rect 486234 60732 486240 60784
rect 486292 60772 486298 60784
rect 487062 60772 487068 60784
rect 486292 60744 487068 60772
rect 486292 60732 486298 60744
rect 487062 60732 487068 60744
rect 487120 60732 487126 60784
rect 489270 60732 489276 60784
rect 489328 60772 489334 60784
rect 489822 60772 489828 60784
rect 489328 60744 489828 60772
rect 489328 60732 489334 60744
rect 489822 60732 489828 60744
rect 489880 60732 489886 60784
rect 493318 60732 493324 60784
rect 493376 60772 493382 60784
rect 493962 60772 493968 60784
rect 493376 60744 493968 60772
rect 493376 60732 493382 60744
rect 493962 60732 493968 60744
rect 494020 60732 494026 60784
rect 494330 60732 494336 60784
rect 494388 60772 494394 60784
rect 495250 60772 495256 60784
rect 494388 60744 495256 60772
rect 494388 60732 494394 60744
rect 495250 60732 495256 60744
rect 495308 60732 495314 60784
rect 498470 60732 498476 60784
rect 498528 60772 498534 60784
rect 499482 60772 499488 60784
rect 498528 60744 499488 60772
rect 498528 60732 498534 60744
rect 499482 60732 499488 60744
rect 499540 60732 499546 60784
rect 501506 60732 501512 60784
rect 501564 60772 501570 60784
rect 502242 60772 502248 60784
rect 501564 60744 502248 60772
rect 501564 60732 501570 60744
rect 502242 60732 502248 60744
rect 502300 60732 502306 60784
rect 504542 60732 504548 60784
rect 504600 60772 504606 60784
rect 505002 60772 505008 60784
rect 504600 60744 505008 60772
rect 504600 60732 504606 60744
rect 505002 60732 505008 60744
rect 505060 60732 505066 60784
rect 506382 60732 506388 60784
rect 506440 60772 506446 60784
rect 507118 60772 507124 60784
rect 506440 60744 507124 60772
rect 506440 60732 506446 60744
rect 507118 60732 507124 60744
rect 507176 60732 507182 60784
rect 509694 60732 509700 60784
rect 509752 60772 509758 60784
rect 511258 60772 511264 60784
rect 509752 60744 511264 60772
rect 509752 60732 509758 60744
rect 511258 60732 511264 60744
rect 511316 60732 511322 60784
rect 513742 60732 513748 60784
rect 513800 60772 513806 60784
rect 514662 60772 514668 60784
rect 513800 60744 514668 60772
rect 513800 60732 513806 60744
rect 514662 60732 514668 60744
rect 514720 60732 514726 60784
rect 528002 60732 528008 60784
rect 528060 60772 528066 60784
rect 528462 60772 528468 60784
rect 528060 60744 528468 60772
rect 528060 60732 528066 60744
rect 528462 60732 528468 60744
rect 528520 60732 528526 60784
rect 532142 60732 532148 60784
rect 532200 60772 532206 60784
rect 532602 60772 532608 60784
rect 532200 60744 532608 60772
rect 532200 60732 532206 60744
rect 532602 60732 532608 60744
rect 532660 60732 532666 60784
rect 533982 60732 533988 60784
rect 534040 60772 534046 60784
rect 536098 60772 536104 60784
rect 534040 60744 536104 60772
rect 534040 60732 534046 60744
rect 536098 60732 536104 60744
rect 536156 60732 536162 60784
rect 536190 60732 536196 60784
rect 536248 60772 536254 60784
rect 536742 60772 536748 60784
rect 536248 60744 536748 60772
rect 536248 60732 536254 60744
rect 536742 60732 536748 60744
rect 536800 60732 536806 60784
rect 42886 60664 42892 60716
rect 42944 60704 42950 60716
rect 43070 60704 43076 60716
rect 42944 60676 43076 60704
rect 42944 60664 42950 60676
rect 43070 60664 43076 60676
rect 43128 60664 43134 60716
rect 76558 60664 76564 60716
rect 76616 60704 76622 60716
rect 76742 60704 76748 60716
rect 76616 60676 76748 60704
rect 76616 60664 76622 60676
rect 76742 60664 76748 60676
rect 76800 60664 76806 60716
rect 520826 60664 520832 60716
rect 520884 60664 520890 60716
rect 520844 60636 520872 60664
rect 520918 60636 520924 60648
rect 520844 60608 520924 60636
rect 520918 60596 520924 60608
rect 520976 60596 520982 60648
rect 40126 59644 40132 59696
rect 40184 59684 40190 59696
rect 40678 59684 40684 59696
rect 40184 59656 40684 59684
rect 40184 59644 40190 59656
rect 40678 59644 40684 59656
rect 40736 59644 40742 59696
rect 42794 57876 42800 57928
rect 42852 57916 42858 57928
rect 43070 57916 43076 57928
rect 42852 57888 43076 57916
rect 42852 57876 42858 57888
rect 43070 57876 43076 57888
rect 43128 57876 43134 57928
rect 76466 57876 76472 57928
rect 76524 57916 76530 57928
rect 76742 57916 76748 57928
rect 76524 57888 76748 57916
rect 76524 57876 76530 57888
rect 76742 57876 76748 57888
rect 76800 57876 76806 57928
rect 74534 56652 74540 56704
rect 74592 56692 74598 56704
rect 75270 56692 75276 56704
rect 74592 56664 75276 56692
rect 74592 56652 74598 56664
rect 75270 56652 75276 56664
rect 75328 56652 75334 56704
rect 74626 56584 74632 56636
rect 74684 56624 74690 56636
rect 74810 56624 74816 56636
rect 74684 56596 74816 56624
rect 74684 56584 74690 56596
rect 74810 56584 74816 56596
rect 74868 56584 74874 56636
rect 74258 56516 74264 56568
rect 74316 56556 74322 56568
rect 74534 56556 74540 56568
rect 74316 56528 74540 56556
rect 74316 56516 74322 56528
rect 74534 56516 74540 56528
rect 74592 56516 74598 56568
rect 520734 53116 520740 53168
rect 520792 53156 520798 53168
rect 520918 53156 520924 53168
rect 520792 53128 520924 53156
rect 520792 53116 520798 53128
rect 520918 53116 520924 53128
rect 520976 53116 520982 53168
rect 113450 51144 113456 51196
rect 113508 51144 113514 51196
rect 516870 51144 516876 51196
rect 516928 51184 516934 51196
rect 516928 51156 517008 51184
rect 516928 51144 516934 51156
rect 113468 51060 113496 51144
rect 516980 51060 517008 51156
rect 113450 51008 113456 51060
rect 113508 51008 113514 51060
rect 516962 51008 516968 51060
rect 517020 51008 517026 51060
rect 42794 48288 42800 48340
rect 42852 48328 42858 48340
rect 42978 48328 42984 48340
rect 42852 48300 42984 48328
rect 42852 48288 42858 48300
rect 42978 48288 42984 48300
rect 43036 48288 43042 48340
rect 76466 48288 76472 48340
rect 76524 48328 76530 48340
rect 76650 48328 76656 48340
rect 76524 48300 76656 48328
rect 76524 48288 76530 48300
rect 76650 48288 76656 48300
rect 76708 48288 76714 48340
rect 113266 48288 113272 48340
rect 113324 48328 113330 48340
rect 113450 48328 113456 48340
rect 113324 48300 113456 48328
rect 113324 48288 113330 48300
rect 113450 48288 113456 48300
rect 113508 48288 113514 48340
rect 520734 48288 520740 48340
rect 520792 48328 520798 48340
rect 520918 48328 520924 48340
rect 520792 48300 520924 48328
rect 520792 48288 520798 48300
rect 520918 48288 520924 48300
rect 520976 48288 520982 48340
rect 516686 48220 516692 48272
rect 516744 48260 516750 48272
rect 516870 48260 516876 48272
rect 516744 48232 516876 48260
rect 516744 48220 516750 48232
rect 516870 48220 516876 48232
rect 516928 48220 516934 48272
rect 74258 46928 74264 46980
rect 74316 46968 74322 46980
rect 74442 46968 74448 46980
rect 74316 46940 74448 46968
rect 74316 46928 74322 46940
rect 74442 46928 74448 46940
rect 74500 46928 74506 46980
rect 76650 41556 76656 41608
rect 76708 41556 76714 41608
rect 76668 41472 76696 41556
rect 42978 41420 42984 41472
rect 43036 41420 43042 41472
rect 76650 41420 76656 41472
rect 76708 41420 76714 41472
rect 113266 41420 113272 41472
rect 113324 41420 113330 41472
rect 42996 41336 43024 41420
rect 113284 41392 113312 41420
rect 113358 41392 113364 41404
rect 113284 41364 113364 41392
rect 113358 41352 113364 41364
rect 113416 41352 113422 41404
rect 577498 41352 577504 41404
rect 577556 41392 577562 41404
rect 580534 41392 580540 41404
rect 577556 41364 580540 41392
rect 577556 41352 577562 41364
rect 580534 41352 580540 41364
rect 580592 41352 580598 41404
rect 42978 41284 42984 41336
rect 43036 41284 43042 41336
rect 76650 38808 76656 38820
rect 76576 38780 76656 38808
rect 76576 38684 76604 38780
rect 76650 38768 76656 38780
rect 76708 38768 76714 38820
rect 42886 38632 42892 38684
rect 42944 38672 42950 38684
rect 42978 38672 42984 38684
rect 42944 38644 42984 38672
rect 42944 38632 42950 38644
rect 42978 38632 42984 38644
rect 43036 38632 43042 38684
rect 76558 38632 76564 38684
rect 76616 38632 76622 38684
rect 113174 38564 113180 38616
rect 113232 38604 113238 38616
rect 113358 38604 113364 38616
rect 113232 38576 113364 38604
rect 113232 38564 113238 38576
rect 113358 38564 113364 38576
rect 113416 38564 113422 38616
rect 74350 37272 74356 37324
rect 74408 37312 74414 37324
rect 74442 37312 74448 37324
rect 74408 37284 74448 37312
rect 74408 37272 74414 37284
rect 74442 37272 74448 37284
rect 74500 37272 74506 37324
rect 74350 37136 74356 37188
rect 74408 37176 74414 37188
rect 74718 37176 74724 37188
rect 74408 37148 74724 37176
rect 74408 37136 74414 37148
rect 74718 37136 74724 37148
rect 74776 37136 74782 37188
rect 42886 33940 42892 33992
rect 42944 33980 42950 33992
rect 43254 33980 43260 33992
rect 42944 33952 43260 33980
rect 42944 33940 42950 33952
rect 43254 33940 43260 33952
rect 43312 33940 43318 33992
rect 521010 31764 521016 31816
rect 521068 31764 521074 31816
rect 516686 31696 516692 31748
rect 516744 31736 516750 31748
rect 516870 31736 516876 31748
rect 516744 31708 516876 31736
rect 516744 31696 516750 31708
rect 516870 31696 516876 31708
rect 516928 31696 516934 31748
rect 521028 31680 521056 31764
rect 521010 31628 521016 31680
rect 521068 31628 521074 31680
rect 39850 30268 39856 30320
rect 39908 30308 39914 30320
rect 579890 30308 579896 30320
rect 39908 30280 579896 30308
rect 39908 30268 39914 30280
rect 579890 30268 579896 30280
rect 579948 30268 579954 30320
rect 43070 28976 43076 29028
rect 43128 29016 43134 29028
rect 43254 29016 43260 29028
rect 43128 28988 43260 29016
rect 43128 28976 43134 28988
rect 43254 28976 43260 28988
rect 43312 28976 43318 29028
rect 113174 28976 113180 29028
rect 113232 29016 113238 29028
rect 113450 29016 113456 29028
rect 113232 28988 113456 29016
rect 113232 28976 113238 28988
rect 113450 28976 113456 28988
rect 113508 28976 113514 29028
rect 516594 28908 516600 28960
rect 516652 28948 516658 28960
rect 516870 28948 516876 28960
rect 516652 28920 516876 28948
rect 516652 28908 516658 28920
rect 516870 28908 516876 28920
rect 516928 28908 516934 28960
rect 520918 28908 520924 28960
rect 520976 28948 520982 28960
rect 521010 28948 521016 28960
rect 520976 28920 521016 28948
rect 520976 28908 520982 28920
rect 521010 28908 521016 28920
rect 521068 28908 521074 28960
rect 74258 27548 74264 27600
rect 74316 27588 74322 27600
rect 74442 27588 74448 27600
rect 74316 27560 74448 27588
rect 74316 27548 74322 27560
rect 74442 27548 74448 27560
rect 74500 27548 74506 27600
rect 3510 22040 3516 22092
rect 3568 22080 3574 22092
rect 538214 22080 538220 22092
rect 3568 22052 538220 22080
rect 3568 22040 3574 22052
rect 538214 22040 538220 22052
rect 538272 22040 538278 22092
rect 42886 19320 42892 19372
rect 42944 19360 42950 19372
rect 42978 19360 42984 19372
rect 42944 19332 42984 19360
rect 42944 19320 42950 19332
rect 42978 19320 42984 19332
rect 43036 19320 43042 19372
rect 516594 19320 516600 19372
rect 516652 19360 516658 19372
rect 516778 19360 516784 19372
rect 516652 19332 516784 19360
rect 516652 19320 516658 19332
rect 516778 19320 516784 19332
rect 516836 19320 516842 19372
rect 74074 17960 74080 18012
rect 74132 18000 74138 18012
rect 74258 18000 74264 18012
rect 74132 17972 74264 18000
rect 74132 17960 74138 17972
rect 74258 17960 74264 17972
rect 74316 17960 74322 18012
rect 74074 9664 74080 9716
rect 74132 9704 74138 9716
rect 74258 9704 74264 9716
rect 74132 9676 74264 9704
rect 74132 9664 74138 9676
rect 74258 9664 74264 9676
rect 74316 9664 74322 9716
rect 518710 6196 518716 6248
rect 518768 6236 518774 6248
rect 558362 6236 558368 6248
rect 518768 6208 558368 6236
rect 518768 6196 518774 6208
rect 558362 6196 558368 6208
rect 558420 6196 558426 6248
rect 528462 6128 528468 6180
rect 528520 6168 528526 6180
rect 569034 6168 569040 6180
rect 528520 6140 569040 6168
rect 528520 6128 528526 6140
rect 569034 6128 569040 6140
rect 569092 6128 569098 6180
rect 501598 5448 501604 5500
rect 501656 5488 501662 5500
rect 533430 5488 533436 5500
rect 501656 5460 533436 5488
rect 501656 5448 501662 5460
rect 533430 5448 533436 5460
rect 533488 5448 533494 5500
rect 531958 5380 531964 5432
rect 532016 5420 532022 5432
rect 565538 5420 565544 5432
rect 532016 5392 565544 5420
rect 532016 5380 532022 5392
rect 565538 5380 565544 5392
rect 565596 5380 565602 5432
rect 37366 5312 37372 5364
rect 37424 5352 37430 5364
rect 70670 5352 70676 5364
rect 37424 5324 70676 5352
rect 37424 5312 37430 5324
rect 70670 5312 70676 5324
rect 70728 5312 70734 5364
rect 482830 5312 482836 5364
rect 482888 5352 482894 5364
rect 515582 5352 515588 5364
rect 482888 5324 515588 5352
rect 482888 5312 482894 5324
rect 515582 5312 515588 5324
rect 515640 5312 515646 5364
rect 522298 5312 522304 5364
rect 522356 5352 522362 5364
rect 554774 5352 554780 5364
rect 522356 5324 554780 5352
rect 522356 5312 522362 5324
rect 554774 5312 554780 5324
rect 554832 5312 554838 5364
rect 33870 5244 33876 5296
rect 33928 5284 33934 5296
rect 67634 5284 67640 5296
rect 33928 5256 67640 5284
rect 33928 5244 33934 5256
rect 67634 5244 67640 5256
rect 67692 5244 67698 5296
rect 473262 5244 473268 5296
rect 473320 5284 473326 5296
rect 504818 5284 504824 5296
rect 473320 5256 504824 5284
rect 473320 5244 473326 5256
rect 504818 5244 504824 5256
rect 504876 5244 504882 5296
rect 505738 5244 505744 5296
rect 505796 5284 505802 5296
rect 540514 5284 540520 5296
rect 505796 5256 540520 5284
rect 505796 5244 505802 5256
rect 540514 5244 540520 5256
rect 540572 5244 540578 5296
rect 40954 5176 40960 5228
rect 41012 5216 41018 5228
rect 74626 5216 74632 5228
rect 41012 5188 74632 5216
rect 41012 5176 41018 5188
rect 74626 5176 74632 5188
rect 74684 5176 74690 5228
rect 478782 5176 478788 5228
rect 478840 5216 478846 5228
rect 511994 5216 512000 5228
rect 478840 5188 512000 5216
rect 478840 5176 478846 5188
rect 511994 5176 512000 5188
rect 512052 5176 512058 5228
rect 515398 5176 515404 5228
rect 515456 5216 515462 5228
rect 551186 5216 551192 5228
rect 515456 5188 551192 5216
rect 515456 5176 515462 5188
rect 551186 5176 551192 5188
rect 551244 5176 551250 5228
rect 30282 5108 30288 5160
rect 30340 5148 30346 5160
rect 64874 5148 64880 5160
rect 30340 5120 64880 5148
rect 30340 5108 30346 5120
rect 64874 5108 64880 5120
rect 64932 5108 64938 5160
rect 476022 5108 476028 5160
rect 476080 5148 476086 5160
rect 508406 5148 508412 5160
rect 476080 5120 508412 5148
rect 476080 5108 476086 5120
rect 508406 5108 508412 5120
rect 508464 5108 508470 5160
rect 511258 5108 511264 5160
rect 511316 5148 511322 5160
rect 547690 5148 547696 5160
rect 511316 5120 547696 5148
rect 511316 5108 511322 5120
rect 547690 5108 547696 5120
rect 547748 5108 547754 5160
rect 26694 5040 26700 5092
rect 26752 5080 26758 5092
rect 62114 5080 62120 5092
rect 26752 5052 62120 5080
rect 26752 5040 26758 5052
rect 62114 5040 62120 5052
rect 62172 5040 62178 5092
rect 500862 5040 500868 5092
rect 500920 5080 500926 5092
rect 536926 5080 536932 5092
rect 500920 5052 536932 5080
rect 500920 5040 500926 5052
rect 536926 5040 536932 5052
rect 536984 5040 536990 5092
rect 21910 4972 21916 5024
rect 21968 5012 21974 5024
rect 57974 5012 57980 5024
rect 21968 4984 57980 5012
rect 21968 4972 21974 4984
rect 57974 4972 57980 4984
rect 58032 4972 58038 5024
rect 470502 4972 470508 5024
rect 470560 5012 470566 5024
rect 501230 5012 501236 5024
rect 470560 4984 501236 5012
rect 470560 4972 470566 4984
rect 501230 4972 501236 4984
rect 501288 4972 501294 5024
rect 507118 4972 507124 5024
rect 507176 5012 507182 5024
rect 544102 5012 544108 5024
rect 507176 4984 544108 5012
rect 507176 4972 507182 4984
rect 544102 4972 544108 4984
rect 544160 4972 544166 5024
rect 12434 4904 12440 4956
rect 12492 4944 12498 4956
rect 49694 4944 49700 4956
rect 12492 4916 49700 4944
rect 12492 4904 12498 4916
rect 49694 4904 49700 4916
rect 49752 4904 49758 4956
rect 69474 4904 69480 4956
rect 69532 4944 69538 4956
rect 98270 4944 98276 4956
rect 69532 4916 98276 4944
rect 69532 4904 69538 4916
rect 98270 4904 98276 4916
rect 98328 4904 98334 4956
rect 485682 4904 485688 4956
rect 485740 4944 485746 4956
rect 519078 4944 519084 4956
rect 485740 4916 519084 4944
rect 485740 4904 485746 4916
rect 519078 4904 519084 4916
rect 519136 4904 519142 4956
rect 533338 4904 533344 4956
rect 533396 4944 533402 4956
rect 572622 4944 572628 4956
rect 533396 4916 572628 4944
rect 533396 4904 533402 4916
rect 572622 4904 572628 4916
rect 572680 4904 572686 4956
rect 17218 4836 17224 4888
rect 17276 4876 17282 4888
rect 53834 4876 53840 4888
rect 17276 4848 53840 4876
rect 17276 4836 17282 4848
rect 53834 4836 53840 4848
rect 53892 4836 53898 4888
rect 65978 4836 65984 4888
rect 66036 4876 66042 4888
rect 95234 4876 95240 4888
rect 66036 4848 95240 4876
rect 66036 4836 66042 4848
rect 95234 4836 95240 4848
rect 95292 4836 95298 4888
rect 488442 4836 488448 4888
rect 488500 4876 488506 4888
rect 522666 4876 522672 4888
rect 488500 4848 522672 4876
rect 488500 4836 488506 4848
rect 522666 4836 522672 4848
rect 522724 4836 522730 4888
rect 522850 4836 522856 4888
rect 522908 4876 522914 4888
rect 561950 4876 561956 4888
rect 522908 4848 561956 4876
rect 522908 4836 522914 4848
rect 561950 4836 561956 4848
rect 562008 4836 562014 4888
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 45554 4808 45560 4820
rect 7708 4780 45560 4808
rect 7708 4768 7714 4780
rect 45554 4768 45560 4780
rect 45612 4768 45618 4820
rect 47394 4768 47400 4820
rect 47452 4808 47458 4820
rect 77294 4808 77300 4820
rect 47452 4780 77300 4808
rect 47452 4768 47458 4780
rect 77294 4768 77300 4780
rect 77352 4768 77358 4820
rect 448330 4768 448336 4820
rect 448388 4808 448394 4820
rect 476298 4808 476304 4820
rect 448388 4780 476304 4808
rect 448388 4768 448394 4780
rect 476298 4768 476304 4780
rect 476356 4768 476362 4820
rect 495250 4768 495256 4820
rect 495308 4808 495314 4820
rect 529842 4808 529848 4820
rect 495308 4780 529848 4808
rect 495308 4768 495314 4780
rect 529842 4768 529848 4780
rect 529900 4768 529906 4820
rect 536098 4768 536104 4820
rect 536156 4808 536162 4820
rect 576210 4808 576216 4820
rect 536156 4780 576216 4808
rect 536156 4768 536162 4780
rect 576210 4768 576216 4780
rect 576268 4768 576274 4820
rect 42150 4088 42156 4140
rect 42208 4128 42214 4140
rect 42702 4128 42708 4140
rect 42208 4100 42708 4128
rect 42208 4088 42214 4100
rect 42702 4088 42708 4100
rect 42760 4088 42766 4140
rect 50522 4088 50528 4140
rect 50580 4128 50586 4140
rect 50982 4128 50988 4140
rect 50580 4100 50988 4128
rect 50580 4088 50586 4100
rect 50982 4088 50988 4100
rect 51040 4088 51046 4140
rect 71866 4088 71872 4140
rect 71924 4128 71930 4140
rect 73062 4128 73068 4140
rect 71924 4100 73068 4128
rect 71924 4088 71930 4100
rect 73062 4088 73068 4100
rect 73120 4088 73126 4140
rect 77846 4088 77852 4140
rect 77904 4128 77910 4140
rect 78582 4128 78588 4140
rect 77904 4100 78588 4128
rect 77904 4088 77910 4100
rect 78582 4088 78588 4100
rect 78640 4088 78646 4140
rect 79042 4088 79048 4140
rect 79100 4128 79106 4140
rect 79962 4128 79968 4140
rect 79100 4100 79968 4128
rect 79100 4088 79106 4100
rect 79962 4088 79968 4100
rect 80020 4088 80026 4140
rect 111150 4088 111156 4140
rect 111208 4128 111214 4140
rect 111702 4128 111708 4140
rect 111208 4100 111708 4128
rect 111208 4088 111214 4100
rect 111702 4088 111708 4100
rect 111760 4088 111766 4140
rect 112346 4088 112352 4140
rect 112404 4128 112410 4140
rect 113082 4128 113088 4140
rect 112404 4100 113088 4128
rect 112404 4088 112410 4100
rect 113082 4088 113088 4100
rect 113140 4088 113146 4140
rect 113542 4088 113548 4140
rect 113600 4128 113606 4140
rect 114462 4128 114468 4140
rect 113600 4100 114468 4128
rect 113600 4088 113606 4100
rect 114462 4088 114468 4100
rect 114520 4088 114526 4140
rect 115934 4088 115940 4140
rect 115992 4128 115998 4140
rect 117130 4128 117136 4140
rect 115992 4100 117136 4128
rect 115992 4088 115998 4100
rect 117130 4088 117136 4100
rect 117188 4088 117194 4140
rect 296622 4088 296628 4140
rect 296680 4128 296686 4140
rect 299106 4128 299112 4140
rect 296680 4100 299112 4128
rect 296680 4088 296686 4100
rect 299106 4088 299112 4100
rect 299164 4088 299170 4140
rect 304902 4088 304908 4140
rect 304960 4128 304966 4140
rect 308582 4128 308588 4140
rect 304960 4100 308588 4128
rect 304960 4088 304966 4100
rect 308582 4088 308588 4100
rect 308640 4088 308646 4140
rect 320082 4088 320088 4140
rect 320140 4128 320146 4140
rect 326430 4128 326436 4140
rect 320140 4100 326436 4128
rect 320140 4088 320146 4100
rect 326430 4088 326436 4100
rect 326488 4088 326494 4140
rect 339402 4088 339408 4140
rect 339460 4128 339466 4140
rect 348970 4128 348976 4140
rect 339460 4100 348976 4128
rect 339460 4088 339466 4100
rect 348970 4088 348976 4100
rect 349028 4088 349034 4140
rect 349062 4088 349068 4140
rect 349120 4128 349126 4140
rect 359734 4128 359740 4140
rect 349120 4100 359740 4128
rect 349120 4088 349126 4100
rect 359734 4088 359740 4100
rect 359792 4088 359798 4140
rect 362862 4088 362868 4140
rect 362920 4128 362926 4140
rect 376386 4128 376392 4140
rect 362920 4100 376392 4128
rect 362920 4088 362926 4100
rect 376386 4088 376392 4100
rect 376444 4088 376450 4140
rect 377950 4088 377956 4140
rect 378008 4128 378014 4140
rect 393038 4128 393044 4140
rect 378008 4100 393044 4128
rect 378008 4088 378014 4100
rect 393038 4088 393044 4100
rect 393096 4088 393102 4140
rect 395982 4088 395988 4140
rect 396040 4128 396046 4140
rect 414474 4128 414480 4140
rect 396040 4100 414480 4128
rect 396040 4088 396046 4100
rect 414474 4088 414480 4100
rect 414532 4088 414538 4140
rect 420822 4088 420828 4140
rect 420880 4128 420886 4140
rect 442994 4128 443000 4140
rect 420880 4100 443000 4128
rect 420880 4088 420886 4100
rect 442994 4088 443000 4100
rect 443052 4088 443058 4140
rect 449802 4088 449808 4140
rect 449860 4128 449866 4140
rect 477494 4128 477500 4140
rect 449860 4100 477500 4128
rect 449860 4088 449866 4100
rect 477494 4088 477500 4100
rect 477552 4088 477558 4140
rect 480162 4088 480168 4140
rect 480220 4128 480226 4140
rect 480220 4100 507532 4128
rect 480220 4088 480226 4100
rect 83826 4020 83832 4072
rect 83884 4060 83890 4072
rect 110506 4060 110512 4072
rect 83884 4032 110512 4060
rect 83884 4020 83890 4032
rect 110506 4020 110512 4032
rect 110564 4020 110570 4072
rect 295150 4020 295156 4072
rect 295208 4060 295214 4072
rect 296714 4060 296720 4072
rect 295208 4032 296720 4060
rect 295208 4020 295214 4032
rect 296714 4020 296720 4032
rect 296772 4020 296778 4072
rect 340782 4020 340788 4072
rect 340840 4060 340846 4072
rect 350258 4060 350264 4072
rect 340840 4032 350264 4060
rect 340840 4020 340846 4032
rect 350258 4020 350264 4032
rect 350316 4020 350322 4072
rect 351822 4020 351828 4072
rect 351880 4060 351886 4072
rect 363322 4060 363328 4072
rect 351880 4032 363328 4060
rect 351880 4020 351886 4032
rect 363322 4020 363328 4032
rect 363380 4020 363386 4072
rect 367002 4020 367008 4072
rect 367060 4060 367066 4072
rect 381170 4060 381176 4072
rect 367060 4032 381176 4060
rect 367060 4020 367066 4032
rect 381170 4020 381176 4032
rect 381228 4020 381234 4072
rect 382182 4020 382188 4072
rect 382240 4060 382246 4072
rect 399018 4060 399024 4072
rect 382240 4032 399024 4060
rect 382240 4020 382246 4032
rect 399018 4020 399024 4032
rect 399076 4020 399082 4072
rect 401410 4020 401416 4072
rect 401468 4060 401474 4072
rect 420362 4060 420368 4072
rect 401468 4032 420368 4060
rect 401468 4020 401474 4032
rect 420362 4020 420368 4032
rect 420420 4020 420426 4072
rect 423582 4020 423588 4072
rect 423640 4060 423646 4072
rect 446582 4060 446588 4072
rect 423640 4032 446588 4060
rect 423640 4020 423646 4032
rect 446582 4020 446588 4032
rect 446640 4020 446646 4072
rect 447042 4020 447048 4072
rect 447100 4060 447106 4072
rect 473906 4060 473912 4072
rect 447100 4032 473912 4060
rect 447100 4020 447106 4032
rect 473906 4020 473912 4032
rect 473964 4020 473970 4072
rect 474642 4020 474648 4072
rect 474700 4060 474706 4072
rect 506014 4060 506020 4072
rect 474700 4032 506020 4060
rect 474700 4020 474706 4032
rect 506014 4020 506020 4032
rect 506072 4020 506078 4072
rect 20714 3952 20720 4004
rect 20772 3992 20778 4004
rect 47578 3992 47584 4004
rect 20772 3964 47584 3992
rect 20772 3952 20778 3964
rect 47578 3952 47584 3964
rect 47636 3952 47642 4004
rect 64690 3952 64696 4004
rect 64748 3992 64754 4004
rect 68278 3992 68284 4004
rect 64748 3964 68284 3992
rect 64748 3952 64754 3964
rect 68278 3952 68284 3964
rect 68336 3952 68342 4004
rect 76650 3992 76656 4004
rect 73540 3964 76656 3992
rect 19518 3884 19524 3936
rect 19576 3924 19582 3936
rect 40678 3924 40684 3936
rect 19576 3896 40684 3924
rect 19576 3884 19582 3896
rect 40678 3884 40684 3896
rect 40736 3884 40742 3936
rect 46934 3884 46940 3936
rect 46992 3924 46998 3936
rect 73540 3924 73568 3964
rect 76650 3952 76656 3964
rect 76708 3952 76714 4004
rect 98086 3952 98092 4004
rect 98144 3992 98150 4004
rect 122834 3992 122840 4004
rect 98144 3964 122840 3992
rect 98144 3952 98150 3964
rect 122834 3952 122840 3964
rect 122892 3952 122898 4004
rect 332502 3952 332508 4004
rect 332560 3992 332566 4004
rect 340690 3992 340696 4004
rect 332560 3964 340696 3992
rect 332560 3952 332566 3964
rect 340690 3952 340696 3964
rect 340748 3952 340754 4004
rect 342070 3952 342076 4004
rect 342128 3992 342134 4004
rect 351362 3992 351368 4004
rect 342128 3964 351368 3992
rect 342128 3952 342134 3964
rect 351362 3952 351368 3964
rect 351420 3952 351426 4004
rect 354582 3952 354588 4004
rect 354640 3992 354646 4004
rect 365714 3992 365720 4004
rect 354640 3964 365720 3992
rect 354640 3952 354646 3964
rect 365714 3952 365720 3964
rect 365772 3952 365778 4004
rect 373902 3952 373908 4004
rect 373960 3992 373966 4004
rect 388254 3992 388260 4004
rect 373960 3964 388260 3992
rect 373960 3952 373966 3964
rect 388254 3952 388260 3964
rect 388312 3952 388318 4004
rect 390462 3952 390468 4004
rect 390520 3992 390526 4004
rect 408494 3992 408500 4004
rect 390520 3964 408500 3992
rect 390520 3952 390526 3964
rect 408494 3952 408500 3964
rect 408552 3952 408558 4004
rect 411162 3952 411168 4004
rect 411220 3992 411226 4004
rect 432322 3992 432328 4004
rect 411220 3964 432328 3992
rect 411220 3952 411226 3964
rect 432322 3952 432328 3964
rect 432380 3952 432386 4004
rect 438762 3952 438768 4004
rect 438820 3992 438826 4004
rect 464430 3992 464436 4004
rect 438820 3964 464436 3992
rect 438820 3952 438826 3964
rect 464430 3952 464436 3964
rect 464488 3952 464494 4004
rect 464982 3952 464988 4004
rect 465040 3992 465046 4004
rect 469490 3992 469496 4004
rect 465040 3964 469496 3992
rect 465040 3952 465046 3964
rect 469490 3952 469496 3964
rect 469548 3952 469554 4004
rect 471882 3952 471888 4004
rect 471940 3992 471946 4004
rect 502426 3992 502432 4004
rect 471940 3964 502432 3992
rect 471940 3952 471946 3964
rect 502426 3952 502432 3964
rect 502484 3952 502490 4004
rect 507302 3992 507308 4004
rect 504376 3964 507308 3992
rect 46992 3896 73568 3924
rect 46992 3884 46998 3896
rect 75178 3884 75184 3936
rect 75236 3924 75242 3936
rect 82998 3924 83004 3936
rect 75236 3896 83004 3924
rect 75236 3884 75242 3896
rect 82998 3884 83004 3896
rect 83056 3884 83062 3936
rect 84838 3884 84844 3936
rect 84896 3924 84902 3936
rect 86954 3924 86960 3936
rect 84896 3896 86960 3924
rect 84896 3884 84902 3896
rect 86954 3884 86960 3896
rect 87012 3884 87018 3936
rect 87322 3884 87328 3936
rect 87380 3924 87386 3936
rect 113358 3924 113364 3936
rect 87380 3896 113364 3924
rect 87380 3884 87386 3896
rect 113358 3884 113364 3896
rect 113416 3884 113422 3936
rect 325602 3884 325608 3936
rect 325660 3924 325666 3936
rect 332410 3924 332416 3936
rect 325660 3896 332416 3924
rect 325660 3884 325666 3896
rect 332410 3884 332416 3896
rect 332468 3884 332474 3936
rect 335262 3884 335268 3936
rect 335320 3924 335326 3936
rect 344278 3924 344284 3936
rect 335320 3896 344284 3924
rect 335320 3884 335326 3896
rect 344278 3884 344284 3896
rect 344336 3884 344342 3936
rect 347682 3884 347688 3936
rect 347740 3924 347746 3936
rect 358538 3924 358544 3936
rect 347740 3896 358544 3924
rect 347740 3884 347746 3896
rect 358538 3884 358544 3896
rect 358596 3884 358602 3936
rect 360102 3884 360108 3936
rect 360160 3924 360166 3936
rect 372798 3924 372804 3936
rect 360160 3896 372804 3924
rect 360160 3884 360166 3896
rect 372798 3884 372804 3896
rect 372856 3884 372862 3936
rect 378042 3884 378048 3936
rect 378100 3924 378106 3936
rect 394234 3924 394240 3936
rect 378100 3896 394240 3924
rect 378100 3884 378106 3896
rect 394234 3884 394240 3896
rect 394292 3884 394298 3936
rect 397270 3884 397276 3936
rect 397328 3924 397334 3936
rect 415670 3924 415676 3936
rect 397328 3896 415676 3924
rect 397328 3884 397334 3896
rect 415670 3884 415676 3896
rect 415728 3884 415734 3936
rect 419442 3884 419448 3936
rect 419500 3924 419506 3936
rect 441798 3924 441804 3936
rect 419500 3896 441804 3924
rect 419500 3884 419506 3896
rect 441798 3884 441804 3896
rect 441856 3884 441862 3936
rect 444190 3884 444196 3936
rect 444248 3924 444254 3936
rect 471514 3924 471520 3936
rect 444248 3896 471520 3924
rect 444248 3884 444254 3896
rect 471514 3884 471520 3896
rect 471572 3884 471578 3936
rect 477402 3884 477408 3936
rect 477460 3924 477466 3936
rect 504376 3924 504404 3964
rect 507302 3952 507308 3964
rect 507360 3952 507366 4004
rect 477460 3896 504404 3924
rect 507504 3924 507532 4100
rect 508498 4088 508504 4140
rect 508556 4128 508562 4140
rect 510798 4128 510804 4140
rect 508556 4100 510804 4128
rect 508556 4088 508562 4100
rect 510798 4088 510804 4100
rect 510856 4088 510862 4140
rect 514662 4088 514668 4140
rect 514720 4128 514726 4140
rect 552382 4128 552388 4140
rect 514720 4100 552388 4128
rect 514720 4088 514726 4100
rect 552382 4088 552388 4100
rect 552440 4088 552446 4140
rect 507762 4020 507768 4072
rect 507820 4060 507826 4072
rect 516870 4060 516876 4072
rect 507820 4032 516876 4060
rect 507820 4020 507826 4032
rect 516870 4020 516876 4032
rect 516928 4020 516934 4072
rect 516962 4020 516968 4072
rect 517020 4060 517026 4072
rect 521470 4060 521476 4072
rect 517020 4032 521476 4060
rect 517020 4020 517026 4032
rect 521470 4020 521476 4032
rect 521528 4020 521534 4072
rect 528462 4020 528468 4072
rect 528520 4060 528526 4072
rect 545298 4060 545304 4072
rect 528520 4032 545304 4060
rect 528520 4020 528526 4032
rect 545298 4020 545304 4032
rect 545356 4020 545362 4072
rect 547138 4020 547144 4072
rect 547196 4060 547202 4072
rect 575014 4060 575020 4072
rect 547196 4032 575020 4060
rect 547196 4020 547202 4032
rect 575014 4020 575020 4032
rect 575072 4020 575078 4072
rect 510522 3952 510528 4004
rect 510580 3992 510586 4004
rect 514846 3992 514852 4004
rect 510580 3964 514852 3992
rect 510580 3952 510586 3964
rect 514846 3952 514852 3964
rect 514904 3952 514910 4004
rect 528370 3952 528376 4004
rect 528428 3992 528434 4004
rect 542998 3992 543004 4004
rect 528428 3964 543004 3992
rect 528428 3952 528434 3964
rect 542998 3952 543004 3964
rect 543056 3952 543062 4004
rect 548518 3952 548524 4004
rect 548576 3992 548582 4004
rect 582190 3992 582196 4004
rect 548576 3964 582196 3992
rect 548576 3952 548582 3964
rect 582190 3952 582196 3964
rect 582248 3952 582254 4004
rect 513190 3924 513196 3936
rect 507504 3896 513196 3924
rect 477460 3884 477466 3896
rect 513190 3884 513196 3896
rect 513248 3884 513254 3936
rect 518802 3884 518808 3936
rect 518860 3924 518866 3936
rect 557166 3924 557172 3936
rect 518860 3896 557172 3924
rect 518860 3884 518866 3896
rect 557166 3884 557172 3896
rect 557224 3884 557230 3936
rect 36170 3816 36176 3868
rect 36228 3856 36234 3868
rect 64138 3856 64144 3868
rect 36228 3828 64144 3856
rect 36228 3816 36234 3828
rect 64138 3816 64144 3828
rect 64196 3816 64202 3868
rect 72970 3816 72976 3868
rect 73028 3856 73034 3868
rect 102134 3856 102140 3868
rect 73028 3828 102140 3856
rect 73028 3816 73034 3828
rect 102134 3816 102140 3828
rect 102192 3816 102198 3868
rect 313182 3816 313188 3868
rect 313240 3856 313246 3868
rect 318058 3856 318064 3868
rect 313240 3828 318064 3856
rect 313240 3816 313246 3828
rect 318058 3816 318064 3828
rect 318116 3816 318122 3868
rect 333882 3816 333888 3868
rect 333940 3856 333946 3868
rect 341886 3856 341892 3868
rect 333940 3828 341892 3856
rect 333940 3816 333946 3828
rect 341886 3816 341892 3828
rect 341944 3816 341950 3868
rect 342162 3816 342168 3868
rect 342220 3856 342226 3868
rect 352558 3856 352564 3868
rect 342220 3828 352564 3856
rect 342220 3816 342226 3828
rect 352558 3816 352564 3828
rect 352616 3816 352622 3868
rect 353202 3816 353208 3868
rect 353260 3856 353266 3868
rect 364518 3856 364524 3868
rect 353260 3828 364524 3856
rect 353260 3816 353266 3828
rect 364518 3816 364524 3828
rect 364576 3816 364582 3868
rect 365530 3816 365536 3868
rect 365588 3856 365594 3868
rect 378778 3856 378784 3868
rect 365588 3828 378784 3856
rect 365588 3816 365594 3828
rect 378778 3816 378784 3828
rect 378836 3816 378842 3868
rect 379422 3816 379428 3868
rect 379480 3856 379486 3868
rect 395430 3856 395436 3868
rect 379480 3828 395436 3856
rect 379480 3816 379486 3828
rect 395430 3816 395436 3828
rect 395488 3816 395494 3868
rect 397362 3816 397368 3868
rect 397420 3856 397426 3868
rect 416866 3856 416872 3868
rect 397420 3828 416872 3856
rect 397420 3816 397426 3828
rect 416866 3816 416872 3828
rect 416924 3816 416930 3868
rect 424962 3816 424968 3868
rect 425020 3856 425026 3868
rect 448974 3856 448980 3868
rect 425020 3828 448980 3856
rect 425020 3816 425026 3828
rect 448974 3816 448980 3828
rect 449032 3816 449038 3868
rect 459462 3816 459468 3868
rect 459520 3856 459526 3868
rect 489362 3856 489368 3868
rect 459520 3828 489368 3856
rect 459520 3816 459526 3828
rect 489362 3816 489368 3828
rect 489420 3816 489426 3868
rect 489822 3816 489828 3868
rect 489880 3856 489886 3868
rect 523862 3856 523868 3868
rect 489880 3828 523868 3856
rect 489880 3816 489886 3828
rect 523862 3816 523868 3828
rect 523920 3816 523926 3868
rect 524322 3816 524328 3868
rect 524380 3856 524386 3868
rect 564342 3856 564348 3868
rect 524380 3828 564348 3856
rect 524380 3816 524386 3828
rect 564342 3816 564348 3828
rect 564400 3816 564406 3868
rect 29086 3748 29092 3800
rect 29144 3788 29150 3800
rect 59998 3788 60004 3800
rect 29144 3760 60004 3788
rect 29144 3748 29150 3760
rect 59998 3748 60004 3760
rect 60056 3748 60062 3800
rect 62390 3748 62396 3800
rect 62448 3788 62454 3800
rect 92474 3788 92480 3800
rect 62448 3760 92480 3788
rect 62448 3748 62454 3760
rect 92474 3748 92480 3760
rect 92532 3748 92538 3800
rect 101582 3748 101588 3800
rect 101640 3788 101646 3800
rect 125778 3788 125784 3800
rect 101640 3760 125784 3788
rect 101640 3748 101646 3760
rect 125778 3748 125784 3760
rect 125836 3748 125842 3800
rect 328362 3748 328368 3800
rect 328420 3788 328426 3800
rect 335906 3788 335912 3800
rect 328420 3760 335912 3788
rect 328420 3748 328426 3760
rect 335906 3748 335912 3760
rect 335964 3748 335970 3800
rect 336642 3748 336648 3800
rect 336700 3788 336706 3800
rect 345474 3788 345480 3800
rect 336700 3760 345480 3788
rect 336700 3748 336706 3760
rect 345474 3748 345480 3760
rect 345532 3748 345538 3800
rect 346302 3748 346308 3800
rect 346360 3788 346366 3800
rect 356146 3788 356152 3800
rect 346360 3760 356152 3788
rect 346360 3748 346366 3760
rect 356146 3748 356152 3760
rect 356204 3748 356210 3800
rect 357250 3748 357256 3800
rect 357308 3788 357314 3800
rect 369210 3788 369216 3800
rect 357308 3760 369216 3788
rect 357308 3748 357314 3760
rect 369210 3748 369216 3760
rect 369268 3748 369274 3800
rect 371142 3748 371148 3800
rect 371200 3788 371206 3800
rect 385862 3788 385868 3800
rect 371200 3760 385868 3788
rect 371200 3748 371206 3760
rect 385862 3748 385868 3760
rect 385920 3748 385926 3800
rect 387702 3748 387708 3800
rect 387760 3788 387766 3800
rect 404906 3788 404912 3800
rect 387760 3760 404912 3788
rect 387760 3748 387766 3760
rect 404906 3748 404912 3760
rect 404964 3748 404970 3800
rect 408402 3748 408408 3800
rect 408460 3788 408466 3800
rect 428734 3788 428740 3800
rect 408460 3760 428740 3788
rect 408460 3748 408466 3760
rect 428734 3748 428740 3760
rect 428792 3748 428798 3800
rect 431862 3748 431868 3800
rect 431920 3788 431926 3800
rect 456058 3788 456064 3800
rect 431920 3760 456064 3788
rect 431920 3748 431926 3760
rect 456058 3748 456064 3760
rect 456116 3748 456122 3800
rect 456702 3748 456708 3800
rect 456760 3788 456766 3800
rect 485774 3788 485780 3800
rect 456760 3760 485780 3788
rect 456760 3748 456766 3760
rect 485774 3748 485780 3760
rect 485832 3748 485838 3800
rect 487062 3748 487068 3800
rect 487120 3788 487126 3800
rect 514478 3788 514484 3800
rect 487120 3760 514484 3788
rect 487120 3748 487126 3760
rect 514478 3748 514484 3760
rect 514536 3748 514542 3800
rect 521562 3748 521568 3800
rect 521620 3788 521626 3800
rect 560754 3788 560760 3800
rect 521620 3760 560760 3788
rect 521620 3748 521626 3760
rect 560754 3748 560760 3760
rect 560812 3748 560818 3800
rect 11238 3680 11244 3732
rect 11296 3720 11302 3732
rect 43438 3720 43444 3732
rect 11296 3692 43444 3720
rect 11296 3680 11302 3692
rect 43438 3680 43444 3692
rect 43496 3680 43502 3732
rect 44542 3680 44548 3732
rect 44600 3720 44606 3732
rect 47394 3720 47400 3732
rect 44600 3692 47400 3720
rect 44600 3680 44606 3692
rect 47394 3680 47400 3692
rect 47452 3680 47458 3732
rect 58802 3680 58808 3732
rect 58860 3720 58866 3732
rect 89806 3720 89812 3732
rect 58860 3692 89812 3720
rect 58860 3680 58866 3692
rect 89806 3680 89812 3692
rect 89864 3680 89870 3732
rect 90910 3680 90916 3732
rect 90968 3720 90974 3732
rect 90968 3692 91140 3720
rect 90968 3680 90974 3692
rect 5258 3612 5264 3664
rect 5316 3652 5322 3664
rect 42978 3652 42984 3664
rect 5316 3624 42984 3652
rect 5316 3612 5322 3624
rect 42978 3612 42984 3624
rect 43036 3612 43042 3664
rect 51626 3612 51632 3664
rect 51684 3652 51690 3664
rect 75178 3652 75184 3664
rect 51684 3624 75184 3652
rect 51684 3612 51690 3624
rect 75178 3612 75184 3624
rect 75236 3612 75242 3664
rect 81434 3612 81440 3664
rect 81492 3652 81498 3664
rect 82630 3652 82636 3664
rect 81492 3624 82636 3652
rect 81492 3612 81498 3624
rect 82630 3612 82636 3624
rect 82688 3612 82694 3664
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 41414 3584 41420 3596
rect 2924 3556 41420 3584
rect 2924 3544 2930 3556
rect 41414 3544 41420 3556
rect 41472 3544 41478 3596
rect 54018 3544 54024 3596
rect 54076 3584 54082 3596
rect 55122 3584 55128 3596
rect 54076 3556 55128 3584
rect 54076 3544 54082 3556
rect 55122 3544 55128 3556
rect 55180 3544 55186 3596
rect 59998 3544 60004 3596
rect 60056 3584 60062 3596
rect 60642 3584 60648 3596
rect 60056 3556 60648 3584
rect 60056 3544 60062 3556
rect 60642 3544 60648 3556
rect 60700 3544 60706 3596
rect 61194 3544 61200 3596
rect 61252 3584 61258 3596
rect 62022 3584 62028 3596
rect 61252 3556 62028 3584
rect 61252 3544 61258 3556
rect 62022 3544 62028 3556
rect 62080 3544 62086 3596
rect 62114 3544 62120 3596
rect 62172 3584 62178 3596
rect 84838 3584 84844 3596
rect 62172 3556 84844 3584
rect 62172 3544 62178 3556
rect 84838 3544 84844 3556
rect 84896 3544 84902 3596
rect 84930 3544 84936 3596
rect 84988 3584 84994 3596
rect 85482 3584 85488 3596
rect 84988 3556 85488 3584
rect 84988 3544 84994 3556
rect 85482 3544 85488 3556
rect 85540 3544 85546 3596
rect 86126 3544 86132 3596
rect 86184 3584 86190 3596
rect 86862 3584 86868 3596
rect 86184 3556 86868 3584
rect 86184 3544 86190 3556
rect 86862 3544 86868 3556
rect 86920 3544 86926 3596
rect 88518 3544 88524 3596
rect 88576 3584 88582 3596
rect 89622 3584 89628 3596
rect 88576 3556 89628 3584
rect 88576 3544 88582 3556
rect 89622 3544 89628 3556
rect 89680 3544 89686 3596
rect 89714 3544 89720 3596
rect 89772 3584 89778 3596
rect 91002 3584 91008 3596
rect 89772 3556 91008 3584
rect 89772 3544 89778 3556
rect 91002 3544 91008 3556
rect 91060 3544 91066 3596
rect 91112 3584 91140 3692
rect 94498 3680 94504 3732
rect 94556 3720 94562 3732
rect 120074 3720 120080 3732
rect 94556 3692 120080 3720
rect 94556 3680 94562 3692
rect 120074 3680 120080 3692
rect 120132 3680 120138 3732
rect 129734 3720 129740 3732
rect 122944 3692 129740 3720
rect 106366 3612 106372 3664
rect 106424 3652 106430 3664
rect 107562 3652 107568 3664
rect 106424 3624 107568 3652
rect 106424 3612 106430 3624
rect 107562 3612 107568 3624
rect 107620 3612 107626 3664
rect 117406 3584 117412 3596
rect 91112 3556 117412 3584
rect 117406 3544 117412 3556
rect 117464 3544 117470 3596
rect 119430 3544 119436 3596
rect 119488 3584 119494 3596
rect 119982 3584 119988 3596
rect 119488 3556 119988 3584
rect 119488 3544 119494 3556
rect 119982 3544 119988 3556
rect 120040 3544 120046 3596
rect 120626 3544 120632 3596
rect 120684 3584 120690 3596
rect 121362 3584 121368 3596
rect 120684 3556 121368 3584
rect 120684 3544 120690 3556
rect 121362 3544 121368 3556
rect 121420 3544 121426 3596
rect 121822 3544 121828 3596
rect 121880 3584 121886 3596
rect 122742 3584 122748 3596
rect 121880 3556 122748 3584
rect 121880 3544 121886 3556
rect 122742 3544 122748 3556
rect 122800 3544 122806 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 40126 3516 40132 3528
rect 1728 3488 40132 3516
rect 1728 3476 1734 3488
rect 40126 3476 40132 3488
rect 40184 3476 40190 3528
rect 45738 3476 45744 3528
rect 45796 3516 45802 3528
rect 46842 3516 46848 3528
rect 45796 3488 46848 3516
rect 45796 3476 45802 3488
rect 46842 3476 46848 3488
rect 46900 3476 46906 3528
rect 75086 3516 75092 3528
rect 46952 3488 75092 3516
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 40218 3448 40224 3460
rect 624 3420 40224 3448
rect 624 3408 630 3420
rect 40218 3408 40224 3420
rect 40276 3408 40282 3460
rect 43346 3408 43352 3460
rect 43404 3448 43410 3460
rect 46952 3448 46980 3488
rect 75086 3476 75092 3488
rect 75144 3476 75150 3528
rect 80072 3488 103928 3516
rect 43404 3420 46980 3448
rect 43404 3408 43410 3420
rect 52822 3408 52828 3460
rect 52880 3448 52886 3460
rect 53742 3448 53748 3460
rect 52880 3420 53748 3448
rect 52880 3408 52886 3420
rect 53742 3408 53748 3420
rect 53800 3408 53806 3460
rect 53852 3420 70624 3448
rect 8846 3340 8852 3392
rect 8904 3380 8910 3392
rect 9582 3380 9588 3392
rect 8904 3352 9588 3380
rect 8904 3340 8910 3352
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 10042 3340 10048 3392
rect 10100 3380 10106 3392
rect 10962 3380 10968 3392
rect 10100 3352 10968 3380
rect 10100 3340 10106 3352
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 16022 3340 16028 3392
rect 16080 3380 16086 3392
rect 16482 3380 16488 3392
rect 16080 3352 16488 3380
rect 16080 3340 16086 3352
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 24302 3340 24308 3392
rect 24360 3380 24366 3392
rect 24762 3380 24768 3392
rect 24360 3352 24768 3380
rect 24360 3340 24366 3352
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 25498 3340 25504 3392
rect 25556 3380 25562 3392
rect 26142 3380 26148 3392
rect 25556 3352 26148 3380
rect 25556 3340 25562 3352
rect 26142 3340 26148 3352
rect 26200 3340 26206 3392
rect 27890 3340 27896 3392
rect 27948 3380 27954 3392
rect 28902 3380 28908 3392
rect 27948 3352 28908 3380
rect 27948 3340 27954 3352
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 34974 3340 34980 3392
rect 35032 3380 35038 3392
rect 35802 3380 35808 3392
rect 35032 3352 35808 3380
rect 35032 3340 35038 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 48130 3340 48136 3392
rect 48188 3380 48194 3392
rect 53852 3380 53880 3420
rect 48188 3352 53880 3380
rect 48188 3340 48194 3352
rect 55214 3340 55220 3392
rect 55272 3380 55278 3392
rect 62114 3380 62120 3392
rect 55272 3352 62120 3380
rect 55272 3340 55278 3352
rect 62114 3340 62120 3352
rect 62172 3340 62178 3392
rect 63586 3340 63592 3392
rect 63644 3380 63650 3392
rect 64782 3380 64788 3392
rect 63644 3352 64788 3380
rect 63644 3340 63650 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 68278 3340 68284 3392
rect 68336 3380 68342 3392
rect 68922 3380 68928 3392
rect 68336 3352 68928 3380
rect 68336 3340 68342 3352
rect 68922 3340 68928 3352
rect 68980 3340 68986 3392
rect 70596 3312 70624 3420
rect 70670 3408 70676 3460
rect 70728 3448 70734 3460
rect 71682 3448 71688 3460
rect 70728 3420 71688 3448
rect 70728 3408 70734 3420
rect 71682 3408 71688 3420
rect 71740 3408 71746 3460
rect 76650 3408 76656 3460
rect 76708 3448 76714 3460
rect 80072 3448 80100 3488
rect 76708 3420 80100 3448
rect 76708 3408 76714 3420
rect 80238 3408 80244 3460
rect 80296 3448 80302 3460
rect 103900 3448 103928 3488
rect 103974 3476 103980 3528
rect 104032 3516 104038 3528
rect 104802 3516 104808 3528
rect 104032 3488 104808 3516
rect 104032 3476 104038 3488
rect 104802 3476 104808 3488
rect 104860 3476 104866 3528
rect 114738 3476 114744 3528
rect 114796 3516 114802 3528
rect 115842 3516 115848 3528
rect 114796 3488 115848 3516
rect 114796 3476 114802 3488
rect 115842 3476 115848 3488
rect 115900 3476 115906 3528
rect 122944 3516 122972 3692
rect 129734 3680 129740 3692
rect 129792 3680 129798 3732
rect 306282 3680 306288 3732
rect 306340 3720 306346 3732
rect 309778 3720 309784 3732
rect 306340 3692 309784 3720
rect 306340 3680 306346 3692
rect 309778 3680 309784 3692
rect 309836 3680 309842 3732
rect 337930 3680 337936 3732
rect 337988 3720 337994 3732
rect 346670 3720 346676 3732
rect 337988 3692 346676 3720
rect 337988 3680 337994 3692
rect 346670 3680 346676 3692
rect 346728 3680 346734 3732
rect 350350 3680 350356 3732
rect 350408 3720 350414 3732
rect 360930 3720 360936 3732
rect 350408 3692 360936 3720
rect 350408 3680 350414 3692
rect 360930 3680 360936 3692
rect 360988 3680 360994 3732
rect 361390 3680 361396 3732
rect 361448 3720 361454 3732
rect 375190 3720 375196 3732
rect 361448 3692 375196 3720
rect 361448 3680 361454 3692
rect 375190 3680 375196 3692
rect 375248 3680 375254 3732
rect 375282 3680 375288 3732
rect 375340 3720 375346 3732
rect 390646 3720 390652 3732
rect 375340 3692 390652 3720
rect 375340 3680 375346 3692
rect 390646 3680 390652 3692
rect 390704 3680 390710 3732
rect 394602 3680 394608 3732
rect 394660 3720 394666 3732
rect 413278 3720 413284 3732
rect 394660 3692 413284 3720
rect 394660 3680 394666 3692
rect 413278 3680 413284 3692
rect 413336 3680 413342 3732
rect 413922 3680 413928 3732
rect 413980 3720 413986 3732
rect 435818 3720 435824 3732
rect 413980 3692 435824 3720
rect 413980 3680 413986 3692
rect 435818 3680 435824 3692
rect 435876 3680 435882 3732
rect 441522 3680 441528 3732
rect 441580 3720 441586 3732
rect 467834 3720 467840 3732
rect 441580 3692 467840 3720
rect 441580 3680 441586 3692
rect 467834 3680 467840 3692
rect 467892 3680 467898 3732
rect 469122 3680 469128 3732
rect 469180 3720 469186 3732
rect 500126 3720 500132 3732
rect 469180 3692 500132 3720
rect 469180 3680 469186 3692
rect 500126 3680 500132 3692
rect 500184 3680 500190 3732
rect 505002 3680 505008 3732
rect 505060 3720 505066 3732
rect 541710 3720 541716 3732
rect 505060 3692 541716 3720
rect 505060 3680 505066 3692
rect 541710 3680 541716 3692
rect 541768 3680 541774 3732
rect 542998 3680 543004 3732
rect 543056 3720 543062 3732
rect 548886 3720 548892 3732
rect 543056 3692 548892 3720
rect 543056 3680 543062 3692
rect 548886 3680 548892 3692
rect 548944 3680 548950 3732
rect 552658 3680 552664 3732
rect 552716 3720 552722 3732
rect 580994 3720 581000 3732
rect 552716 3692 581000 3720
rect 552716 3680 552722 3692
rect 580994 3680 581000 3692
rect 581052 3680 581058 3732
rect 126606 3612 126612 3664
rect 126664 3652 126670 3664
rect 147674 3652 147680 3664
rect 126664 3624 147680 3652
rect 126664 3612 126670 3624
rect 147674 3612 147680 3624
rect 147732 3612 147738 3664
rect 314470 3612 314476 3664
rect 314528 3652 314534 3664
rect 319254 3652 319260 3664
rect 314528 3624 319260 3652
rect 314528 3612 314534 3624
rect 319254 3612 319260 3624
rect 319312 3612 319318 3664
rect 322842 3612 322848 3664
rect 322900 3652 322906 3664
rect 328822 3652 328828 3664
rect 322900 3624 328828 3652
rect 322900 3612 322906 3624
rect 328822 3612 328828 3624
rect 328880 3612 328886 3664
rect 331122 3612 331128 3664
rect 331180 3652 331186 3664
rect 338298 3652 338304 3664
rect 331180 3624 338304 3652
rect 331180 3612 331186 3624
rect 338298 3612 338304 3624
rect 338356 3612 338362 3664
rect 343542 3612 343548 3664
rect 343600 3652 343606 3664
rect 353754 3652 353760 3664
rect 343600 3624 353760 3652
rect 343600 3612 343606 3624
rect 353754 3612 353760 3624
rect 353812 3612 353818 3664
rect 354490 3612 354496 3664
rect 354548 3652 354554 3664
rect 366910 3652 366916 3664
rect 354548 3624 366916 3652
rect 354548 3612 354554 3624
rect 366910 3612 366916 3624
rect 366968 3612 366974 3664
rect 368382 3612 368388 3664
rect 368440 3652 368446 3664
rect 382366 3652 382372 3664
rect 368440 3624 382372 3652
rect 368440 3612 368446 3624
rect 382366 3612 382372 3624
rect 382424 3612 382430 3664
rect 383562 3612 383568 3664
rect 383620 3652 383626 3664
rect 400214 3652 400220 3664
rect 383620 3624 400220 3652
rect 383620 3612 383626 3624
rect 400214 3612 400220 3624
rect 400272 3612 400278 3664
rect 401502 3612 401508 3664
rect 401560 3652 401566 3664
rect 421558 3652 421564 3664
rect 401560 3624 421564 3652
rect 401560 3612 401566 3624
rect 421558 3612 421564 3624
rect 421616 3612 421622 3664
rect 429102 3612 429108 3664
rect 429160 3652 429166 3664
rect 453666 3652 453672 3664
rect 429160 3624 453672 3652
rect 429160 3612 429166 3624
rect 453666 3612 453672 3624
rect 453724 3612 453730 3664
rect 453942 3612 453948 3664
rect 454000 3652 454006 3664
rect 482278 3652 482284 3664
rect 454000 3624 482284 3652
rect 454000 3612 454006 3624
rect 482278 3612 482284 3624
rect 482336 3612 482342 3664
rect 482922 3612 482928 3664
rect 482980 3652 482986 3664
rect 516778 3652 516784 3664
rect 482980 3624 516784 3652
rect 482980 3612 482986 3624
rect 516778 3612 516784 3624
rect 516836 3612 516842 3664
rect 519446 3612 519452 3664
rect 519504 3652 519510 3664
rect 520366 3652 520372 3664
rect 519504 3624 520372 3652
rect 519504 3612 519510 3624
rect 520366 3612 520372 3624
rect 520424 3612 520430 3664
rect 522942 3612 522948 3664
rect 523000 3652 523006 3664
rect 563146 3652 563152 3664
rect 523000 3624 563152 3652
rect 523000 3612 523006 3624
rect 563146 3612 563152 3624
rect 563204 3612 563210 3664
rect 567838 3612 567844 3664
rect 567896 3652 567902 3664
rect 579798 3652 579804 3664
rect 567896 3624 579804 3652
rect 567896 3612 567902 3624
rect 579798 3612 579804 3624
rect 579856 3612 579862 3664
rect 127802 3544 127808 3596
rect 127860 3584 127866 3596
rect 149054 3584 149060 3596
rect 127860 3556 149060 3584
rect 127860 3544 127866 3556
rect 149054 3544 149060 3556
rect 149112 3544 149118 3596
rect 158714 3544 158720 3596
rect 158772 3584 158778 3596
rect 159910 3584 159916 3596
rect 158772 3556 159916 3584
rect 158772 3544 158778 3556
rect 159910 3544 159916 3556
rect 159968 3544 159974 3596
rect 167086 3544 167092 3596
rect 167144 3584 167150 3596
rect 168190 3584 168196 3596
rect 167144 3556 168196 3584
rect 167144 3544 167150 3556
rect 168190 3544 168196 3556
rect 168248 3544 168254 3596
rect 201494 3544 201500 3596
rect 201552 3584 201558 3596
rect 202690 3584 202696 3596
rect 201552 3556 202696 3584
rect 201552 3544 201558 3556
rect 202690 3544 202696 3556
rect 202748 3544 202754 3596
rect 227714 3544 227720 3596
rect 227772 3584 227778 3596
rect 228910 3584 228916 3596
rect 227772 3556 228916 3584
rect 227772 3544 227778 3556
rect 228910 3544 228916 3556
rect 228968 3544 228974 3596
rect 244366 3544 244372 3596
rect 244424 3584 244430 3596
rect 245562 3584 245568 3596
rect 244424 3556 245568 3584
rect 244424 3544 244430 3556
rect 245562 3544 245568 3556
rect 245620 3544 245626 3596
rect 252646 3544 252652 3596
rect 252704 3584 252710 3596
rect 253842 3584 253848 3596
rect 252704 3556 253848 3584
rect 252704 3544 252710 3556
rect 253842 3544 253848 3556
rect 253900 3544 253906 3596
rect 278866 3544 278872 3596
rect 278924 3584 278930 3596
rect 280062 3584 280068 3596
rect 278924 3556 280068 3584
rect 278924 3544 278930 3556
rect 280062 3544 280068 3556
rect 280120 3544 280126 3596
rect 293862 3544 293868 3596
rect 293920 3584 293926 3596
rect 295518 3584 295524 3596
rect 293920 3556 295524 3584
rect 293920 3544 293926 3556
rect 295518 3544 295524 3556
rect 295576 3544 295582 3596
rect 303430 3544 303436 3596
rect 303488 3584 303494 3596
rect 307386 3584 307392 3596
rect 303488 3556 307392 3584
rect 303488 3544 303494 3556
rect 307386 3544 307392 3556
rect 307444 3544 307450 3596
rect 314562 3544 314568 3596
rect 314620 3584 314626 3596
rect 320450 3584 320456 3596
rect 314620 3556 320456 3584
rect 314620 3544 314626 3556
rect 320450 3544 320456 3556
rect 320508 3544 320514 3596
rect 324222 3544 324228 3596
rect 324280 3584 324286 3596
rect 331214 3584 331220 3596
rect 324280 3556 331220 3584
rect 324280 3544 324286 3556
rect 331214 3544 331220 3556
rect 331272 3544 331278 3596
rect 333790 3544 333796 3596
rect 333848 3584 333854 3596
rect 343082 3584 343088 3596
rect 333848 3556 343088 3584
rect 333848 3544 333854 3556
rect 343082 3544 343088 3556
rect 343140 3544 343146 3596
rect 344922 3544 344928 3596
rect 344980 3584 344986 3596
rect 354950 3584 354956 3596
rect 344980 3556 354956 3584
rect 344980 3544 344986 3556
rect 354950 3544 354956 3556
rect 355008 3544 355014 3596
rect 357250 3544 357256 3596
rect 357308 3584 357314 3596
rect 370406 3584 370412 3596
rect 357308 3556 370412 3584
rect 357308 3544 357314 3556
rect 370406 3544 370412 3556
rect 370464 3544 370470 3596
rect 372522 3544 372528 3596
rect 372580 3584 372586 3596
rect 387058 3584 387064 3596
rect 372580 3556 387064 3584
rect 372580 3544 372586 3556
rect 387058 3544 387064 3556
rect 387116 3544 387122 3596
rect 388990 3544 388996 3596
rect 389048 3584 389054 3596
rect 407298 3584 407304 3596
rect 389048 3556 407304 3584
rect 389048 3544 389054 3556
rect 407298 3544 407304 3556
rect 407356 3544 407362 3596
rect 409782 3544 409788 3596
rect 409840 3584 409846 3596
rect 431126 3584 431132 3596
rect 409840 3556 431132 3584
rect 409840 3544 409846 3556
rect 431126 3544 431132 3556
rect 431184 3544 431190 3596
rect 431770 3544 431776 3596
rect 431828 3584 431834 3596
rect 457254 3584 457260 3596
rect 431828 3556 457260 3584
rect 431828 3544 431834 3556
rect 457254 3544 457260 3556
rect 457312 3544 457318 3596
rect 467742 3544 467748 3596
rect 467800 3584 467806 3596
rect 467800 3556 469260 3584
rect 467800 3544 467806 3556
rect 115952 3488 122972 3516
rect 104894 3448 104900 3460
rect 80296 3420 103836 3448
rect 103900 3420 104900 3448
rect 80296 3408 80302 3420
rect 93302 3340 93308 3392
rect 93360 3380 93366 3392
rect 93762 3380 93768 3392
rect 93360 3352 93768 3380
rect 93360 3340 93366 3352
rect 93762 3340 93768 3352
rect 93820 3340 93826 3392
rect 95694 3340 95700 3392
rect 95752 3380 95758 3392
rect 96522 3380 96528 3392
rect 95752 3352 96528 3380
rect 95752 3340 95758 3352
rect 96522 3340 96528 3352
rect 96580 3340 96586 3392
rect 96890 3340 96896 3392
rect 96948 3380 96954 3392
rect 97902 3380 97908 3392
rect 96948 3352 97908 3380
rect 96948 3340 96954 3352
rect 97902 3340 97908 3352
rect 97960 3340 97966 3392
rect 102778 3340 102784 3392
rect 102836 3380 102842 3392
rect 103422 3380 103428 3392
rect 102836 3352 103428 3380
rect 102836 3340 102842 3352
rect 103422 3340 103428 3352
rect 103480 3340 103486 3392
rect 103808 3380 103836 3420
rect 104894 3408 104900 3420
rect 104952 3408 104958 3460
rect 107654 3448 107660 3460
rect 105004 3420 107660 3448
rect 105004 3380 105032 3420
rect 107654 3408 107660 3420
rect 107712 3408 107718 3460
rect 103808 3352 105032 3380
rect 105170 3340 105176 3392
rect 105228 3380 105234 3392
rect 115952 3380 115980 3488
rect 123018 3476 123024 3528
rect 123076 3516 123082 3528
rect 124122 3516 124128 3528
rect 123076 3488 124128 3516
rect 123076 3476 123082 3488
rect 124122 3476 124128 3488
rect 124180 3476 124186 3528
rect 128998 3476 129004 3528
rect 129056 3516 129062 3528
rect 129642 3516 129648 3528
rect 129056 3488 129648 3516
rect 129056 3476 129062 3488
rect 129642 3476 129648 3488
rect 129700 3476 129706 3528
rect 130194 3476 130200 3528
rect 130252 3516 130258 3528
rect 130252 3488 145604 3516
rect 130252 3476 130258 3488
rect 105228 3352 115980 3380
rect 116044 3420 132540 3448
rect 105228 3340 105234 3352
rect 80054 3312 80060 3324
rect 70596 3284 80060 3312
rect 80054 3272 80060 3284
rect 80112 3272 80118 3324
rect 108758 3272 108764 3324
rect 108816 3312 108822 3324
rect 116044 3312 116072 3420
rect 131390 3340 131396 3392
rect 131448 3380 131454 3392
rect 132402 3380 132408 3392
rect 131448 3352 132408 3380
rect 131448 3340 131454 3352
rect 132402 3340 132408 3352
rect 132460 3340 132466 3392
rect 108816 3284 116072 3312
rect 108816 3272 108822 3284
rect 124214 3272 124220 3324
rect 124272 3312 124278 3324
rect 125502 3312 125508 3324
rect 124272 3284 125508 3312
rect 124272 3272 124278 3284
rect 125502 3272 125508 3284
rect 125560 3272 125566 3324
rect 132512 3312 132540 3420
rect 132586 3408 132592 3460
rect 132644 3448 132650 3460
rect 133690 3448 133696 3460
rect 132644 3420 133696 3448
rect 132644 3408 132650 3420
rect 133690 3408 133696 3420
rect 133748 3408 133754 3460
rect 136082 3408 136088 3460
rect 136140 3448 136146 3460
rect 136542 3448 136548 3460
rect 136140 3420 136548 3448
rect 136140 3408 136146 3420
rect 136542 3408 136548 3420
rect 136600 3408 136606 3460
rect 137278 3408 137284 3460
rect 137336 3448 137342 3460
rect 137922 3448 137928 3460
rect 137336 3420 137928 3448
rect 137336 3408 137342 3420
rect 137922 3408 137928 3420
rect 137980 3408 137986 3460
rect 138474 3408 138480 3460
rect 138532 3448 138538 3460
rect 139302 3448 139308 3460
rect 138532 3420 139308 3448
rect 138532 3408 138538 3420
rect 139302 3408 139308 3420
rect 139360 3408 139366 3460
rect 139670 3408 139676 3460
rect 139728 3448 139734 3460
rect 140682 3448 140688 3460
rect 139728 3420 140688 3448
rect 139728 3408 139734 3420
rect 140682 3408 140688 3420
rect 140740 3408 140746 3460
rect 145576 3380 145604 3488
rect 145650 3476 145656 3528
rect 145708 3516 145714 3528
rect 146202 3516 146208 3528
rect 145708 3488 146208 3516
rect 145708 3476 145714 3488
rect 146202 3476 146208 3488
rect 146260 3476 146266 3528
rect 146846 3476 146852 3528
rect 146904 3516 146910 3528
rect 147582 3516 147588 3528
rect 146904 3488 147588 3516
rect 146904 3476 146910 3488
rect 147582 3476 147588 3488
rect 147640 3476 147646 3528
rect 148042 3476 148048 3528
rect 148100 3516 148106 3528
rect 148962 3516 148968 3528
rect 148100 3488 148968 3516
rect 148100 3476 148106 3488
rect 148962 3476 148968 3488
rect 149020 3476 149026 3528
rect 150434 3476 150440 3528
rect 150492 3516 150498 3528
rect 151722 3516 151728 3528
rect 150492 3488 151728 3516
rect 150492 3476 150498 3488
rect 151722 3476 151728 3488
rect 151780 3476 151786 3528
rect 153930 3476 153936 3528
rect 153988 3516 153994 3528
rect 154482 3516 154488 3528
rect 153988 3488 154488 3516
rect 153988 3476 153994 3488
rect 154482 3476 154488 3488
rect 154540 3476 154546 3528
rect 155126 3476 155132 3528
rect 155184 3516 155190 3528
rect 155862 3516 155868 3528
rect 155184 3488 155868 3516
rect 155184 3476 155190 3488
rect 155862 3476 155868 3488
rect 155920 3476 155926 3528
rect 156322 3476 156328 3528
rect 156380 3516 156386 3528
rect 157242 3516 157248 3528
rect 156380 3488 157248 3516
rect 156380 3476 156386 3488
rect 157242 3476 157248 3488
rect 157300 3476 157306 3528
rect 162302 3476 162308 3528
rect 162360 3516 162366 3528
rect 162762 3516 162768 3528
rect 162360 3488 162768 3516
rect 162360 3476 162366 3488
rect 162762 3476 162768 3488
rect 162820 3476 162826 3528
rect 163498 3476 163504 3528
rect 163556 3516 163562 3528
rect 164142 3516 164148 3528
rect 163556 3488 164148 3516
rect 163556 3476 163562 3488
rect 164142 3476 164148 3488
rect 164200 3476 164206 3528
rect 165890 3476 165896 3528
rect 165948 3516 165954 3528
rect 166902 3516 166908 3528
rect 165948 3488 166908 3516
rect 165948 3476 165954 3488
rect 166902 3476 166908 3488
rect 166960 3476 166966 3528
rect 171778 3476 171784 3528
rect 171836 3516 171842 3528
rect 172422 3516 172428 3528
rect 171836 3488 172428 3516
rect 171836 3476 171842 3488
rect 172422 3476 172428 3488
rect 172480 3476 172486 3528
rect 172974 3476 172980 3528
rect 173032 3516 173038 3528
rect 173802 3516 173808 3528
rect 173032 3488 173808 3516
rect 173032 3476 173038 3488
rect 173802 3476 173808 3488
rect 173860 3476 173866 3528
rect 180150 3476 180156 3528
rect 180208 3516 180214 3528
rect 180702 3516 180708 3528
rect 180208 3488 180708 3516
rect 180208 3476 180214 3488
rect 180702 3476 180708 3488
rect 180760 3476 180766 3528
rect 182542 3476 182548 3528
rect 182600 3516 182606 3528
rect 183462 3516 183468 3528
rect 182600 3488 183468 3516
rect 182600 3476 182606 3488
rect 183462 3476 183468 3488
rect 183520 3476 183526 3528
rect 183738 3476 183744 3528
rect 183796 3516 183802 3528
rect 184750 3516 184756 3528
rect 183796 3488 184756 3516
rect 183796 3476 183802 3488
rect 184750 3476 184756 3488
rect 184808 3476 184814 3528
rect 188430 3476 188436 3528
rect 188488 3516 188494 3528
rect 188982 3516 188988 3528
rect 188488 3488 188988 3516
rect 188488 3476 188494 3488
rect 188982 3476 188988 3488
rect 189040 3476 189046 3528
rect 189626 3476 189632 3528
rect 189684 3516 189690 3528
rect 190362 3516 190368 3528
rect 189684 3488 190368 3516
rect 189684 3476 189690 3488
rect 190362 3476 190368 3488
rect 190420 3476 190426 3528
rect 192018 3476 192024 3528
rect 192076 3516 192082 3528
rect 193122 3516 193128 3528
rect 192076 3488 193128 3516
rect 192076 3476 192082 3488
rect 193122 3476 193128 3488
rect 193180 3476 193186 3528
rect 193214 3476 193220 3528
rect 193272 3516 193278 3528
rect 194502 3516 194508 3528
rect 193272 3488 194508 3516
rect 193272 3476 193278 3488
rect 194502 3476 194508 3488
rect 194560 3476 194566 3528
rect 196802 3476 196808 3528
rect 196860 3516 196866 3528
rect 197262 3516 197268 3528
rect 196860 3488 197268 3516
rect 196860 3476 196866 3488
rect 197262 3476 197268 3488
rect 197320 3476 197326 3528
rect 197998 3476 198004 3528
rect 198056 3516 198062 3528
rect 198642 3516 198648 3528
rect 198056 3488 198648 3516
rect 198056 3476 198062 3488
rect 198642 3476 198648 3488
rect 198700 3476 198706 3528
rect 199194 3476 199200 3528
rect 199252 3516 199258 3528
rect 200022 3516 200028 3528
rect 199252 3488 200028 3516
rect 199252 3476 199258 3488
rect 200022 3476 200028 3488
rect 200080 3476 200086 3528
rect 200390 3476 200396 3528
rect 200448 3516 200454 3528
rect 201402 3516 201408 3528
rect 200448 3488 201408 3516
rect 200448 3476 200454 3488
rect 201402 3476 201408 3488
rect 201460 3476 201466 3528
rect 205082 3476 205088 3528
rect 205140 3516 205146 3528
rect 205542 3516 205548 3528
rect 205140 3488 205548 3516
rect 205140 3476 205146 3488
rect 205542 3476 205548 3488
rect 205600 3476 205606 3528
rect 207474 3476 207480 3528
rect 207532 3516 207538 3528
rect 208302 3516 208308 3528
rect 207532 3488 208308 3516
rect 207532 3476 207538 3488
rect 208302 3476 208308 3488
rect 208360 3476 208366 3528
rect 208670 3476 208676 3528
rect 208728 3516 208734 3528
rect 209682 3516 209688 3528
rect 208728 3488 209688 3516
rect 208728 3476 208734 3488
rect 209682 3476 209688 3488
rect 209740 3476 209746 3528
rect 209866 3476 209872 3528
rect 209924 3516 209930 3528
rect 211062 3516 211068 3528
rect 209924 3488 211068 3516
rect 209924 3476 209930 3488
rect 211062 3476 211068 3488
rect 211120 3476 211126 3528
rect 214650 3476 214656 3528
rect 214708 3516 214714 3528
rect 215202 3516 215208 3528
rect 214708 3488 215208 3516
rect 214708 3476 214714 3488
rect 215202 3476 215208 3488
rect 215260 3476 215266 3528
rect 215846 3476 215852 3528
rect 215904 3516 215910 3528
rect 216582 3516 216588 3528
rect 215904 3488 216588 3516
rect 215904 3476 215910 3488
rect 216582 3476 216588 3488
rect 216640 3476 216646 3528
rect 217042 3476 217048 3528
rect 217100 3516 217106 3528
rect 217962 3516 217968 3528
rect 217100 3488 217968 3516
rect 217100 3476 217106 3488
rect 217962 3476 217968 3488
rect 218020 3476 218026 3528
rect 218146 3476 218152 3528
rect 218204 3516 218210 3528
rect 219250 3516 219256 3528
rect 218204 3488 219256 3516
rect 218204 3476 218210 3488
rect 219250 3476 219256 3488
rect 219308 3476 219314 3528
rect 222930 3476 222936 3528
rect 222988 3516 222994 3528
rect 223482 3516 223488 3528
rect 222988 3488 223488 3516
rect 222988 3476 222994 3488
rect 223482 3476 223488 3488
rect 223540 3476 223546 3528
rect 224126 3476 224132 3528
rect 224184 3516 224190 3528
rect 224862 3516 224868 3528
rect 224184 3488 224868 3516
rect 224184 3476 224190 3488
rect 224862 3476 224868 3488
rect 224920 3476 224926 3528
rect 225322 3476 225328 3528
rect 225380 3516 225386 3528
rect 226242 3516 226248 3528
rect 225380 3488 226248 3516
rect 225380 3476 225386 3488
rect 226242 3476 226248 3488
rect 226300 3476 226306 3528
rect 226518 3476 226524 3528
rect 226576 3516 226582 3528
rect 227622 3516 227628 3528
rect 226576 3488 227628 3516
rect 226576 3476 226582 3488
rect 227622 3476 227628 3488
rect 227680 3476 227686 3528
rect 231302 3476 231308 3528
rect 231360 3516 231366 3528
rect 231762 3516 231768 3528
rect 231360 3488 231768 3516
rect 231360 3476 231366 3488
rect 231762 3476 231768 3488
rect 231820 3476 231826 3528
rect 232498 3476 232504 3528
rect 232556 3516 232562 3528
rect 233142 3516 233148 3528
rect 232556 3488 233148 3516
rect 232556 3476 232562 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 233694 3476 233700 3528
rect 233752 3516 233758 3528
rect 234522 3516 234528 3528
rect 233752 3488 234528 3516
rect 233752 3476 233758 3488
rect 234522 3476 234528 3488
rect 234580 3476 234586 3528
rect 239582 3476 239588 3528
rect 239640 3516 239646 3528
rect 240042 3516 240048 3528
rect 239640 3488 240048 3516
rect 239640 3476 239646 3488
rect 240042 3476 240048 3488
rect 240100 3476 240106 3528
rect 240778 3476 240784 3528
rect 240836 3516 240842 3528
rect 241422 3516 241428 3528
rect 240836 3488 241428 3516
rect 240836 3476 240842 3488
rect 241422 3476 241428 3488
rect 241480 3476 241486 3528
rect 243170 3476 243176 3528
rect 243228 3516 243234 3528
rect 244182 3516 244188 3528
rect 243228 3488 244188 3516
rect 243228 3476 243234 3488
rect 244182 3476 244188 3488
rect 244240 3476 244246 3528
rect 249150 3476 249156 3528
rect 249208 3516 249214 3528
rect 249702 3516 249708 3528
rect 249208 3488 249708 3516
rect 249208 3476 249214 3488
rect 249702 3476 249708 3488
rect 249760 3476 249766 3528
rect 251450 3476 251456 3528
rect 251508 3516 251514 3528
rect 252462 3516 252468 3528
rect 251508 3488 252468 3516
rect 251508 3476 251514 3488
rect 252462 3476 252468 3488
rect 252520 3476 252526 3528
rect 257430 3476 257436 3528
rect 257488 3516 257494 3528
rect 257982 3516 257988 3528
rect 257488 3488 257988 3516
rect 257488 3476 257494 3488
rect 257982 3476 257988 3488
rect 258040 3476 258046 3528
rect 258626 3476 258632 3528
rect 258684 3516 258690 3528
rect 259362 3516 259368 3528
rect 258684 3488 259368 3516
rect 258684 3476 258690 3488
rect 259362 3476 259368 3488
rect 259420 3476 259426 3528
rect 262214 3476 262220 3528
rect 262272 3516 262278 3528
rect 263686 3516 263692 3528
rect 262272 3488 263692 3516
rect 262272 3476 262278 3488
rect 263686 3476 263692 3488
rect 263744 3476 263750 3528
rect 265802 3476 265808 3528
rect 265860 3516 265866 3528
rect 266262 3516 266268 3528
rect 265860 3488 266268 3516
rect 265860 3476 265866 3488
rect 266262 3476 266268 3488
rect 266320 3476 266326 3528
rect 268102 3476 268108 3528
rect 268160 3516 268166 3528
rect 269022 3516 269028 3528
rect 268160 3488 269028 3516
rect 268160 3476 268166 3488
rect 269022 3476 269028 3488
rect 269080 3476 269086 3528
rect 269298 3476 269304 3528
rect 269356 3516 269362 3528
rect 270402 3516 270408 3528
rect 269356 3488 270408 3516
rect 269356 3476 269362 3488
rect 270402 3476 270408 3488
rect 270460 3476 270466 3528
rect 272886 3476 272892 3528
rect 272944 3516 272950 3528
rect 273346 3516 273352 3528
rect 272944 3488 273352 3516
rect 272944 3476 272950 3488
rect 273346 3476 273352 3488
rect 273404 3476 273410 3528
rect 276014 3476 276020 3528
rect 276072 3516 276078 3528
rect 276474 3516 276480 3528
rect 276072 3488 276480 3516
rect 276072 3476 276078 3488
rect 276474 3476 276480 3488
rect 276532 3476 276538 3528
rect 281534 3476 281540 3528
rect 281592 3516 281598 3528
rect 282454 3516 282460 3528
rect 281592 3488 282460 3516
rect 281592 3476 281598 3488
rect 282454 3476 282460 3488
rect 282512 3476 282518 3528
rect 291102 3476 291108 3528
rect 291160 3516 291166 3528
rect 291930 3516 291936 3528
rect 291160 3488 291936 3516
rect 291160 3476 291166 3488
rect 291930 3476 291936 3488
rect 291988 3476 291994 3528
rect 292482 3476 292488 3528
rect 292540 3516 292546 3528
rect 294322 3516 294328 3528
rect 292540 3488 294328 3516
rect 292540 3476 292546 3488
rect 294322 3476 294328 3488
rect 294380 3476 294386 3528
rect 298002 3476 298008 3528
rect 298060 3516 298066 3528
rect 300302 3516 300308 3528
rect 298060 3488 300308 3516
rect 298060 3476 298066 3488
rect 300302 3476 300308 3488
rect 300360 3476 300366 3528
rect 302142 3476 302148 3528
rect 302200 3516 302206 3528
rect 304994 3516 305000 3528
rect 302200 3488 305000 3516
rect 302200 3476 302206 3488
rect 304994 3476 305000 3488
rect 305052 3476 305058 3528
rect 309042 3476 309048 3528
rect 309100 3516 309106 3528
rect 313366 3516 313372 3528
rect 309100 3488 313372 3516
rect 309100 3476 309106 3488
rect 313366 3476 313372 3488
rect 313424 3476 313430 3528
rect 317322 3476 317328 3528
rect 317380 3516 317386 3528
rect 322842 3516 322848 3528
rect 317380 3488 322848 3516
rect 317380 3476 317386 3488
rect 322842 3476 322848 3488
rect 322900 3476 322906 3528
rect 331030 3476 331036 3528
rect 331088 3516 331094 3528
rect 339494 3516 339500 3528
rect 331088 3488 339500 3516
rect 331088 3476 331094 3488
rect 339494 3476 339500 3488
rect 339552 3476 339558 3528
rect 346210 3476 346216 3528
rect 346268 3516 346274 3528
rect 357342 3516 357348 3528
rect 346268 3488 357348 3516
rect 346268 3476 346274 3488
rect 357342 3476 357348 3488
rect 357400 3476 357406 3528
rect 358722 3476 358728 3528
rect 358780 3516 358786 3528
rect 371602 3516 371608 3528
rect 358780 3488 371608 3516
rect 358780 3476 358786 3488
rect 371602 3476 371608 3488
rect 371660 3476 371666 3528
rect 373810 3476 373816 3528
rect 373868 3516 373874 3528
rect 389450 3516 389456 3528
rect 373868 3488 389456 3516
rect 373868 3476 373874 3488
rect 389450 3476 389456 3488
rect 389508 3476 389514 3528
rect 393130 3476 393136 3528
rect 393188 3516 393194 3528
rect 412082 3516 412088 3528
rect 393188 3488 412088 3516
rect 393188 3476 393194 3488
rect 412082 3476 412088 3488
rect 412140 3476 412146 3528
rect 416590 3476 416596 3528
rect 416648 3516 416654 3528
rect 439406 3516 439412 3528
rect 416648 3488 439412 3516
rect 416648 3476 416654 3488
rect 439406 3476 439412 3488
rect 439464 3476 439470 3528
rect 440142 3476 440148 3528
rect 440200 3516 440206 3528
rect 466822 3516 466828 3528
rect 440200 3488 466828 3516
rect 440200 3476 440206 3488
rect 466822 3476 466828 3488
rect 466880 3476 466886 3528
rect 467926 3476 467932 3528
rect 467984 3516 467990 3528
rect 469122 3516 469128 3528
rect 467984 3488 469128 3516
rect 467984 3476 467990 3488
rect 469122 3476 469128 3488
rect 469180 3476 469186 3528
rect 469232 3516 469260 3556
rect 469306 3544 469312 3596
rect 469364 3584 469370 3596
rect 492950 3584 492956 3596
rect 469364 3556 492956 3584
rect 469364 3544 469370 3556
rect 492950 3544 492956 3556
rect 493008 3544 493014 3596
rect 495342 3544 495348 3596
rect 495400 3584 495406 3596
rect 531038 3584 531044 3596
rect 495400 3556 531044 3584
rect 495400 3544 495406 3556
rect 531038 3544 531044 3556
rect 531096 3544 531102 3596
rect 532602 3544 532608 3596
rect 532660 3584 532666 3596
rect 573818 3584 573824 3596
rect 532660 3556 573824 3584
rect 532660 3544 532666 3556
rect 573818 3544 573824 3556
rect 573876 3544 573882 3596
rect 498930 3516 498936 3528
rect 469232 3488 498936 3516
rect 498930 3476 498936 3488
rect 498988 3476 498994 3528
rect 499390 3476 499396 3528
rect 499448 3516 499454 3528
rect 535730 3516 535736 3528
rect 499448 3488 535736 3516
rect 499448 3476 499454 3488
rect 535730 3476 535736 3488
rect 535788 3476 535794 3528
rect 536742 3476 536748 3528
rect 536800 3516 536806 3528
rect 578602 3516 578608 3528
rect 536800 3488 578608 3516
rect 536800 3476 536806 3488
rect 578602 3476 578608 3488
rect 578660 3476 578666 3528
rect 164694 3408 164700 3460
rect 164752 3448 164758 3460
rect 165522 3448 165528 3460
rect 164752 3420 165528 3448
rect 164752 3408 164758 3420
rect 165522 3408 165528 3420
rect 165580 3408 165586 3460
rect 241974 3408 241980 3460
rect 242032 3448 242038 3460
rect 242802 3448 242808 3460
rect 242032 3420 242808 3448
rect 242032 3408 242038 3420
rect 242802 3408 242808 3420
rect 242860 3408 242866 3460
rect 250346 3408 250352 3460
rect 250404 3448 250410 3460
rect 251082 3448 251088 3460
rect 250404 3420 251088 3448
rect 250404 3408 250410 3420
rect 251082 3408 251088 3420
rect 251140 3408 251146 3460
rect 295242 3408 295248 3460
rect 295300 3448 295306 3460
rect 297910 3448 297916 3460
rect 295300 3420 297916 3448
rect 295300 3408 295306 3420
rect 297910 3408 297916 3420
rect 297968 3408 297974 3460
rect 300762 3408 300768 3460
rect 300820 3448 300826 3460
rect 303798 3448 303804 3460
rect 300820 3420 303804 3448
rect 300820 3408 300826 3420
rect 303798 3408 303804 3420
rect 303856 3408 303862 3460
rect 306190 3408 306196 3460
rect 306248 3448 306254 3460
rect 310974 3448 310980 3460
rect 306248 3420 310980 3448
rect 306248 3408 306254 3420
rect 310974 3408 310980 3420
rect 311032 3408 311038 3460
rect 315942 3408 315948 3460
rect 316000 3448 316006 3460
rect 321646 3448 321652 3460
rect 316000 3420 321652 3448
rect 316000 3408 316006 3420
rect 321646 3408 321652 3420
rect 321704 3408 321710 3460
rect 322750 3408 322756 3460
rect 322808 3448 322814 3460
rect 330018 3448 330024 3460
rect 322808 3420 330024 3448
rect 322808 3408 322814 3420
rect 330018 3408 330024 3420
rect 330076 3408 330082 3460
rect 338022 3408 338028 3460
rect 338080 3448 338086 3460
rect 347866 3448 347872 3460
rect 338080 3420 347872 3448
rect 338080 3408 338086 3420
rect 347866 3408 347872 3420
rect 347924 3408 347930 3460
rect 350442 3408 350448 3460
rect 350500 3448 350506 3460
rect 362126 3448 362132 3460
rect 350500 3420 362132 3448
rect 350500 3408 350506 3420
rect 362126 3408 362132 3420
rect 362184 3408 362190 3460
rect 365622 3408 365628 3460
rect 365680 3448 365686 3460
rect 379974 3448 379980 3460
rect 365680 3420 379980 3448
rect 365680 3408 365686 3420
rect 379974 3408 379980 3420
rect 380032 3408 380038 3460
rect 380710 3408 380716 3460
rect 380768 3448 380774 3460
rect 397822 3448 397828 3460
rect 380768 3420 397828 3448
rect 380768 3408 380774 3420
rect 397822 3408 397828 3420
rect 397880 3408 397886 3460
rect 404170 3408 404176 3460
rect 404228 3448 404234 3460
rect 425054 3448 425060 3460
rect 404228 3420 425060 3448
rect 404228 3408 404234 3420
rect 425054 3408 425060 3420
rect 425112 3408 425118 3460
rect 425146 3408 425152 3460
rect 425204 3448 425210 3460
rect 426342 3448 426348 3460
rect 425204 3420 426348 3448
rect 425204 3408 425210 3420
rect 426342 3408 426348 3420
rect 426400 3408 426406 3460
rect 426434 3408 426440 3460
rect 426492 3448 426498 3460
rect 450170 3448 450176 3460
rect 426492 3420 450176 3448
rect 426492 3408 426498 3420
rect 450170 3408 450176 3420
rect 450228 3408 450234 3460
rect 455322 3408 455328 3460
rect 455380 3448 455386 3460
rect 484578 3448 484584 3460
rect 455380 3420 484584 3448
rect 455380 3408 455386 3420
rect 484578 3408 484584 3420
rect 484636 3408 484642 3460
rect 492582 3408 492588 3460
rect 492640 3448 492646 3460
rect 527450 3448 527456 3460
rect 492640 3420 527456 3448
rect 492640 3408 492646 3420
rect 527450 3408 527456 3420
rect 527508 3408 527514 3460
rect 529658 3408 529664 3460
rect 529716 3448 529722 3460
rect 571426 3448 571432 3460
rect 529716 3420 571432 3448
rect 529716 3408 529722 3420
rect 571426 3408 571432 3420
rect 571484 3408 571490 3460
rect 150618 3380 150624 3392
rect 145576 3352 150624 3380
rect 150618 3340 150624 3352
rect 150676 3340 150682 3392
rect 170582 3340 170588 3392
rect 170640 3380 170646 3392
rect 171042 3380 171048 3392
rect 170640 3352 171048 3380
rect 170640 3340 170646 3352
rect 171042 3340 171048 3352
rect 171100 3340 171106 3392
rect 247954 3340 247960 3392
rect 248012 3380 248018 3392
rect 249058 3380 249064 3392
rect 248012 3352 249064 3380
rect 248012 3340 248018 3352
rect 249058 3340 249064 3352
rect 249116 3340 249122 3392
rect 310330 3340 310336 3392
rect 310388 3380 310394 3392
rect 315758 3380 315764 3392
rect 310388 3352 315764 3380
rect 310388 3340 310394 3352
rect 315758 3340 315764 3352
rect 315816 3340 315822 3392
rect 318610 3340 318616 3392
rect 318668 3380 318674 3392
rect 325234 3380 325240 3392
rect 318668 3352 325240 3380
rect 318668 3340 318674 3352
rect 325234 3340 325240 3352
rect 325292 3340 325298 3392
rect 326890 3340 326896 3392
rect 326948 3380 326954 3392
rect 333606 3380 333612 3392
rect 326948 3352 333612 3380
rect 326948 3340 326954 3352
rect 333606 3340 333612 3352
rect 333664 3340 333670 3392
rect 355962 3340 355968 3392
rect 356020 3380 356026 3392
rect 368014 3380 368020 3392
rect 356020 3352 368020 3380
rect 356020 3340 356026 3352
rect 368014 3340 368020 3352
rect 368072 3340 368078 3392
rect 369762 3340 369768 3392
rect 369820 3380 369826 3392
rect 384666 3380 384672 3392
rect 369820 3352 384672 3380
rect 369820 3340 369826 3352
rect 384666 3340 384672 3352
rect 384724 3340 384730 3392
rect 391842 3340 391848 3392
rect 391900 3380 391906 3392
rect 409690 3380 409696 3392
rect 391900 3352 409696 3380
rect 391900 3340 391906 3352
rect 409690 3340 409696 3352
rect 409748 3340 409754 3392
rect 412542 3340 412548 3392
rect 412600 3380 412606 3392
rect 422294 3380 422300 3392
rect 412600 3352 422300 3380
rect 412600 3340 412606 3352
rect 422294 3340 422300 3352
rect 422352 3340 422358 3392
rect 434714 3340 434720 3392
rect 434772 3380 434778 3392
rect 459646 3380 459652 3392
rect 434772 3352 459652 3380
rect 434772 3340 434778 3352
rect 459646 3340 459652 3352
rect 459704 3340 459710 3392
rect 463602 3340 463608 3392
rect 463660 3380 463666 3392
rect 469306 3380 469312 3392
rect 463660 3352 469312 3380
rect 463660 3340 463666 3352
rect 469306 3340 469312 3352
rect 469364 3340 469370 3392
rect 469398 3340 469404 3392
rect 469456 3380 469462 3392
rect 491754 3380 491760 3392
rect 469456 3352 491760 3380
rect 469456 3340 469462 3352
rect 491754 3340 491760 3352
rect 491812 3340 491818 3392
rect 496078 3340 496084 3392
rect 496136 3380 496142 3392
rect 507210 3380 507216 3392
rect 496136 3352 507216 3380
rect 496136 3340 496142 3352
rect 507210 3340 507216 3352
rect 507268 3340 507274 3392
rect 507302 3340 507308 3392
rect 507360 3380 507366 3392
rect 509602 3380 509608 3392
rect 507360 3352 509608 3380
rect 507360 3340 507366 3352
rect 509602 3340 509608 3352
rect 509660 3340 509666 3392
rect 511902 3340 511908 3392
rect 511960 3380 511966 3392
rect 550082 3380 550088 3392
rect 511960 3352 550088 3380
rect 511960 3340 511966 3352
rect 550082 3340 550088 3352
rect 550140 3340 550146 3392
rect 132678 3312 132684 3324
rect 132512 3284 132684 3312
rect 132678 3272 132684 3284
rect 132736 3272 132742 3324
rect 149238 3272 149244 3324
rect 149296 3312 149302 3324
rect 150342 3312 150348 3324
rect 149296 3284 150348 3312
rect 149296 3272 149302 3284
rect 150342 3272 150348 3284
rect 150400 3272 150406 3324
rect 157518 3272 157524 3324
rect 157576 3312 157582 3324
rect 158622 3312 158628 3324
rect 157576 3284 158628 3312
rect 157576 3272 157582 3284
rect 158622 3272 158628 3284
rect 158680 3272 158686 3324
rect 174170 3272 174176 3324
rect 174228 3312 174234 3324
rect 175182 3312 175188 3324
rect 174228 3284 175188 3312
rect 174228 3272 174234 3284
rect 175182 3272 175188 3284
rect 175240 3272 175246 3324
rect 234798 3272 234804 3324
rect 234856 3312 234862 3324
rect 235902 3312 235908 3324
rect 234856 3284 235908 3312
rect 234856 3272 234862 3284
rect 235902 3272 235908 3284
rect 235960 3272 235966 3324
rect 280154 3272 280160 3324
rect 280212 3312 280218 3324
rect 281258 3312 281264 3324
rect 280212 3284 281264 3312
rect 280212 3272 280218 3284
rect 281258 3272 281264 3284
rect 281316 3272 281322 3324
rect 310422 3272 310428 3324
rect 310480 3312 310486 3324
rect 314562 3312 314568 3324
rect 310480 3284 314568 3312
rect 310480 3272 310486 3284
rect 314562 3272 314568 3284
rect 314620 3272 314626 3324
rect 369670 3272 369676 3324
rect 369728 3312 369734 3324
rect 383562 3312 383568 3324
rect 369728 3284 383568 3312
rect 369728 3272 369734 3284
rect 383562 3272 383568 3284
rect 383620 3272 383626 3324
rect 389082 3272 389088 3324
rect 389140 3312 389146 3324
rect 406102 3312 406108 3324
rect 389140 3284 406108 3312
rect 389140 3272 389146 3284
rect 406102 3272 406108 3284
rect 406160 3272 406166 3324
rect 407022 3272 407028 3324
rect 407080 3312 407086 3324
rect 427538 3312 427544 3324
rect 407080 3284 427544 3312
rect 407080 3272 407086 3284
rect 427538 3272 427544 3284
rect 427596 3272 427602 3324
rect 434622 3312 434628 3324
rect 427648 3284 434628 3312
rect 235994 3204 236000 3256
rect 236052 3244 236058 3256
rect 237282 3244 237288 3256
rect 236052 3216 237288 3244
rect 236052 3204 236058 3216
rect 237282 3204 237288 3216
rect 237340 3204 237346 3256
rect 266998 3204 267004 3256
rect 267056 3244 267062 3256
rect 267826 3244 267832 3256
rect 267056 3216 267832 3244
rect 267056 3204 267062 3216
rect 267826 3204 267832 3216
rect 267884 3204 267890 3256
rect 274818 3204 274824 3256
rect 274876 3244 274882 3256
rect 275278 3244 275284 3256
rect 274876 3216 275284 3244
rect 274876 3204 274882 3216
rect 275278 3204 275284 3216
rect 275336 3204 275342 3256
rect 307662 3204 307668 3256
rect 307720 3244 307726 3256
rect 312170 3244 312176 3256
rect 307720 3216 312176 3244
rect 307720 3204 307726 3216
rect 312170 3204 312176 3216
rect 312228 3204 312234 3256
rect 364242 3204 364248 3256
rect 364300 3244 364306 3256
rect 377582 3244 377588 3256
rect 364300 3216 377588 3244
rect 364300 3204 364306 3216
rect 377582 3204 377588 3216
rect 377640 3204 377646 3256
rect 386322 3204 386328 3256
rect 386380 3244 386386 3256
rect 403710 3244 403716 3256
rect 386380 3216 403716 3244
rect 386380 3204 386386 3216
rect 403710 3204 403716 3216
rect 403768 3204 403774 3256
rect 404262 3204 404268 3256
rect 404320 3244 404326 3256
rect 423950 3244 423956 3256
rect 404320 3216 423956 3244
rect 404320 3204 404326 3216
rect 423950 3204 423956 3216
rect 424008 3204 424014 3256
rect 303522 3136 303528 3188
rect 303580 3176 303586 3188
rect 306190 3176 306196 3188
rect 303580 3148 306196 3176
rect 303580 3136 303586 3148
rect 306190 3136 306196 3148
rect 306248 3136 306254 3188
rect 361482 3136 361488 3188
rect 361540 3176 361546 3188
rect 373994 3176 374000 3188
rect 361540 3148 374000 3176
rect 361540 3136 361546 3148
rect 373994 3136 374000 3148
rect 374052 3136 374058 3188
rect 380802 3136 380808 3188
rect 380860 3176 380866 3188
rect 396626 3176 396632 3188
rect 380860 3148 396632 3176
rect 380860 3136 380866 3148
rect 396626 3136 396632 3148
rect 396684 3136 396690 3188
rect 398742 3136 398748 3188
rect 398800 3176 398806 3188
rect 417970 3176 417976 3188
rect 398800 3148 417976 3176
rect 398800 3136 398806 3148
rect 417970 3136 417976 3148
rect 418028 3136 418034 3188
rect 422294 3136 422300 3188
rect 422352 3176 422358 3188
rect 427648 3176 427676 3284
rect 434622 3272 434628 3284
rect 434680 3272 434686 3324
rect 437382 3272 437388 3324
rect 437440 3312 437446 3324
rect 463234 3312 463240 3324
rect 437440 3284 463240 3312
rect 437440 3272 437446 3284
rect 463234 3272 463240 3284
rect 463292 3272 463298 3324
rect 466362 3272 466368 3324
rect 466420 3312 466426 3324
rect 496538 3312 496544 3324
rect 466420 3284 496544 3312
rect 466420 3272 466426 3284
rect 496538 3272 496544 3284
rect 496596 3272 496602 3324
rect 502242 3272 502248 3324
rect 502300 3312 502306 3324
rect 538122 3312 538128 3324
rect 502300 3284 538128 3312
rect 502300 3272 502306 3284
rect 538122 3272 538128 3284
rect 538180 3272 538186 3324
rect 544378 3272 544384 3324
rect 544436 3312 544442 3324
rect 546494 3312 546500 3324
rect 544436 3284 546500 3312
rect 544436 3272 544442 3284
rect 546494 3272 546500 3284
rect 546552 3272 546558 3324
rect 546586 3272 546592 3324
rect 546644 3312 546650 3324
rect 577406 3312 577412 3324
rect 546644 3284 577412 3312
rect 546644 3272 546650 3284
rect 577406 3272 577412 3284
rect 577464 3272 577470 3324
rect 427722 3204 427728 3256
rect 427780 3244 427786 3256
rect 452470 3244 452476 3256
rect 427780 3216 452476 3244
rect 427780 3204 427786 3216
rect 452470 3204 452476 3216
rect 452528 3204 452534 3256
rect 452562 3204 452568 3256
rect 452620 3244 452626 3256
rect 481082 3244 481088 3256
rect 452620 3216 481088 3244
rect 452620 3204 452626 3216
rect 481082 3204 481088 3216
rect 481140 3204 481146 3256
rect 481542 3204 481548 3256
rect 481600 3244 481606 3256
rect 514386 3244 514392 3256
rect 481600 3216 514392 3244
rect 481600 3204 481606 3216
rect 514386 3204 514392 3216
rect 514444 3204 514450 3256
rect 514478 3204 514484 3256
rect 514536 3244 514542 3256
rect 520274 3244 520280 3256
rect 514536 3216 520280 3244
rect 514536 3204 514542 3216
rect 520274 3204 520280 3216
rect 520332 3204 520338 3256
rect 520366 3204 520372 3256
rect 520424 3244 520430 3256
rect 555970 3244 555976 3256
rect 520424 3216 555976 3244
rect 520424 3204 520430 3216
rect 555970 3204 555976 3216
rect 556028 3204 556034 3256
rect 422352 3148 427676 3176
rect 422352 3136 422358 3148
rect 436002 3136 436008 3188
rect 436060 3176 436066 3188
rect 460842 3176 460848 3188
rect 436060 3148 460848 3176
rect 436060 3136 436066 3148
rect 460842 3136 460848 3148
rect 460900 3136 460906 3188
rect 462222 3136 462228 3188
rect 462280 3176 462286 3188
rect 469398 3176 469404 3188
rect 462280 3148 469404 3176
rect 462280 3136 462286 3148
rect 469398 3136 469404 3148
rect 469456 3136 469462 3188
rect 469490 3136 469496 3188
rect 469548 3176 469554 3188
rect 495342 3176 495348 3188
rect 469548 3148 495348 3176
rect 469548 3136 469554 3148
rect 495342 3136 495348 3148
rect 495400 3136 495406 3188
rect 499482 3136 499488 3188
rect 499540 3176 499546 3188
rect 534534 3176 534540 3188
rect 499540 3148 534540 3176
rect 499540 3136 499546 3148
rect 534534 3136 534540 3148
rect 534592 3136 534598 3188
rect 537478 3136 537484 3188
rect 537536 3176 537542 3188
rect 570230 3176 570236 3188
rect 537536 3148 570236 3176
rect 537536 3136 537542 3148
rect 570230 3136 570236 3148
rect 570288 3136 570294 3188
rect 181346 3068 181352 3120
rect 181404 3108 181410 3120
rect 182082 3108 182088 3120
rect 181404 3080 182088 3108
rect 181404 3068 181410 3080
rect 182082 3068 182088 3080
rect 182140 3068 182146 3120
rect 376662 3068 376668 3120
rect 376720 3108 376726 3120
rect 391842 3108 391848 3120
rect 376720 3080 391848 3108
rect 376720 3068 376726 3080
rect 391842 3068 391848 3080
rect 391900 3068 391906 3120
rect 393222 3068 393228 3120
rect 393280 3108 393286 3120
rect 410886 3108 410892 3120
rect 393280 3080 410892 3108
rect 393280 3068 393286 3080
rect 410886 3068 410892 3080
rect 410944 3068 410950 3120
rect 422202 3068 422208 3120
rect 422260 3108 422266 3120
rect 445386 3108 445392 3120
rect 422260 3080 445392 3108
rect 422260 3068 422266 3080
rect 445386 3068 445392 3080
rect 445444 3068 445450 3120
rect 459370 3068 459376 3120
rect 459428 3108 459434 3120
rect 488166 3108 488172 3120
rect 459428 3080 488172 3108
rect 459428 3068 459434 3080
rect 488166 3068 488172 3080
rect 488224 3068 488230 3120
rect 493962 3068 493968 3120
rect 494020 3108 494026 3120
rect 528646 3108 528652 3120
rect 494020 3080 528652 3108
rect 494020 3068 494026 3080
rect 528646 3068 528652 3080
rect 528704 3068 528710 3120
rect 534718 3068 534724 3120
rect 534776 3108 534782 3120
rect 566734 3108 566740 3120
rect 534776 3080 566740 3108
rect 534776 3068 534782 3080
rect 566734 3068 566740 3080
rect 566792 3068 566798 3120
rect 18322 3000 18328 3052
rect 18380 3040 18386 3052
rect 19242 3040 19248 3052
rect 18380 3012 19248 3040
rect 18380 3000 18386 3012
rect 19242 3000 19248 3012
rect 19300 3000 19306 3052
rect 140866 3000 140872 3052
rect 140924 3040 140930 3052
rect 142062 3040 142068 3052
rect 140924 3012 142068 3040
rect 140924 3000 140930 3012
rect 142062 3000 142068 3012
rect 142120 3000 142126 3052
rect 175366 3000 175372 3052
rect 175424 3040 175430 3052
rect 176470 3040 176476 3052
rect 175424 3012 176476 3040
rect 175424 3000 175430 3012
rect 176470 3000 176476 3012
rect 176528 3000 176534 3052
rect 190822 3000 190828 3052
rect 190880 3040 190886 3052
rect 191742 3040 191748 3052
rect 190880 3012 191748 3040
rect 190880 3000 190886 3012
rect 191742 3000 191748 3012
rect 191800 3000 191806 3052
rect 206278 3000 206284 3052
rect 206336 3040 206342 3052
rect 206922 3040 206928 3052
rect 206336 3012 206928 3040
rect 206336 3000 206342 3012
rect 206922 3000 206928 3012
rect 206980 3000 206986 3052
rect 259822 3000 259828 3052
rect 259880 3040 259886 3052
rect 260742 3040 260748 3052
rect 259880 3012 260748 3040
rect 259880 3000 259886 3012
rect 260742 3000 260748 3012
rect 260800 3000 260806 3052
rect 261018 3000 261024 3052
rect 261076 3040 261082 3052
rect 262122 3040 262128 3052
rect 261076 3012 262128 3040
rect 261076 3000 261082 3012
rect 262122 3000 262128 3012
rect 262180 3000 262186 3052
rect 299382 3000 299388 3052
rect 299440 3040 299446 3052
rect 301406 3040 301412 3052
rect 299440 3012 301412 3040
rect 299440 3000 299446 3012
rect 301406 3000 301412 3012
rect 301464 3000 301470 3052
rect 311802 3000 311808 3052
rect 311860 3040 311866 3052
rect 316954 3040 316960 3052
rect 311860 3012 316960 3040
rect 311860 3000 311866 3012
rect 316954 3000 316960 3012
rect 317012 3000 317018 3052
rect 321462 3000 321468 3052
rect 321520 3040 321526 3052
rect 327626 3040 327632 3052
rect 321520 3012 327632 3040
rect 321520 3000 321526 3012
rect 327626 3000 327632 3012
rect 327684 3000 327690 3052
rect 384942 3000 384948 3052
rect 385000 3040 385006 3052
rect 402514 3040 402520 3052
rect 385000 3012 402520 3040
rect 385000 3000 385006 3012
rect 402514 3000 402520 3012
rect 402572 3000 402578 3052
rect 416682 3000 416688 3052
rect 416740 3040 416746 3052
rect 438210 3040 438216 3052
rect 416740 3012 438216 3040
rect 416740 3000 416746 3012
rect 438210 3000 438216 3012
rect 438268 3000 438274 3052
rect 452286 3000 452292 3052
rect 452344 3040 452350 3052
rect 479886 3040 479892 3052
rect 452344 3012 479892 3040
rect 452344 3000 452350 3012
rect 479886 3000 479892 3012
rect 479944 3000 479950 3052
rect 483658 3000 483664 3052
rect 483716 3040 483722 3052
rect 503622 3040 503628 3052
rect 483716 3012 503628 3040
rect 483716 3000 483722 3012
rect 503622 3000 503628 3012
rect 503680 3000 503686 3052
rect 512638 3000 512644 3052
rect 512696 3040 512702 3052
rect 517882 3040 517888 3052
rect 512696 3012 517888 3040
rect 512696 3000 512702 3012
rect 517882 3000 517888 3012
rect 517940 3000 517946 3052
rect 521102 3000 521108 3052
rect 521160 3040 521166 3052
rect 525058 3040 525064 3052
rect 521160 3012 525064 3040
rect 521160 3000 521166 3012
rect 525058 3000 525064 3012
rect 525116 3000 525122 3052
rect 526438 3000 526444 3052
rect 526496 3040 526502 3052
rect 559558 3040 559564 3052
rect 526496 3012 559564 3040
rect 526496 3000 526502 3012
rect 559558 3000 559564 3012
rect 559616 3000 559622 3052
rect 291010 2932 291016 2984
rect 291068 2972 291074 2984
rect 293126 2972 293132 2984
rect 291068 2944 293132 2972
rect 291068 2932 291074 2944
rect 293126 2932 293132 2944
rect 293184 2932 293190 2984
rect 299290 2932 299296 2984
rect 299348 2972 299354 2984
rect 302602 2972 302608 2984
rect 299348 2944 302608 2972
rect 299348 2932 299354 2944
rect 302602 2932 302608 2944
rect 302660 2932 302666 2984
rect 329742 2932 329748 2984
rect 329800 2972 329806 2984
rect 337102 2972 337108 2984
rect 329800 2944 337108 2972
rect 329800 2932 329806 2944
rect 337102 2932 337108 2944
rect 337160 2932 337166 2984
rect 384850 2932 384856 2984
rect 384908 2972 384914 2984
rect 401318 2972 401324 2984
rect 384908 2944 401324 2972
rect 384908 2932 384914 2944
rect 401318 2932 401324 2944
rect 401376 2932 401382 2984
rect 451182 2932 451188 2984
rect 451240 2972 451246 2984
rect 478690 2972 478696 2984
rect 451240 2944 478696 2972
rect 451240 2932 451246 2944
rect 478690 2932 478696 2944
rect 478748 2932 478754 2984
rect 516870 2932 516876 2984
rect 516928 2972 516934 2984
rect 528462 2972 528468 2984
rect 516928 2944 528468 2972
rect 516928 2932 516934 2944
rect 528462 2932 528468 2944
rect 528520 2932 528526 2984
rect 540238 2932 540244 2984
rect 540296 2972 540302 2984
rect 546586 2972 546592 2984
rect 540296 2944 546592 2972
rect 540296 2932 540302 2944
rect 546586 2932 546592 2944
rect 546644 2932 546650 2984
rect 552658 2972 552664 2984
rect 546696 2944 552664 2972
rect 274082 2864 274088 2916
rect 274140 2904 274146 2916
rect 274542 2904 274548 2916
rect 274140 2876 274548 2904
rect 274140 2864 274146 2876
rect 274542 2864 274548 2876
rect 274600 2864 274606 2916
rect 318702 2864 318708 2916
rect 318760 2904 318766 2916
rect 324038 2904 324044 2916
rect 318760 2876 324044 2904
rect 318760 2864 318766 2876
rect 324038 2864 324044 2876
rect 324096 2864 324102 2916
rect 326982 2864 326988 2916
rect 327040 2904 327046 2916
rect 334710 2904 334716 2916
rect 327040 2876 334716 2904
rect 327040 2864 327046 2876
rect 334710 2864 334716 2876
rect 334768 2864 334774 2916
rect 448422 2864 448428 2916
rect 448480 2904 448486 2916
rect 475102 2904 475108 2916
rect 448480 2876 475108 2904
rect 448480 2864 448486 2876
rect 475102 2864 475108 2876
rect 475160 2864 475166 2916
rect 514846 2864 514852 2916
rect 514904 2904 514910 2916
rect 528370 2904 528376 2916
rect 514904 2876 528376 2904
rect 514904 2864 514910 2876
rect 528370 2864 528376 2876
rect 528428 2864 528434 2916
rect 529198 2864 529204 2916
rect 529256 2904 529262 2916
rect 532234 2904 532240 2916
rect 529256 2876 532240 2904
rect 529256 2864 529262 2876
rect 532234 2864 532240 2876
rect 532292 2864 532298 2916
rect 541618 2864 541624 2916
rect 541676 2904 541682 2916
rect 546696 2904 546724 2944
rect 552658 2932 552664 2944
rect 552716 2932 552722 2984
rect 567838 2972 567844 2984
rect 552768 2944 567844 2972
rect 541676 2876 546724 2904
rect 541676 2864 541682 2876
rect 547230 2864 547236 2916
rect 547288 2904 547294 2916
rect 552768 2904 552796 2944
rect 567838 2932 567844 2944
rect 567896 2932 567902 2984
rect 547288 2876 552796 2904
rect 547288 2864 547294 2876
rect 118234 2796 118240 2848
rect 118292 2836 118298 2848
rect 118602 2836 118608 2848
rect 118292 2808 118608 2836
rect 118292 2796 118298 2808
rect 118602 2796 118608 2808
rect 118660 2796 118666 2848
rect 444282 2796 444288 2848
rect 444340 2836 444346 2848
rect 470318 2836 470324 2848
rect 444340 2808 470324 2836
rect 444340 2796 444346 2808
rect 470318 2796 470324 2808
rect 470376 2796 470382 2848
rect 545758 2796 545764 2848
rect 545816 2836 545822 2848
rect 553578 2836 553584 2848
rect 545816 2808 553584 2836
rect 545816 2796 545822 2808
rect 553578 2796 553584 2808
rect 553636 2796 553642 2848
rect 109954 552 109960 604
rect 110012 592 110018 604
rect 110322 592 110328 604
rect 110012 564 110328 592
rect 110012 552 110018 564
rect 110322 552 110328 564
rect 110380 552 110386 604
rect 418246 552 418252 604
rect 418304 592 418310 604
rect 419166 592 419172 604
rect 418304 564 419172 592
rect 418304 552 418310 564
rect 419166 552 419172 564
rect 419224 552 419230 604
rect 429194 552 429200 604
rect 429252 592 429258 604
rect 429930 592 429936 604
rect 429252 564 429936 592
rect 429252 552 429258 564
rect 429930 552 429936 564
rect 429988 552 429994 604
rect 436186 552 436192 604
rect 436244 592 436250 604
rect 437014 592 437020 604
rect 436244 564 437020 592
rect 436244 552 436250 564
rect 437014 552 437020 564
rect 437072 552 437078 604
rect 447134 552 447140 604
rect 447192 592 447198 604
rect 447778 592 447784 604
rect 447192 564 447784 592
rect 447192 552 447198 564
rect 447778 552 447784 564
rect 447836 552 447842 604
rect 454218 552 454224 604
rect 454276 592 454282 604
rect 454862 592 454868 604
rect 454276 564 454868 592
rect 454276 552 454282 564
rect 454862 552 454868 564
rect 454920 552 454926 604
rect 461026 552 461032 604
rect 461084 592 461090 604
rect 462038 592 462044 604
rect 461084 564 462044 592
rect 461084 552 461090 564
rect 462038 552 462044 564
rect 462096 552 462102 604
rect 472066 552 472072 604
rect 472124 592 472130 604
rect 472710 592 472716 604
rect 472124 564 472716 592
rect 472124 552 472130 564
rect 472710 552 472716 564
rect 472768 552 472774 604
rect 485866 552 485872 604
rect 485924 592 485930 604
rect 486970 592 486976 604
rect 485924 564 486976 592
rect 485924 552 485930 564
rect 486970 552 486976 564
rect 487028 552 487034 604
rect 489914 552 489920 604
rect 489972 592 489978 604
rect 490558 592 490564 604
rect 489972 564 490564 592
rect 489972 552 489978 564
rect 490558 552 490564 564
rect 490616 552 490622 604
rect 496814 552 496820 604
rect 496872 592 496878 604
rect 497734 592 497740 604
rect 496872 564 497740 592
rect 496872 552 496878 564
rect 497734 552 497740 564
rect 497792 552 497798 604
rect 525794 552 525800 604
rect 525852 592 525858 604
rect 526254 592 526260 604
rect 525852 564 526260 592
rect 525852 552 525858 564
rect 526254 552 526260 564
rect 526312 552 526318 604
rect 538306 552 538312 604
rect 538364 592 538370 604
rect 539318 592 539324 604
rect 538364 564 539324 592
rect 538364 552 538370 564
rect 539318 552 539324 564
rect 539376 552 539382 604
rect 542354 552 542360 604
rect 542412 592 542418 604
rect 542906 592 542912 604
rect 542412 564 542912 592
rect 542412 552 542418 564
rect 542906 552 542912 564
rect 542964 552 542970 604
<< via1 >>
rect 154120 700952 154172 701004
rect 325700 700952 325752 701004
rect 137836 700884 137888 700936
rect 321560 700884 321612 700936
rect 256608 700816 256660 700868
rect 462320 700816 462372 700868
rect 262128 700748 262180 700800
rect 478512 700748 478564 700800
rect 89168 700680 89220 700732
rect 339500 700680 339552 700732
rect 72976 700612 73028 700664
rect 335360 700612 335412 700664
rect 244188 700544 244240 700596
rect 527180 700544 527232 700596
rect 248328 700476 248380 700528
rect 543464 700476 543516 700528
rect 40500 700408 40552 700460
rect 343640 700408 343692 700460
rect 24308 700340 24360 700392
rect 351920 700340 351972 700392
rect 8116 700272 8168 700324
rect 347780 700272 347832 700324
rect 274548 700204 274600 700256
rect 413652 700204 413704 700256
rect 270408 700136 270460 700188
rect 397460 700136 397512 700188
rect 202788 700068 202840 700120
rect 309140 700068 309192 700120
rect 218980 700000 219032 700052
rect 313280 700000 313332 700052
rect 288348 699932 288400 699984
rect 348792 699932 348844 699984
rect 284208 699864 284260 699916
rect 332508 699864 332560 699916
rect 267648 699796 267700 699848
rect 295340 699796 295392 699848
rect 283840 699728 283892 699780
rect 299480 699728 299532 699780
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 230388 696940 230440 696992
rect 580172 696940 580224 696992
rect 299572 692792 299624 692844
rect 300216 692792 300268 692844
rect 364340 692792 364392 692844
rect 365076 692792 365128 692844
rect 429200 692792 429252 692844
rect 429936 692792 429988 692844
rect 494060 692792 494112 692844
rect 494888 692792 494940 692844
rect 558920 692792 558972 692844
rect 559748 692792 559800 692844
rect 229100 690684 229152 690736
rect 230388 690684 230440 690736
rect 242900 690684 242952 690736
rect 244188 690684 244240 690736
rect 247040 690684 247092 690736
rect 248328 690684 248380 690736
rect 255320 690684 255372 690736
rect 256608 690684 256660 690736
rect 260840 690684 260892 690736
rect 262128 690684 262180 690736
rect 269120 690684 269172 690736
rect 270408 690684 270460 690736
rect 273260 690684 273312 690736
rect 274548 690684 274600 690736
rect 291936 688372 291988 688424
rect 299572 688372 299624 688424
rect 235908 688304 235960 688356
rect 304448 688304 304500 688356
rect 278688 688236 278740 688288
rect 364340 688236 364392 688288
rect 171048 688168 171100 688220
rect 317604 688168 317656 688220
rect 264980 688100 265032 688152
rect 429200 688100 429252 688152
rect 106188 688032 106240 688084
rect 330760 688032 330812 688084
rect 251180 687964 251232 688016
rect 494060 687964 494112 688016
rect 238760 687896 238812 687948
rect 558920 687896 558972 687948
rect 229008 687216 229060 687268
rect 230020 687216 230072 687268
rect 283196 687216 283248 687268
rect 284208 687216 284260 687268
rect 124220 687148 124272 687200
rect 379428 687148 379480 687200
rect 111800 687080 111852 687132
rect 365904 687080 365956 687132
rect 150440 687012 150492 687064
rect 411168 687012 411220 687064
rect 63868 686944 63920 686996
rect 229008 686944 229060 686996
rect 229100 686944 229152 686996
rect 229928 686944 229980 686996
rect 230020 686944 230072 686996
rect 233240 686944 233292 686996
rect 234620 686944 234672 686996
rect 580172 686944 580224 686996
rect 168380 686876 168432 686928
rect 539324 686876 539376 686928
rect 164240 686808 164292 686860
rect 540336 686808 540388 686860
rect 154580 686740 154632 686792
rect 541716 686740 541768 686792
rect 2872 686672 2924 686724
rect 405740 686672 405792 686724
rect 128360 686604 128412 686656
rect 539048 686604 539100 686656
rect 4988 686536 5040 686588
rect 418528 686536 418580 686588
rect 115940 686468 115992 686520
rect 538956 686468 539008 686520
rect 102140 686400 102192 686452
rect 538864 686400 538916 686452
rect 7564 686332 7616 686384
rect 444840 686332 444892 686384
rect 3056 686264 3108 686316
rect 440424 686264 440476 686316
rect 132500 686196 132552 686248
rect 577780 686196 577832 686248
rect 3240 686128 3292 686180
rect 453580 686128 453632 686180
rect 3332 686060 3384 686112
rect 471152 686060 471204 686112
rect 106280 685992 106332 686044
rect 577688 685992 577740 686044
rect 4068 685924 4120 685976
rect 484400 685924 484452 685976
rect 39856 685856 39908 685908
rect 49700 685856 49752 685908
rect 93860 685856 93912 685908
rect 577596 685856 577648 685908
rect 226156 685788 226208 685840
rect 540888 685788 540940 685840
rect 213000 685720 213052 685772
rect 540704 685720 540756 685772
rect 199844 685652 199896 685704
rect 540520 685652 540572 685704
rect 5540 685584 5592 685636
rect 357440 685584 357492 685636
rect 186688 685516 186740 685568
rect 539508 685516 539560 685568
rect 217416 685448 217468 685500
rect 578148 685448 578200 685500
rect 6736 685380 6788 685432
rect 370228 685380 370280 685432
rect 173532 685312 173584 685364
rect 539416 685312 539468 685364
rect 204168 685244 204220 685296
rect 578056 685244 578108 685296
rect 6644 685176 6696 685228
rect 383752 685176 383804 685228
rect 411168 685176 411220 685228
rect 579988 685176 580040 685228
rect 191012 685108 191064 685160
rect 577964 685108 578016 685160
rect 25596 685040 25648 685092
rect 414112 685040 414164 685092
rect 6552 684972 6604 685024
rect 396540 684972 396592 685024
rect 147220 684904 147272 684956
rect 541624 684904 541676 684956
rect 177856 684836 177908 684888
rect 579804 684836 579856 684888
rect 6460 684768 6512 684820
rect 409880 684768 409932 684820
rect 6368 684700 6420 684752
rect 422852 684700 422904 684752
rect 160376 684632 160428 684684
rect 577872 684632 577924 684684
rect 25504 684564 25556 684616
rect 449164 684564 449216 684616
rect 6276 684496 6328 684548
rect 436100 684496 436152 684548
rect 221740 684428 221792 684480
rect 543096 684428 543148 684480
rect 38108 684360 38160 684412
rect 361580 684360 361632 684412
rect 398748 684360 398800 684412
rect 405648 684360 405700 684412
rect 418068 684360 418120 684412
rect 424968 684360 425020 684412
rect 437388 684360 437440 684412
rect 444288 684360 444340 684412
rect 456708 684360 456760 684412
rect 463608 684360 463660 684412
rect 33784 684292 33836 684344
rect 365812 684292 365864 684344
rect 365904 684292 365956 684344
rect 580908 684292 580960 684344
rect 208308 684224 208360 684276
rect 543004 684224 543056 684276
rect 38016 684156 38068 684208
rect 374644 684156 374696 684208
rect 379336 684156 379388 684208
rect 386328 684156 386380 684208
rect 476028 684156 476080 684208
rect 482928 684156 482980 684208
rect 195106 684088 195158 684140
rect 541808 684088 541860 684140
rect 39488 684020 39540 684072
rect 387800 684020 387852 684072
rect 495348 684020 495400 684072
rect 497924 684020 497976 684072
rect 39580 683952 39632 684004
rect 392216 683952 392268 684004
rect 37924 683884 37976 683936
rect 400956 683884 401008 683936
rect 5080 683816 5132 683868
rect 379060 683816 379112 683868
rect 379520 683816 379572 683868
rect 580172 683816 580224 683868
rect 32404 683748 32456 683800
rect 427268 683748 427320 683800
rect 142804 683680 142856 683732
rect 539140 683680 539192 683732
rect 182088 683612 182140 683664
rect 579896 683612 579948 683664
rect 138388 683544 138440 683596
rect 539232 683544 539284 683596
rect 2964 683476 3016 683528
rect 431868 683476 431920 683528
rect 29644 683408 29696 683460
rect 466736 683408 466788 683460
rect 3148 683340 3200 683392
rect 458180 683340 458232 683392
rect 4896 683272 4948 683324
rect 475476 683272 475528 683324
rect 521660 683272 521712 683324
rect 523776 683272 523828 683324
rect 89858 683204 89910 683256
rect 98598 683204 98650 683256
rect 580724 683204 580776 683256
rect 580540 683136 580592 683188
rect 2780 682252 2832 682304
rect 5540 682252 5592 682304
rect 540888 674772 540940 674824
rect 579712 674772 579764 674824
rect 2780 669264 2832 669316
rect 33784 669264 33836 669316
rect 2780 654032 2832 654084
rect 38108 654032 38160 654084
rect 578148 651312 578200 651364
rect 579620 651312 579672 651364
rect 543096 640228 543148 640280
rect 579712 640228 579764 640280
rect 540704 627852 540756 627904
rect 579712 627852 579764 627904
rect 2780 624860 2832 624912
rect 6736 624860 6788 624912
rect 2780 610444 2832 610496
rect 5080 610444 5132 610496
rect 578056 604392 578108 604444
rect 579620 604392 579672 604444
rect 2780 596096 2832 596148
rect 38016 596096 38068 596148
rect 543004 593308 543056 593360
rect 579712 593308 579764 593360
rect 540520 580932 540572 580984
rect 579712 580932 579764 580984
rect 2780 567332 2832 567384
rect 6644 567332 6696 567384
rect 577964 557336 578016 557388
rect 579620 557336 579672 557388
rect 2780 553324 2832 553376
rect 39580 553324 39632 553376
rect 541808 546388 541860 546440
rect 579712 546388 579764 546440
rect 2780 539520 2832 539572
rect 39488 539520 39540 539572
rect 539508 534012 539560 534064
rect 579712 534012 579764 534064
rect 2780 509940 2832 509992
rect 6552 509940 6604 509992
rect 539416 487092 539468 487144
rect 579896 487092 579948 487144
rect 2872 481584 2924 481636
rect 37924 481584 37976 481636
rect 540336 463632 540388 463684
rect 579896 463632 579948 463684
rect 539324 452548 539376 452600
rect 579896 452548 579948 452600
rect 2872 452412 2924 452464
rect 6460 452412 6512 452464
rect 577872 440172 577924 440224
rect 579896 440172 579948 440224
rect 2780 438676 2832 438728
rect 4988 438676 5040 438728
rect 2872 425008 2924 425060
rect 25596 425008 25648 425060
rect 541716 405628 541768 405680
rect 579988 405628 580040 405680
rect 2872 395020 2924 395072
rect 6368 395020 6420 395072
rect 541624 393252 541676 393304
rect 579988 393252 580040 393304
rect 539232 369792 539284 369844
rect 579988 369792 580040 369844
rect 2964 367004 3016 367056
rect 32404 367004 32456 367056
rect 539140 358708 539192 358760
rect 579988 358708 580040 358760
rect 577780 346332 577832 346384
rect 579896 346332 579948 346384
rect 2964 337560 3016 337612
rect 6276 337560 6328 337612
rect 2964 323076 3016 323128
rect 7564 323076 7616 323128
rect 539048 311788 539100 311840
rect 580172 311788 580224 311840
rect 540796 299412 540848 299464
rect 580172 299412 580224 299464
rect 3056 295264 3108 295316
rect 25504 295264 25556 295316
rect 538956 264868 539008 264920
rect 580172 264868 580224 264920
rect 577688 252492 577740 252544
rect 579988 252492 580040 252544
rect 3148 251268 3200 251320
rect 6184 251268 6236 251320
rect 3332 223524 3384 223576
rect 29644 223524 29696 223576
rect 538864 217948 538916 218000
rect 580172 217948 580224 218000
rect 2780 208156 2832 208208
rect 4896 208156 4948 208208
rect 577596 205572 577648 205624
rect 580724 205572 580776 205624
rect 2780 179460 2832 179512
rect 4804 179460 4856 179512
rect 3148 165520 3200 165572
rect 39396 165520 39448 165572
rect 540612 158652 540664 158704
rect 580172 158652 580224 158704
rect 3332 136552 3384 136604
rect 22744 136552 22796 136604
rect 3332 122748 3384 122800
rect 24124 122748 24176 122800
rect 540428 111732 540480 111784
rect 580172 111732 580224 111784
rect 3332 79976 3384 80028
rect 39304 79976 39356 80028
rect 540244 64812 540296 64864
rect 580172 64812 580224 64864
rect 26148 62024 26200 62076
rect 61016 62024 61068 62076
rect 64788 62024 64840 62076
rect 93860 62024 93912 62076
rect 107476 62024 107528 62076
rect 131488 62024 131540 62076
rect 132408 62024 132460 62076
rect 151912 62024 151964 62076
rect 153108 62024 153160 62076
rect 170220 62024 170272 62076
rect 171048 62024 171100 62076
rect 185584 62024 185636 62076
rect 198648 62024 198700 62076
rect 209044 62024 209096 62076
rect 517796 62024 517848 62076
rect 518808 62024 518860 62076
rect 521936 62024 521988 62076
rect 522856 62024 522908 62076
rect 24768 61956 24820 62008
rect 60004 61956 60056 62008
rect 60648 61956 60700 62008
rect 90640 61956 90692 62008
rect 96528 61956 96580 62008
rect 121460 61956 121512 62008
rect 124128 61956 124180 62008
rect 144920 61956 144972 62008
rect 146208 61956 146260 62008
rect 164240 61956 164292 62008
rect 168288 61956 168340 62008
rect 183560 61956 183612 62008
rect 186228 61956 186280 62008
rect 198832 61956 198884 62008
rect 202696 61956 202748 62008
rect 212080 61956 212132 62008
rect 216588 61956 216640 62008
rect 224316 61956 224368 62008
rect 475016 61956 475068 62008
rect 496084 61956 496136 62008
rect 516784 61956 516836 62008
rect 519544 61956 519596 62008
rect 524972 61956 525024 62008
rect 531964 61956 532016 62008
rect 19248 61888 19300 61940
rect 55312 61888 55364 61940
rect 59912 61888 59964 61940
rect 67180 61888 67232 61940
rect 68928 61888 68980 61940
rect 98000 61888 98052 61940
rect 99288 61888 99340 61940
rect 124312 61888 124364 61940
rect 133788 61888 133840 61940
rect 153936 61888 153988 61940
rect 158628 61888 158680 61940
rect 174360 61888 174412 61940
rect 175188 61888 175240 61940
rect 188620 61888 188672 61940
rect 197268 61888 197320 61940
rect 208400 61888 208452 61940
rect 209688 61888 209740 61940
rect 218244 61888 218296 61940
rect 229008 61888 229060 61940
rect 235540 61888 235592 61940
rect 423956 61888 424008 61940
rect 447140 61888 447192 61940
rect 484124 61888 484176 61940
rect 512644 61888 512696 61940
rect 515772 61888 515824 61940
rect 522304 61888 522356 61940
rect 23388 61820 23440 61872
rect 59360 61820 59412 61872
rect 62028 61820 62080 61872
rect 91652 61820 91704 61872
rect 92388 61820 92440 61872
rect 118240 61820 118292 61872
rect 122748 61820 122800 61872
rect 143724 61820 143776 61872
rect 144828 61820 144880 61872
rect 163136 61820 163188 61872
rect 165528 61820 165580 61872
rect 180800 61820 180852 61872
rect 184848 61820 184900 61872
rect 197820 61820 197872 61872
rect 200028 61820 200080 61872
rect 210056 61820 210108 61872
rect 217968 61820 218020 61872
rect 225328 61820 225380 61872
rect 226248 61820 226300 61872
rect 232504 61820 232556 61872
rect 439228 61820 439280 61872
rect 465172 61820 465224 61872
rect 487068 61820 487120 61872
rect 516876 61820 516928 61872
rect 525708 61820 525760 61872
rect 534724 61820 534776 61872
rect 538036 61820 538088 61872
rect 541624 61820 541676 61872
rect 15108 61752 15160 61804
rect 51908 61752 51960 61804
rect 56508 61752 56560 61804
rect 87604 61752 87656 61804
rect 100668 61752 100720 61804
rect 125692 61752 125744 61804
rect 133696 61752 133748 61804
rect 153292 61752 153344 61804
rect 154488 61752 154540 61804
rect 171324 61752 171376 61804
rect 173808 61752 173860 61804
rect 187700 61752 187752 61804
rect 188988 61752 189040 61804
rect 200856 61752 200908 61804
rect 201408 61752 201460 61804
rect 211160 61752 211212 61804
rect 212448 61752 212500 61804
rect 221280 61752 221332 61804
rect 222108 61752 222160 61804
rect 229468 61752 229520 61804
rect 414756 61752 414808 61804
rect 436192 61752 436244 61804
rect 442356 61752 442408 61804
rect 467932 61752 467984 61804
rect 471888 61752 471940 61804
rect 483664 61752 483716 61804
rect 490288 61752 490340 61804
rect 520832 61752 520884 61804
rect 526996 61752 527048 61804
rect 547236 61752 547288 61804
rect 10968 61684 11020 61736
rect 47768 61684 47820 61736
rect 53748 61684 53800 61736
rect 84568 61684 84620 61736
rect 85488 61684 85540 61736
rect 112076 61684 112128 61736
rect 113088 61684 113140 61736
rect 135536 61684 135588 61736
rect 136548 61684 136600 61736
rect 155960 61684 156012 61736
rect 159916 61684 159968 61736
rect 175372 61684 175424 61736
rect 176476 61684 176528 61736
rect 189632 61684 189684 61736
rect 190368 61684 190420 61736
rect 201868 61684 201920 61736
rect 211068 61684 211120 61736
rect 219440 61684 219492 61736
rect 399484 61684 399536 61736
rect 418252 61684 418304 61736
rect 420828 61684 420880 61736
rect 443184 61684 443236 61736
rect 445392 61684 445444 61736
rect 472072 61684 472124 61736
rect 478052 61684 478104 61736
rect 508504 61684 508556 61736
rect 514668 61684 514720 61736
rect 545764 61684 545816 61736
rect 16488 61616 16540 61668
rect 52920 61616 52972 61668
rect 57888 61616 57940 61668
rect 88616 61616 88668 61668
rect 91008 61616 91060 61668
rect 116124 61616 116176 61668
rect 117228 61616 117280 61668
rect 139676 61616 139728 61668
rect 142068 61616 142120 61668
rect 160100 61616 160152 61668
rect 164148 61616 164200 61668
rect 179420 61616 179472 61668
rect 182088 61616 182140 61668
rect 194692 61616 194744 61668
rect 195888 61616 195940 61668
rect 207020 61616 207072 61668
rect 208308 61616 208360 61668
rect 217140 61616 217192 61668
rect 219256 61616 219308 61668
rect 226340 61616 226392 61668
rect 227628 61616 227680 61668
rect 233516 61616 233568 61668
rect 417792 61616 417844 61668
rect 440332 61616 440384 61668
rect 454592 61616 454644 61668
rect 483020 61616 483072 61668
rect 496452 61616 496504 61668
rect 529204 61616 529256 61668
rect 533160 61616 533212 61668
rect 547144 61616 547196 61668
rect 9588 61548 9640 61600
rect 46940 61548 46992 61600
rect 49608 61548 49660 61600
rect 81440 61548 81492 61600
rect 82636 61548 82688 61600
rect 109132 61548 109184 61600
rect 110328 61548 110380 61600
rect 133880 61548 133932 61600
rect 135168 61548 135220 61600
rect 154948 61548 155000 61600
rect 155868 61548 155920 61600
rect 172612 61548 172664 61600
rect 176568 61548 176620 61600
rect 190736 61548 190788 61600
rect 191748 61548 191800 61600
rect 202880 61548 202932 61600
rect 204168 61548 204220 61600
rect 214104 61548 214156 61600
rect 215208 61548 215260 61600
rect 223672 61548 223724 61600
rect 238668 61548 238720 61600
rect 243728 61548 243780 61600
rect 402520 61548 402572 61600
rect 422392 61548 422444 61600
rect 430120 61548 430172 61600
rect 454224 61548 454276 61600
rect 457628 61548 457680 61600
rect 485872 61548 485924 61600
rect 491208 61548 491260 61600
rect 525800 61548 525852 61600
rect 537208 61548 537260 61600
rect 567844 61548 567896 61600
rect 13636 61480 13688 61532
rect 51080 61480 51132 61532
rect 55128 61480 55180 61532
rect 85580 61480 85632 61532
rect 93768 61480 93820 61532
rect 119252 61480 119304 61532
rect 125416 61480 125468 61532
rect 146760 61480 146812 61532
rect 151636 61480 151688 61532
rect 169208 61480 169260 61532
rect 169668 61480 169720 61532
rect 184940 61480 184992 61532
rect 187608 61480 187660 61532
rect 200212 61480 200264 61532
rect 202788 61480 202840 61532
rect 213092 61480 213144 61532
rect 213828 61480 213880 61532
rect 222292 61480 222344 61532
rect 224868 61480 224920 61532
rect 231860 61480 231912 61532
rect 246948 61480 247000 61532
rect 251272 61480 251324 61532
rect 411720 61480 411772 61532
rect 433432 61480 433484 61532
rect 436008 61480 436060 61532
rect 461032 61480 461084 61532
rect 466828 61480 466880 61532
rect 496820 61480 496872 61532
rect 508688 61480 508740 61532
rect 544384 61480 544436 61532
rect 6828 61412 6880 61464
rect 44732 61412 44784 61464
rect 46848 61412 46900 61464
rect 74540 61412 74592 61464
rect 76564 61412 76616 61464
rect 79416 61412 79468 61464
rect 82728 61412 82780 61464
rect 110420 61412 110472 61464
rect 111708 61412 111760 61464
rect 134524 61412 134576 61464
rect 137928 61412 137980 61464
rect 157340 61412 157392 61464
rect 160008 61412 160060 61464
rect 176752 61412 176804 61464
rect 177948 61412 178000 61464
rect 191840 61412 191892 61464
rect 193128 61412 193180 61464
rect 204260 61412 204312 61464
rect 205548 61412 205600 61464
rect 215300 61412 215352 61464
rect 219348 61412 219400 61464
rect 227720 61412 227772 61464
rect 228916 61412 228968 61464
rect 234620 61412 234672 61464
rect 237288 61412 237340 61464
rect 241704 61412 241756 61464
rect 405556 61412 405608 61464
rect 425152 61412 425204 61464
rect 426992 61412 427044 61464
rect 451464 61412 451516 61464
rect 460664 61412 460716 61464
rect 489920 61412 489972 61464
rect 505560 61412 505612 61464
rect 542360 61412 542412 61464
rect 4068 61344 4120 61396
rect 42800 61344 42852 61396
rect 43444 61344 43496 61396
rect 48780 61344 48832 61396
rect 50988 61344 51040 61396
rect 82820 61344 82872 61396
rect 86868 61344 86920 61396
rect 113180 61344 113232 61396
rect 118608 61344 118660 61396
rect 140780 61344 140832 61396
rect 141976 61344 142028 61396
rect 161020 61344 161072 61396
rect 162768 61344 162820 61396
rect 178408 61344 178460 61396
rect 180708 61344 180760 61396
rect 193680 61344 193732 61396
rect 194416 61344 194468 61396
rect 205916 61344 205968 61396
rect 210976 61344 211028 61396
rect 220268 61344 220320 61396
rect 237196 61344 237248 61396
rect 242900 61344 242952 61396
rect 408408 61344 408460 61396
rect 429200 61344 429252 61396
rect 433156 61344 433208 61396
rect 458364 61344 458416 61396
rect 463608 61344 463660 61396
rect 494244 61344 494296 61396
rect 502248 61344 502300 61396
rect 538312 61344 538364 61396
rect 539232 61344 539284 61396
rect 548524 61344 548576 61396
rect 31668 61276 31720 61328
rect 66260 61276 66312 61328
rect 67548 61276 67600 61328
rect 96804 61276 96856 61328
rect 97908 61276 97960 61328
rect 122288 61276 122340 61328
rect 125508 61276 125560 61328
rect 145748 61276 145800 61328
rect 148968 61276 149020 61328
rect 166172 61276 166224 61328
rect 168196 61276 168248 61328
rect 182456 61276 182508 61328
rect 183468 61276 183520 61328
rect 195980 61276 196032 61328
rect 206928 61276 206980 61328
rect 216128 61276 216180 61328
rect 28908 61208 28960 61260
rect 63500 61208 63552 61260
rect 64144 61208 64196 61260
rect 70400 61208 70452 61260
rect 73068 61208 73120 61260
rect 100852 61208 100904 61260
rect 104808 61208 104860 61260
rect 128360 61208 128412 61260
rect 129648 61208 129700 61260
rect 149796 61208 149848 61260
rect 150348 61208 150400 61260
rect 167184 61208 167236 61260
rect 172428 61208 172480 61260
rect 186596 61208 186648 61260
rect 194508 61208 194560 61260
rect 204904 61208 204956 61260
rect 520924 61208 520976 61260
rect 521568 61208 521620 61260
rect 33048 61140 33100 61192
rect 59912 61140 59964 61192
rect 71596 61140 71648 61192
rect 75368 61140 75420 61192
rect 75828 61140 75880 61192
rect 103888 61140 103940 61192
rect 107568 61140 107620 61192
rect 130476 61140 130528 61192
rect 139308 61140 139360 61192
rect 157984 61140 158036 61192
rect 161388 61140 161440 61192
rect 177396 61140 177448 61192
rect 179328 61140 179380 61192
rect 192668 61140 192720 61192
rect 39948 61072 40000 61124
rect 73344 61072 73396 61124
rect 75184 61072 75236 61124
rect 76380 61072 76432 61124
rect 78588 61072 78640 61124
rect 106280 61072 106332 61124
rect 114468 61072 114520 61124
rect 136640 61072 136692 61124
rect 143448 61072 143500 61124
rect 162124 61072 162176 61124
rect 166908 61072 166960 61124
rect 181444 61072 181496 61124
rect 184756 61072 184808 61124
rect 196808 61072 196860 61124
rect 233148 61072 233200 61124
rect 238760 61072 238812 61124
rect 245476 61072 245528 61124
rect 249800 61072 249852 61124
rect 256608 61072 256660 61124
rect 259000 61072 259052 61124
rect 497464 61072 497516 61124
rect 501604 61072 501656 61124
rect 38476 61004 38528 61056
rect 72240 61004 72292 61056
rect 75276 61004 75328 61056
rect 102876 61004 102928 61056
rect 103428 61004 103480 61056
rect 127348 61004 127400 61056
rect 140688 61004 140740 61056
rect 158996 61004 159048 61056
rect 223488 61004 223540 61056
rect 230480 61004 230532 61056
rect 234528 61004 234580 61056
rect 239680 61004 239732 61056
rect 241428 61004 241480 61056
rect 245752 61004 245804 61056
rect 257988 61004 258040 61056
rect 260012 61004 260064 61056
rect 535184 61004 535236 61056
rect 540244 61004 540296 61056
rect 35808 60936 35860 60988
rect 69204 60936 69256 60988
rect 42708 60868 42760 60920
rect 71596 60936 71648 60988
rect 71688 60936 71740 60988
rect 99840 60936 99892 60988
rect 117136 60936 117188 60988
rect 138572 60936 138624 60988
rect 151728 60936 151780 60988
rect 168380 60936 168432 60988
rect 235908 60936 235960 60988
rect 240692 60936 240744 60988
rect 245568 60936 245620 60988
rect 248788 60936 248840 60988
rect 251088 60936 251140 60988
rect 253940 60936 253992 60988
rect 255228 60936 255280 60988
rect 258172 60936 258224 60988
rect 74540 60868 74592 60920
rect 78772 60868 78824 60920
rect 79968 60868 80020 60920
rect 107016 60868 107068 60920
rect 115848 60868 115900 60920
rect 137560 60868 137612 60920
rect 147588 60868 147640 60920
rect 165160 60868 165212 60920
rect 242808 60868 242860 60920
rect 247132 60868 247184 60920
rect 249708 60868 249760 60920
rect 252928 60868 252980 60920
rect 253756 60868 253808 60920
rect 256976 60868 257028 60920
rect 529020 60868 529072 60920
rect 537484 60868 537536 60920
rect 40776 60800 40828 60852
rect 55956 60800 56008 60852
rect 68284 60800 68336 60852
rect 94688 60800 94740 60852
rect 119988 60800 120040 60852
rect 141700 60800 141752 60852
rect 157248 60800 157300 60852
rect 173348 60800 173400 60852
rect 231768 60800 231820 60852
rect 237564 60800 237616 60852
rect 240048 60800 240100 60852
rect 244740 60800 244792 60852
rect 252468 60800 252520 60852
rect 255320 60800 255372 60852
rect 260748 60800 260800 60852
rect 262220 60800 262272 60852
rect 264888 60800 264940 60852
rect 266360 60800 266412 60852
rect 503536 60800 503588 60852
rect 505744 60800 505796 60852
rect 512736 60800 512788 60852
rect 515404 60800 515456 60852
rect 519912 60800 519964 60852
rect 526444 60800 526496 60852
rect 531136 60800 531188 60852
rect 533344 60800 533396 60852
rect 47584 60732 47636 60784
rect 56968 60732 57020 60784
rect 60004 60732 60056 60784
rect 64236 60732 64288 60784
rect 89628 60732 89680 60784
rect 115112 60732 115164 60784
rect 121368 60732 121420 60784
rect 142712 60732 142764 60784
rect 220728 60732 220780 60784
rect 228364 60732 228416 60784
rect 230388 60732 230440 60784
rect 236552 60732 236604 60784
rect 244188 60732 244240 60784
rect 247776 60732 247828 60784
rect 249064 60732 249116 60784
rect 251916 60732 251968 60784
rect 253848 60732 253900 60784
rect 255964 60732 256016 60784
rect 259368 60732 259420 60784
rect 261024 60732 261076 60784
rect 262128 60732 262180 60784
rect 263140 60732 263192 60784
rect 263508 60732 263560 60784
rect 265164 60732 265216 60784
rect 266268 60732 266320 60784
rect 267188 60732 267240 60784
rect 286232 60732 286284 60784
rect 286968 60732 287020 60784
rect 289268 60732 289320 60784
rect 290004 60732 290056 60784
rect 290280 60732 290332 60784
rect 291108 60732 291160 60784
rect 293316 60732 293368 60784
rect 293868 60732 293920 60784
rect 294328 60732 294380 60784
rect 295156 60732 295208 60784
rect 297456 60732 297508 60784
rect 298008 60732 298060 60784
rect 298468 60732 298520 60784
rect 299388 60732 299440 60784
rect 301504 60732 301556 60784
rect 302148 60732 302200 60784
rect 302516 60732 302568 60784
rect 303528 60732 303580 60784
rect 305552 60732 305604 60784
rect 306288 60732 306340 60784
rect 309692 60732 309744 60784
rect 310428 60732 310480 60784
rect 312728 60732 312780 60784
rect 313188 60732 313240 60784
rect 313740 60732 313792 60784
rect 314476 60732 314528 60784
rect 316776 60732 316828 60784
rect 317328 60732 317380 60784
rect 317788 60732 317840 60784
rect 318708 60732 318760 60784
rect 320916 60732 320968 60784
rect 321468 60732 321520 60784
rect 321928 60732 321980 60784
rect 322848 60732 322900 60784
rect 324964 60732 325016 60784
rect 325608 60732 325660 60784
rect 325976 60732 326028 60784
rect 326896 60732 326948 60784
rect 329012 60732 329064 60784
rect 329748 60732 329800 60784
rect 330116 60732 330168 60784
rect 331128 60732 331180 60784
rect 333152 60732 333204 60784
rect 333888 60732 333940 60784
rect 336188 60732 336240 60784
rect 336648 60732 336700 60784
rect 337200 60732 337252 60784
rect 337936 60732 337988 60784
rect 340328 60732 340380 60784
rect 340788 60732 340840 60784
rect 341340 60732 341392 60784
rect 342076 60732 342128 60784
rect 344376 60732 344428 60784
rect 344928 60732 344980 60784
rect 345388 60732 345440 60784
rect 346308 60732 346360 60784
rect 348424 60732 348476 60784
rect 349068 60732 349120 60784
rect 349436 60732 349488 60784
rect 350356 60732 350408 60784
rect 352564 60732 352616 60784
rect 353208 60732 353260 60784
rect 353576 60732 353628 60784
rect 354588 60732 354640 60784
rect 356612 60732 356664 60784
rect 357256 60732 357308 60784
rect 359648 60732 359700 60784
rect 360108 60732 360160 60784
rect 360660 60732 360712 60784
rect 361488 60732 361540 60784
rect 363788 60732 363840 60784
rect 364248 60732 364300 60784
rect 364800 60732 364852 60784
rect 365536 60732 365588 60784
rect 367836 60732 367888 60784
rect 368388 60732 368440 60784
rect 368848 60732 368900 60784
rect 369676 60732 369728 60784
rect 371884 60732 371936 60784
rect 372528 60732 372580 60784
rect 372896 60732 372948 60784
rect 373908 60732 373960 60784
rect 376024 60732 376076 60784
rect 376668 60732 376720 60784
rect 377036 60732 377088 60784
rect 377956 60732 378008 60784
rect 380072 60732 380124 60784
rect 380808 60732 380860 60784
rect 383108 60732 383160 60784
rect 383568 60732 383620 60784
rect 384120 60732 384172 60784
rect 384856 60732 384908 60784
rect 387248 60732 387300 60784
rect 387708 60732 387760 60784
rect 388260 60732 388312 60784
rect 389088 60732 389140 60784
rect 391296 60732 391348 60784
rect 391848 60732 391900 60784
rect 392308 60732 392360 60784
rect 393228 60732 393280 60784
rect 395344 60732 395396 60784
rect 395988 60732 396040 60784
rect 396448 60732 396500 60784
rect 397276 60732 397328 60784
rect 400496 60732 400548 60784
rect 401416 60732 401468 60784
rect 403532 60732 403584 60784
rect 404268 60732 404320 60784
rect 406568 60732 406620 60784
rect 407028 60732 407080 60784
rect 407672 60732 407724 60784
rect 408408 60732 408460 60784
rect 410708 60732 410760 60784
rect 411168 60732 411220 60784
rect 415768 60732 415820 60784
rect 416688 60732 416740 60784
rect 418896 60732 418948 60784
rect 419448 60732 419500 60784
rect 419908 60732 419960 60784
rect 420828 60732 420880 60784
rect 422944 60732 422996 60784
rect 423588 60732 423640 60784
rect 431132 60732 431184 60784
rect 431868 60732 431920 60784
rect 434168 60732 434220 60784
rect 434628 60732 434680 60784
rect 435180 60732 435232 60784
rect 436008 60732 436060 60784
rect 438216 60732 438268 60784
rect 438768 60732 438820 60784
rect 443368 60732 443420 60784
rect 444288 60732 444340 60784
rect 446404 60732 446456 60784
rect 447048 60732 447100 60784
rect 447416 60732 447468 60784
rect 448428 60732 448480 60784
rect 450452 60732 450504 60784
rect 451188 60732 451240 60784
rect 451556 60732 451608 60784
rect 452476 60732 452528 60784
rect 458640 60732 458692 60784
rect 459376 60732 459428 60784
rect 461676 60732 461728 60784
rect 462228 60732 462280 60784
rect 462780 60732 462832 60784
rect 463608 60732 463660 60784
rect 465816 60732 465868 60784
rect 466368 60732 466420 60784
rect 469864 60732 469916 60784
rect 470508 60732 470560 60784
rect 470876 60732 470928 60784
rect 471888 60732 471940 60784
rect 474004 60732 474056 60784
rect 474648 60732 474700 60784
rect 481088 60732 481140 60784
rect 481548 60732 481600 60784
rect 482100 60732 482152 60784
rect 482836 60732 482888 60784
rect 485228 60732 485280 60784
rect 485688 60732 485740 60784
rect 486240 60732 486292 60784
rect 487068 60732 487120 60784
rect 489276 60732 489328 60784
rect 489828 60732 489880 60784
rect 493324 60732 493376 60784
rect 493968 60732 494020 60784
rect 494336 60732 494388 60784
rect 495256 60732 495308 60784
rect 498476 60732 498528 60784
rect 499488 60732 499540 60784
rect 501512 60732 501564 60784
rect 502248 60732 502300 60784
rect 504548 60732 504600 60784
rect 505008 60732 505060 60784
rect 506388 60732 506440 60784
rect 507124 60732 507176 60784
rect 509700 60732 509752 60784
rect 511264 60732 511316 60784
rect 513748 60732 513800 60784
rect 514668 60732 514720 60784
rect 528008 60732 528060 60784
rect 528468 60732 528520 60784
rect 532148 60732 532200 60784
rect 532608 60732 532660 60784
rect 533988 60732 534040 60784
rect 536104 60732 536156 60784
rect 536196 60732 536248 60784
rect 536748 60732 536800 60784
rect 42892 60664 42944 60716
rect 43076 60664 43128 60716
rect 76564 60664 76616 60716
rect 76748 60664 76800 60716
rect 520832 60664 520884 60716
rect 520924 60596 520976 60648
rect 40132 59644 40184 59696
rect 40684 59644 40736 59696
rect 42800 57876 42852 57928
rect 43076 57876 43128 57928
rect 76472 57876 76524 57928
rect 76748 57876 76800 57928
rect 74540 56652 74592 56704
rect 75276 56652 75328 56704
rect 74632 56584 74684 56636
rect 74816 56584 74868 56636
rect 74264 56516 74316 56568
rect 74540 56516 74592 56568
rect 520740 53116 520792 53168
rect 520924 53116 520976 53168
rect 113456 51144 113508 51196
rect 516876 51144 516928 51196
rect 113456 51008 113508 51060
rect 516968 51008 517020 51060
rect 42800 48288 42852 48340
rect 42984 48288 43036 48340
rect 76472 48288 76524 48340
rect 76656 48288 76708 48340
rect 113272 48288 113324 48340
rect 113456 48288 113508 48340
rect 520740 48288 520792 48340
rect 520924 48288 520976 48340
rect 516692 48220 516744 48272
rect 516876 48220 516928 48272
rect 74264 46928 74316 46980
rect 74448 46928 74500 46980
rect 76656 41556 76708 41608
rect 42984 41420 43036 41472
rect 76656 41420 76708 41472
rect 113272 41420 113324 41472
rect 113364 41352 113416 41404
rect 577504 41352 577556 41404
rect 580540 41352 580592 41404
rect 42984 41284 43036 41336
rect 76656 38768 76708 38820
rect 42892 38632 42944 38684
rect 42984 38632 43036 38684
rect 76564 38632 76616 38684
rect 113180 38564 113232 38616
rect 113364 38564 113416 38616
rect 74356 37272 74408 37324
rect 74448 37272 74500 37324
rect 74356 37136 74408 37188
rect 74724 37136 74776 37188
rect 42892 33940 42944 33992
rect 43260 33940 43312 33992
rect 521016 31764 521068 31816
rect 516692 31696 516744 31748
rect 516876 31696 516928 31748
rect 521016 31628 521068 31680
rect 39856 30268 39908 30320
rect 579896 30268 579948 30320
rect 43076 28976 43128 29028
rect 43260 28976 43312 29028
rect 113180 28976 113232 29028
rect 113456 28976 113508 29028
rect 516600 28908 516652 28960
rect 516876 28908 516928 28960
rect 520924 28908 520976 28960
rect 521016 28908 521068 28960
rect 74264 27548 74316 27600
rect 74448 27548 74500 27600
rect 3516 22040 3568 22092
rect 538220 22040 538272 22092
rect 42892 19320 42944 19372
rect 42984 19320 43036 19372
rect 516600 19320 516652 19372
rect 516784 19320 516836 19372
rect 74080 17960 74132 18012
rect 74264 17960 74316 18012
rect 74080 9664 74132 9716
rect 74264 9664 74316 9716
rect 518716 6196 518768 6248
rect 558368 6196 558420 6248
rect 528468 6128 528520 6180
rect 569040 6128 569092 6180
rect 501604 5448 501656 5500
rect 533436 5448 533488 5500
rect 531964 5380 532016 5432
rect 565544 5380 565596 5432
rect 37372 5312 37424 5364
rect 70676 5312 70728 5364
rect 482836 5312 482888 5364
rect 515588 5312 515640 5364
rect 522304 5312 522356 5364
rect 554780 5312 554832 5364
rect 33876 5244 33928 5296
rect 67640 5244 67692 5296
rect 473268 5244 473320 5296
rect 504824 5244 504876 5296
rect 505744 5244 505796 5296
rect 540520 5244 540572 5296
rect 40960 5176 41012 5228
rect 74632 5176 74684 5228
rect 478788 5176 478840 5228
rect 512000 5176 512052 5228
rect 515404 5176 515456 5228
rect 551192 5176 551244 5228
rect 30288 5108 30340 5160
rect 64880 5108 64932 5160
rect 476028 5108 476080 5160
rect 508412 5108 508464 5160
rect 511264 5108 511316 5160
rect 547696 5108 547748 5160
rect 26700 5040 26752 5092
rect 62120 5040 62172 5092
rect 500868 5040 500920 5092
rect 536932 5040 536984 5092
rect 21916 4972 21968 5024
rect 57980 4972 58032 5024
rect 470508 4972 470560 5024
rect 501236 4972 501288 5024
rect 507124 4972 507176 5024
rect 544108 4972 544160 5024
rect 12440 4904 12492 4956
rect 49700 4904 49752 4956
rect 69480 4904 69532 4956
rect 98276 4904 98328 4956
rect 485688 4904 485740 4956
rect 519084 4904 519136 4956
rect 533344 4904 533396 4956
rect 572628 4904 572680 4956
rect 17224 4836 17276 4888
rect 53840 4836 53892 4888
rect 65984 4836 66036 4888
rect 95240 4836 95292 4888
rect 488448 4836 488500 4888
rect 522672 4836 522724 4888
rect 522856 4836 522908 4888
rect 561956 4836 562008 4888
rect 7656 4768 7708 4820
rect 45560 4768 45612 4820
rect 47400 4768 47452 4820
rect 77300 4768 77352 4820
rect 448336 4768 448388 4820
rect 476304 4768 476356 4820
rect 495256 4768 495308 4820
rect 529848 4768 529900 4820
rect 536104 4768 536156 4820
rect 576216 4768 576268 4820
rect 42156 4088 42208 4140
rect 42708 4088 42760 4140
rect 50528 4088 50580 4140
rect 50988 4088 51040 4140
rect 71872 4088 71924 4140
rect 73068 4088 73120 4140
rect 77852 4088 77904 4140
rect 78588 4088 78640 4140
rect 79048 4088 79100 4140
rect 79968 4088 80020 4140
rect 111156 4088 111208 4140
rect 111708 4088 111760 4140
rect 112352 4088 112404 4140
rect 113088 4088 113140 4140
rect 113548 4088 113600 4140
rect 114468 4088 114520 4140
rect 115940 4088 115992 4140
rect 117136 4088 117188 4140
rect 296628 4088 296680 4140
rect 299112 4088 299164 4140
rect 304908 4088 304960 4140
rect 308588 4088 308640 4140
rect 320088 4088 320140 4140
rect 326436 4088 326488 4140
rect 339408 4088 339460 4140
rect 348976 4088 349028 4140
rect 349068 4088 349120 4140
rect 359740 4088 359792 4140
rect 362868 4088 362920 4140
rect 376392 4088 376444 4140
rect 377956 4088 378008 4140
rect 393044 4088 393096 4140
rect 395988 4088 396040 4140
rect 414480 4088 414532 4140
rect 420828 4088 420880 4140
rect 443000 4088 443052 4140
rect 449808 4088 449860 4140
rect 477500 4088 477552 4140
rect 480168 4088 480220 4140
rect 83832 4020 83884 4072
rect 110512 4020 110564 4072
rect 295156 4020 295208 4072
rect 296720 4020 296772 4072
rect 340788 4020 340840 4072
rect 350264 4020 350316 4072
rect 351828 4020 351880 4072
rect 363328 4020 363380 4072
rect 367008 4020 367060 4072
rect 381176 4020 381228 4072
rect 382188 4020 382240 4072
rect 399024 4020 399076 4072
rect 401416 4020 401468 4072
rect 420368 4020 420420 4072
rect 423588 4020 423640 4072
rect 446588 4020 446640 4072
rect 447048 4020 447100 4072
rect 473912 4020 473964 4072
rect 474648 4020 474700 4072
rect 506020 4020 506072 4072
rect 20720 3952 20772 4004
rect 47584 3952 47636 4004
rect 64696 3952 64748 4004
rect 68284 3952 68336 4004
rect 19524 3884 19576 3936
rect 40684 3884 40736 3936
rect 46940 3884 46992 3936
rect 76656 3952 76708 4004
rect 98092 3952 98144 4004
rect 122840 3952 122892 4004
rect 332508 3952 332560 4004
rect 340696 3952 340748 4004
rect 342076 3952 342128 4004
rect 351368 3952 351420 4004
rect 354588 3952 354640 4004
rect 365720 3952 365772 4004
rect 373908 3952 373960 4004
rect 388260 3952 388312 4004
rect 390468 3952 390520 4004
rect 408500 3952 408552 4004
rect 411168 3952 411220 4004
rect 432328 3952 432380 4004
rect 438768 3952 438820 4004
rect 464436 3952 464488 4004
rect 464988 3952 465040 4004
rect 469496 3952 469548 4004
rect 471888 3952 471940 4004
rect 502432 3952 502484 4004
rect 75184 3884 75236 3936
rect 83004 3884 83056 3936
rect 84844 3884 84896 3936
rect 86960 3884 87012 3936
rect 87328 3884 87380 3936
rect 113364 3884 113416 3936
rect 325608 3884 325660 3936
rect 332416 3884 332468 3936
rect 335268 3884 335320 3936
rect 344284 3884 344336 3936
rect 347688 3884 347740 3936
rect 358544 3884 358596 3936
rect 360108 3884 360160 3936
rect 372804 3884 372856 3936
rect 378048 3884 378100 3936
rect 394240 3884 394292 3936
rect 397276 3884 397328 3936
rect 415676 3884 415728 3936
rect 419448 3884 419500 3936
rect 441804 3884 441856 3936
rect 444196 3884 444248 3936
rect 471520 3884 471572 3936
rect 477408 3884 477460 3936
rect 507308 3952 507360 4004
rect 508504 4088 508556 4140
rect 510804 4088 510856 4140
rect 514668 4088 514720 4140
rect 552388 4088 552440 4140
rect 507768 4020 507820 4072
rect 516876 4020 516928 4072
rect 516968 4020 517020 4072
rect 521476 4020 521528 4072
rect 528468 4020 528520 4072
rect 545304 4020 545356 4072
rect 547144 4020 547196 4072
rect 575020 4020 575072 4072
rect 510528 3952 510580 4004
rect 514852 3952 514904 4004
rect 528376 3952 528428 4004
rect 543004 3952 543056 4004
rect 548524 3952 548576 4004
rect 582196 3952 582248 4004
rect 513196 3884 513248 3936
rect 518808 3884 518860 3936
rect 557172 3884 557224 3936
rect 36176 3816 36228 3868
rect 64144 3816 64196 3868
rect 72976 3816 73028 3868
rect 102140 3816 102192 3868
rect 313188 3816 313240 3868
rect 318064 3816 318116 3868
rect 333888 3816 333940 3868
rect 341892 3816 341944 3868
rect 342168 3816 342220 3868
rect 352564 3816 352616 3868
rect 353208 3816 353260 3868
rect 364524 3816 364576 3868
rect 365536 3816 365588 3868
rect 378784 3816 378836 3868
rect 379428 3816 379480 3868
rect 395436 3816 395488 3868
rect 397368 3816 397420 3868
rect 416872 3816 416924 3868
rect 424968 3816 425020 3868
rect 448980 3816 449032 3868
rect 459468 3816 459520 3868
rect 489368 3816 489420 3868
rect 489828 3816 489880 3868
rect 523868 3816 523920 3868
rect 524328 3816 524380 3868
rect 564348 3816 564400 3868
rect 29092 3748 29144 3800
rect 60004 3748 60056 3800
rect 62396 3748 62448 3800
rect 92480 3748 92532 3800
rect 101588 3748 101640 3800
rect 125784 3748 125836 3800
rect 328368 3748 328420 3800
rect 335912 3748 335964 3800
rect 336648 3748 336700 3800
rect 345480 3748 345532 3800
rect 346308 3748 346360 3800
rect 356152 3748 356204 3800
rect 357256 3748 357308 3800
rect 369216 3748 369268 3800
rect 371148 3748 371200 3800
rect 385868 3748 385920 3800
rect 387708 3748 387760 3800
rect 404912 3748 404964 3800
rect 408408 3748 408460 3800
rect 428740 3748 428792 3800
rect 431868 3748 431920 3800
rect 456064 3748 456116 3800
rect 456708 3748 456760 3800
rect 485780 3748 485832 3800
rect 487068 3748 487120 3800
rect 514484 3748 514536 3800
rect 521568 3748 521620 3800
rect 560760 3748 560812 3800
rect 11244 3680 11296 3732
rect 43444 3680 43496 3732
rect 44548 3680 44600 3732
rect 47400 3680 47452 3732
rect 58808 3680 58860 3732
rect 89812 3680 89864 3732
rect 90916 3680 90968 3732
rect 5264 3612 5316 3664
rect 42984 3612 43036 3664
rect 51632 3612 51684 3664
rect 75184 3612 75236 3664
rect 81440 3612 81492 3664
rect 82636 3612 82688 3664
rect 2872 3544 2924 3596
rect 41420 3544 41472 3596
rect 54024 3544 54076 3596
rect 55128 3544 55180 3596
rect 60004 3544 60056 3596
rect 60648 3544 60700 3596
rect 61200 3544 61252 3596
rect 62028 3544 62080 3596
rect 62120 3544 62172 3596
rect 84844 3544 84896 3596
rect 84936 3544 84988 3596
rect 85488 3544 85540 3596
rect 86132 3544 86184 3596
rect 86868 3544 86920 3596
rect 88524 3544 88576 3596
rect 89628 3544 89680 3596
rect 89720 3544 89772 3596
rect 91008 3544 91060 3596
rect 94504 3680 94556 3732
rect 120080 3680 120132 3732
rect 106372 3612 106424 3664
rect 107568 3612 107620 3664
rect 117412 3544 117464 3596
rect 119436 3544 119488 3596
rect 119988 3544 120040 3596
rect 120632 3544 120684 3596
rect 121368 3544 121420 3596
rect 121828 3544 121880 3596
rect 122748 3544 122800 3596
rect 1676 3476 1728 3528
rect 40132 3476 40184 3528
rect 45744 3476 45796 3528
rect 46848 3476 46900 3528
rect 572 3408 624 3460
rect 40224 3408 40276 3460
rect 43352 3408 43404 3460
rect 75092 3476 75144 3528
rect 52828 3408 52880 3460
rect 53748 3408 53800 3460
rect 8852 3340 8904 3392
rect 9588 3340 9640 3392
rect 10048 3340 10100 3392
rect 10968 3340 11020 3392
rect 16028 3340 16080 3392
rect 16488 3340 16540 3392
rect 24308 3340 24360 3392
rect 24768 3340 24820 3392
rect 25504 3340 25556 3392
rect 26148 3340 26200 3392
rect 27896 3340 27948 3392
rect 28908 3340 28960 3392
rect 34980 3340 35032 3392
rect 35808 3340 35860 3392
rect 48136 3340 48188 3392
rect 55220 3340 55272 3392
rect 62120 3340 62172 3392
rect 63592 3340 63644 3392
rect 64788 3340 64840 3392
rect 68284 3340 68336 3392
rect 68928 3340 68980 3392
rect 70676 3408 70728 3460
rect 71688 3408 71740 3460
rect 76656 3408 76708 3460
rect 80244 3408 80296 3460
rect 103980 3476 104032 3528
rect 104808 3476 104860 3528
rect 114744 3476 114796 3528
rect 115848 3476 115900 3528
rect 129740 3680 129792 3732
rect 306288 3680 306340 3732
rect 309784 3680 309836 3732
rect 337936 3680 337988 3732
rect 346676 3680 346728 3732
rect 350356 3680 350408 3732
rect 360936 3680 360988 3732
rect 361396 3680 361448 3732
rect 375196 3680 375248 3732
rect 375288 3680 375340 3732
rect 390652 3680 390704 3732
rect 394608 3680 394660 3732
rect 413284 3680 413336 3732
rect 413928 3680 413980 3732
rect 435824 3680 435876 3732
rect 441528 3680 441580 3732
rect 467840 3680 467892 3732
rect 469128 3680 469180 3732
rect 500132 3680 500184 3732
rect 505008 3680 505060 3732
rect 541716 3680 541768 3732
rect 543004 3680 543056 3732
rect 548892 3680 548944 3732
rect 552664 3680 552716 3732
rect 581000 3680 581052 3732
rect 126612 3612 126664 3664
rect 147680 3612 147732 3664
rect 314476 3612 314528 3664
rect 319260 3612 319312 3664
rect 322848 3612 322900 3664
rect 328828 3612 328880 3664
rect 331128 3612 331180 3664
rect 338304 3612 338356 3664
rect 343548 3612 343600 3664
rect 353760 3612 353812 3664
rect 354496 3612 354548 3664
rect 366916 3612 366968 3664
rect 368388 3612 368440 3664
rect 382372 3612 382424 3664
rect 383568 3612 383620 3664
rect 400220 3612 400272 3664
rect 401508 3612 401560 3664
rect 421564 3612 421616 3664
rect 429108 3612 429160 3664
rect 453672 3612 453724 3664
rect 453948 3612 454000 3664
rect 482284 3612 482336 3664
rect 482928 3612 482980 3664
rect 516784 3612 516836 3664
rect 519452 3612 519504 3664
rect 520372 3612 520424 3664
rect 522948 3612 523000 3664
rect 563152 3612 563204 3664
rect 567844 3612 567896 3664
rect 579804 3612 579856 3664
rect 127808 3544 127860 3596
rect 149060 3544 149112 3596
rect 158720 3544 158772 3596
rect 159916 3544 159968 3596
rect 167092 3544 167144 3596
rect 168196 3544 168248 3596
rect 201500 3544 201552 3596
rect 202696 3544 202748 3596
rect 227720 3544 227772 3596
rect 228916 3544 228968 3596
rect 244372 3544 244424 3596
rect 245568 3544 245620 3596
rect 252652 3544 252704 3596
rect 253848 3544 253900 3596
rect 278872 3544 278924 3596
rect 280068 3544 280120 3596
rect 293868 3544 293920 3596
rect 295524 3544 295576 3596
rect 303436 3544 303488 3596
rect 307392 3544 307444 3596
rect 314568 3544 314620 3596
rect 320456 3544 320508 3596
rect 324228 3544 324280 3596
rect 331220 3544 331272 3596
rect 333796 3544 333848 3596
rect 343088 3544 343140 3596
rect 344928 3544 344980 3596
rect 354956 3544 355008 3596
rect 357256 3544 357308 3596
rect 370412 3544 370464 3596
rect 372528 3544 372580 3596
rect 387064 3544 387116 3596
rect 388996 3544 389048 3596
rect 407304 3544 407356 3596
rect 409788 3544 409840 3596
rect 431132 3544 431184 3596
rect 431776 3544 431828 3596
rect 457260 3544 457312 3596
rect 467748 3544 467800 3596
rect 93308 3340 93360 3392
rect 93768 3340 93820 3392
rect 95700 3340 95752 3392
rect 96528 3340 96580 3392
rect 96896 3340 96948 3392
rect 97908 3340 97960 3392
rect 102784 3340 102836 3392
rect 103428 3340 103480 3392
rect 104900 3408 104952 3460
rect 107660 3408 107712 3460
rect 105176 3340 105228 3392
rect 123024 3476 123076 3528
rect 124128 3476 124180 3528
rect 129004 3476 129056 3528
rect 129648 3476 129700 3528
rect 130200 3476 130252 3528
rect 80060 3272 80112 3324
rect 108764 3272 108816 3324
rect 131396 3340 131448 3392
rect 132408 3340 132460 3392
rect 124220 3272 124272 3324
rect 125508 3272 125560 3324
rect 132592 3408 132644 3460
rect 133696 3408 133748 3460
rect 136088 3408 136140 3460
rect 136548 3408 136600 3460
rect 137284 3408 137336 3460
rect 137928 3408 137980 3460
rect 138480 3408 138532 3460
rect 139308 3408 139360 3460
rect 139676 3408 139728 3460
rect 140688 3408 140740 3460
rect 145656 3476 145708 3528
rect 146208 3476 146260 3528
rect 146852 3476 146904 3528
rect 147588 3476 147640 3528
rect 148048 3476 148100 3528
rect 148968 3476 149020 3528
rect 150440 3476 150492 3528
rect 151728 3476 151780 3528
rect 153936 3476 153988 3528
rect 154488 3476 154540 3528
rect 155132 3476 155184 3528
rect 155868 3476 155920 3528
rect 156328 3476 156380 3528
rect 157248 3476 157300 3528
rect 162308 3476 162360 3528
rect 162768 3476 162820 3528
rect 163504 3476 163556 3528
rect 164148 3476 164200 3528
rect 165896 3476 165948 3528
rect 166908 3476 166960 3528
rect 171784 3476 171836 3528
rect 172428 3476 172480 3528
rect 172980 3476 173032 3528
rect 173808 3476 173860 3528
rect 180156 3476 180208 3528
rect 180708 3476 180760 3528
rect 182548 3476 182600 3528
rect 183468 3476 183520 3528
rect 183744 3476 183796 3528
rect 184756 3476 184808 3528
rect 188436 3476 188488 3528
rect 188988 3476 189040 3528
rect 189632 3476 189684 3528
rect 190368 3476 190420 3528
rect 192024 3476 192076 3528
rect 193128 3476 193180 3528
rect 193220 3476 193272 3528
rect 194508 3476 194560 3528
rect 196808 3476 196860 3528
rect 197268 3476 197320 3528
rect 198004 3476 198056 3528
rect 198648 3476 198700 3528
rect 199200 3476 199252 3528
rect 200028 3476 200080 3528
rect 200396 3476 200448 3528
rect 201408 3476 201460 3528
rect 205088 3476 205140 3528
rect 205548 3476 205600 3528
rect 207480 3476 207532 3528
rect 208308 3476 208360 3528
rect 208676 3476 208728 3528
rect 209688 3476 209740 3528
rect 209872 3476 209924 3528
rect 211068 3476 211120 3528
rect 214656 3476 214708 3528
rect 215208 3476 215260 3528
rect 215852 3476 215904 3528
rect 216588 3476 216640 3528
rect 217048 3476 217100 3528
rect 217968 3476 218020 3528
rect 218152 3476 218204 3528
rect 219256 3476 219308 3528
rect 222936 3476 222988 3528
rect 223488 3476 223540 3528
rect 224132 3476 224184 3528
rect 224868 3476 224920 3528
rect 225328 3476 225380 3528
rect 226248 3476 226300 3528
rect 226524 3476 226576 3528
rect 227628 3476 227680 3528
rect 231308 3476 231360 3528
rect 231768 3476 231820 3528
rect 232504 3476 232556 3528
rect 233148 3476 233200 3528
rect 233700 3476 233752 3528
rect 234528 3476 234580 3528
rect 239588 3476 239640 3528
rect 240048 3476 240100 3528
rect 240784 3476 240836 3528
rect 241428 3476 241480 3528
rect 243176 3476 243228 3528
rect 244188 3476 244240 3528
rect 249156 3476 249208 3528
rect 249708 3476 249760 3528
rect 251456 3476 251508 3528
rect 252468 3476 252520 3528
rect 257436 3476 257488 3528
rect 257988 3476 258040 3528
rect 258632 3476 258684 3528
rect 259368 3476 259420 3528
rect 262220 3476 262272 3528
rect 263692 3476 263744 3528
rect 265808 3476 265860 3528
rect 266268 3476 266320 3528
rect 268108 3476 268160 3528
rect 269028 3476 269080 3528
rect 269304 3476 269356 3528
rect 270408 3476 270460 3528
rect 272892 3476 272944 3528
rect 273352 3476 273404 3528
rect 276020 3476 276072 3528
rect 276480 3476 276532 3528
rect 281540 3476 281592 3528
rect 282460 3476 282512 3528
rect 291108 3476 291160 3528
rect 291936 3476 291988 3528
rect 292488 3476 292540 3528
rect 294328 3476 294380 3528
rect 298008 3476 298060 3528
rect 300308 3476 300360 3528
rect 302148 3476 302200 3528
rect 305000 3476 305052 3528
rect 309048 3476 309100 3528
rect 313372 3476 313424 3528
rect 317328 3476 317380 3528
rect 322848 3476 322900 3528
rect 331036 3476 331088 3528
rect 339500 3476 339552 3528
rect 346216 3476 346268 3528
rect 357348 3476 357400 3528
rect 358728 3476 358780 3528
rect 371608 3476 371660 3528
rect 373816 3476 373868 3528
rect 389456 3476 389508 3528
rect 393136 3476 393188 3528
rect 412088 3476 412140 3528
rect 416596 3476 416648 3528
rect 439412 3476 439464 3528
rect 440148 3476 440200 3528
rect 466828 3476 466880 3528
rect 467932 3476 467984 3528
rect 469128 3476 469180 3528
rect 469312 3544 469364 3596
rect 492956 3544 493008 3596
rect 495348 3544 495400 3596
rect 531044 3544 531096 3596
rect 532608 3544 532660 3596
rect 573824 3544 573876 3596
rect 498936 3476 498988 3528
rect 499396 3476 499448 3528
rect 535736 3476 535788 3528
rect 536748 3476 536800 3528
rect 578608 3476 578660 3528
rect 164700 3408 164752 3460
rect 165528 3408 165580 3460
rect 241980 3408 242032 3460
rect 242808 3408 242860 3460
rect 250352 3408 250404 3460
rect 251088 3408 251140 3460
rect 295248 3408 295300 3460
rect 297916 3408 297968 3460
rect 300768 3408 300820 3460
rect 303804 3408 303856 3460
rect 306196 3408 306248 3460
rect 310980 3408 311032 3460
rect 315948 3408 316000 3460
rect 321652 3408 321704 3460
rect 322756 3408 322808 3460
rect 330024 3408 330076 3460
rect 338028 3408 338080 3460
rect 347872 3408 347924 3460
rect 350448 3408 350500 3460
rect 362132 3408 362184 3460
rect 365628 3408 365680 3460
rect 379980 3408 380032 3460
rect 380716 3408 380768 3460
rect 397828 3408 397880 3460
rect 404176 3408 404228 3460
rect 425060 3408 425112 3460
rect 425152 3408 425204 3460
rect 426348 3408 426400 3460
rect 426440 3408 426492 3460
rect 450176 3408 450228 3460
rect 455328 3408 455380 3460
rect 484584 3408 484636 3460
rect 492588 3408 492640 3460
rect 527456 3408 527508 3460
rect 529664 3408 529716 3460
rect 571432 3408 571484 3460
rect 150624 3340 150676 3392
rect 170588 3340 170640 3392
rect 171048 3340 171100 3392
rect 247960 3340 248012 3392
rect 249064 3340 249116 3392
rect 310336 3340 310388 3392
rect 315764 3340 315816 3392
rect 318616 3340 318668 3392
rect 325240 3340 325292 3392
rect 326896 3340 326948 3392
rect 333612 3340 333664 3392
rect 355968 3340 356020 3392
rect 368020 3340 368072 3392
rect 369768 3340 369820 3392
rect 384672 3340 384724 3392
rect 391848 3340 391900 3392
rect 409696 3340 409748 3392
rect 412548 3340 412600 3392
rect 422300 3340 422352 3392
rect 434720 3340 434772 3392
rect 459652 3340 459704 3392
rect 463608 3340 463660 3392
rect 469312 3340 469364 3392
rect 469404 3340 469456 3392
rect 491760 3340 491812 3392
rect 496084 3340 496136 3392
rect 507216 3340 507268 3392
rect 507308 3340 507360 3392
rect 509608 3340 509660 3392
rect 511908 3340 511960 3392
rect 550088 3340 550140 3392
rect 132684 3272 132736 3324
rect 149244 3272 149296 3324
rect 150348 3272 150400 3324
rect 157524 3272 157576 3324
rect 158628 3272 158680 3324
rect 174176 3272 174228 3324
rect 175188 3272 175240 3324
rect 234804 3272 234856 3324
rect 235908 3272 235960 3324
rect 280160 3272 280212 3324
rect 281264 3272 281316 3324
rect 310428 3272 310480 3324
rect 314568 3272 314620 3324
rect 369676 3272 369728 3324
rect 383568 3272 383620 3324
rect 389088 3272 389140 3324
rect 406108 3272 406160 3324
rect 407028 3272 407080 3324
rect 427544 3272 427596 3324
rect 236000 3204 236052 3256
rect 237288 3204 237340 3256
rect 267004 3204 267056 3256
rect 267832 3204 267884 3256
rect 274824 3204 274876 3256
rect 275284 3204 275336 3256
rect 307668 3204 307720 3256
rect 312176 3204 312228 3256
rect 364248 3204 364300 3256
rect 377588 3204 377640 3256
rect 386328 3204 386380 3256
rect 403716 3204 403768 3256
rect 404268 3204 404320 3256
rect 423956 3204 424008 3256
rect 303528 3136 303580 3188
rect 306196 3136 306248 3188
rect 361488 3136 361540 3188
rect 374000 3136 374052 3188
rect 380808 3136 380860 3188
rect 396632 3136 396684 3188
rect 398748 3136 398800 3188
rect 417976 3136 418028 3188
rect 422300 3136 422352 3188
rect 434628 3272 434680 3324
rect 437388 3272 437440 3324
rect 463240 3272 463292 3324
rect 466368 3272 466420 3324
rect 496544 3272 496596 3324
rect 502248 3272 502300 3324
rect 538128 3272 538180 3324
rect 544384 3272 544436 3324
rect 546500 3272 546552 3324
rect 546592 3272 546644 3324
rect 577412 3272 577464 3324
rect 427728 3204 427780 3256
rect 452476 3204 452528 3256
rect 452568 3204 452620 3256
rect 481088 3204 481140 3256
rect 481548 3204 481600 3256
rect 514392 3204 514444 3256
rect 514484 3204 514536 3256
rect 520280 3204 520332 3256
rect 520372 3204 520424 3256
rect 555976 3204 556028 3256
rect 436008 3136 436060 3188
rect 460848 3136 460900 3188
rect 462228 3136 462280 3188
rect 469404 3136 469456 3188
rect 469496 3136 469548 3188
rect 495348 3136 495400 3188
rect 499488 3136 499540 3188
rect 534540 3136 534592 3188
rect 537484 3136 537536 3188
rect 570236 3136 570288 3188
rect 181352 3068 181404 3120
rect 182088 3068 182140 3120
rect 376668 3068 376720 3120
rect 391848 3068 391900 3120
rect 393228 3068 393280 3120
rect 410892 3068 410944 3120
rect 422208 3068 422260 3120
rect 445392 3068 445444 3120
rect 459376 3068 459428 3120
rect 488172 3068 488224 3120
rect 493968 3068 494020 3120
rect 528652 3068 528704 3120
rect 534724 3068 534776 3120
rect 566740 3068 566792 3120
rect 18328 3000 18380 3052
rect 19248 3000 19300 3052
rect 140872 3000 140924 3052
rect 142068 3000 142120 3052
rect 175372 3000 175424 3052
rect 176476 3000 176528 3052
rect 190828 3000 190880 3052
rect 191748 3000 191800 3052
rect 206284 3000 206336 3052
rect 206928 3000 206980 3052
rect 259828 3000 259880 3052
rect 260748 3000 260800 3052
rect 261024 3000 261076 3052
rect 262128 3000 262180 3052
rect 299388 3000 299440 3052
rect 301412 3000 301464 3052
rect 311808 3000 311860 3052
rect 316960 3000 317012 3052
rect 321468 3000 321520 3052
rect 327632 3000 327684 3052
rect 384948 3000 385000 3052
rect 402520 3000 402572 3052
rect 416688 3000 416740 3052
rect 438216 3000 438268 3052
rect 452292 3000 452344 3052
rect 479892 3000 479944 3052
rect 483664 3000 483716 3052
rect 503628 3000 503680 3052
rect 512644 3000 512696 3052
rect 517888 3000 517940 3052
rect 521108 3000 521160 3052
rect 525064 3000 525116 3052
rect 526444 3000 526496 3052
rect 559564 3000 559616 3052
rect 291016 2932 291068 2984
rect 293132 2932 293184 2984
rect 299296 2932 299348 2984
rect 302608 2932 302660 2984
rect 329748 2932 329800 2984
rect 337108 2932 337160 2984
rect 384856 2932 384908 2984
rect 401324 2932 401376 2984
rect 451188 2932 451240 2984
rect 478696 2932 478748 2984
rect 516876 2932 516928 2984
rect 528468 2932 528520 2984
rect 540244 2932 540296 2984
rect 546592 2932 546644 2984
rect 274088 2864 274140 2916
rect 274548 2864 274600 2916
rect 318708 2864 318760 2916
rect 324044 2864 324096 2916
rect 326988 2864 327040 2916
rect 334716 2864 334768 2916
rect 448428 2864 448480 2916
rect 475108 2864 475160 2916
rect 514852 2864 514904 2916
rect 528376 2864 528428 2916
rect 529204 2864 529256 2916
rect 532240 2864 532292 2916
rect 541624 2864 541676 2916
rect 552664 2932 552716 2984
rect 547236 2864 547288 2916
rect 567844 2932 567896 2984
rect 118240 2796 118292 2848
rect 118608 2796 118660 2848
rect 444288 2796 444340 2848
rect 470324 2796 470376 2848
rect 545764 2796 545816 2848
rect 553584 2796 553636 2848
rect 109960 552 110012 604
rect 110328 552 110380 604
rect 418252 552 418304 604
rect 419172 552 419224 604
rect 429200 552 429252 604
rect 429936 552 429988 604
rect 436192 552 436244 604
rect 437020 552 437072 604
rect 447140 552 447192 604
rect 447784 552 447836 604
rect 454224 552 454276 604
rect 454868 552 454920 604
rect 461032 552 461084 604
rect 462044 552 462096 604
rect 472072 552 472124 604
rect 472716 552 472768 604
rect 485872 552 485924 604
rect 486976 552 487028 604
rect 489920 552 489972 604
rect 490564 552 490616 604
rect 496820 552 496872 604
rect 497740 552 497792 604
rect 525800 552 525852 604
rect 526260 552 526312 604
rect 538312 552 538364 604
rect 539324 552 539376 604
rect 542360 552 542412 604
rect 542912 552 542964 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 40512 700466 40540 703520
rect 72988 700670 73016 703520
rect 89180 700738 89208 703520
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 72976 700664 73028 700670
rect 72976 700606 73028 700612
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 105464 699718 105492 703520
rect 137848 700942 137876 703520
rect 154132 701010 154160 703520
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 137836 700936 137888 700942
rect 137836 700878 137888 700884
rect 170324 699718 170352 703520
rect 202800 700126 202828 703520
rect 202788 700120 202840 700126
rect 202788 700062 202840 700068
rect 218992 700058 219020 703520
rect 218980 700052 219032 700058
rect 218980 699994 219032 700000
rect 235184 699718 235212 703520
rect 256608 700868 256660 700874
rect 256608 700810 256660 700816
rect 244188 700596 244240 700602
rect 244188 700538 244240 700544
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 106200 688090 106228 699654
rect 171060 688226 171088 699654
rect 230388 696992 230440 696998
rect 230388 696934 230440 696940
rect 230400 690742 230428 696934
rect 229100 690736 229152 690742
rect 229100 690678 229152 690684
rect 230388 690736 230440 690742
rect 230388 690678 230440 690684
rect 171048 688220 171100 688226
rect 171048 688162 171100 688168
rect 106188 688084 106240 688090
rect 106188 688026 106240 688032
rect 229008 687268 229060 687274
rect 229008 687210 229060 687216
rect 124220 687200 124272 687206
rect 4802 687168 4858 687177
rect 124220 687142 124272 687148
rect 4802 687103 4858 687112
rect 111800 687132 111852 687138
rect 3698 686896 3754 686905
rect 3698 686831 3754 686840
rect 2872 686724 2924 686730
rect 2872 686666 2924 686672
rect 2780 682304 2832 682310
rect 2778 682272 2780 682281
rect 2832 682272 2834 682281
rect 2778 682207 2834 682216
rect 2780 669316 2832 669322
rect 2780 669258 2832 669264
rect 2792 668001 2820 669258
rect 2778 667992 2834 668001
rect 2778 667927 2834 667936
rect 2780 654084 2832 654090
rect 2780 654026 2832 654032
rect 2792 653585 2820 654026
rect 2778 653576 2834 653585
rect 2778 653511 2834 653520
rect 2780 624912 2832 624918
rect 2778 624880 2780 624889
rect 2832 624880 2834 624889
rect 2778 624815 2834 624824
rect 2780 610496 2832 610502
rect 2778 610464 2780 610473
rect 2832 610464 2834 610473
rect 2778 610399 2834 610408
rect 2780 596148 2832 596154
rect 2780 596090 2832 596096
rect 2792 596057 2820 596090
rect 2778 596048 2834 596057
rect 2778 595983 2834 595992
rect 2780 567384 2832 567390
rect 2778 567352 2780 567361
rect 2832 567352 2834 567361
rect 2778 567287 2834 567296
rect 2780 553376 2832 553382
rect 2780 553318 2832 553324
rect 2792 553081 2820 553318
rect 2778 553072 2834 553081
rect 2778 553007 2834 553016
rect 2780 539572 2832 539578
rect 2780 539514 2832 539520
rect 2792 538665 2820 539514
rect 2778 538656 2834 538665
rect 2778 538591 2834 538600
rect 2780 509992 2832 509998
rect 2778 509960 2780 509969
rect 2832 509960 2834 509969
rect 2778 509895 2834 509904
rect 2884 495553 2912 686666
rect 3056 686316 3108 686322
rect 3056 686258 3108 686264
rect 2964 683528 3016 683534
rect 2964 683470 3016 683476
rect 2870 495544 2926 495553
rect 2870 495479 2926 495488
rect 2872 481636 2924 481642
rect 2872 481578 2924 481584
rect 2884 481137 2912 481578
rect 2870 481128 2926 481137
rect 2870 481063 2926 481072
rect 2872 452464 2924 452470
rect 2870 452432 2872 452441
rect 2924 452432 2926 452441
rect 2870 452367 2926 452376
rect 2780 438728 2832 438734
rect 2780 438670 2832 438676
rect 2792 438025 2820 438670
rect 2778 438016 2834 438025
rect 2778 437951 2834 437960
rect 2872 425060 2924 425066
rect 2872 425002 2924 425008
rect 2884 423745 2912 425002
rect 2870 423736 2926 423745
rect 2870 423671 2926 423680
rect 2872 395072 2924 395078
rect 2870 395040 2872 395049
rect 2924 395040 2926 395049
rect 2870 394975 2926 394984
rect 2976 380633 3004 683470
rect 2962 380624 3018 380633
rect 2962 380559 3018 380568
rect 2964 367056 3016 367062
rect 2964 366998 3016 367004
rect 2976 366217 3004 366998
rect 2962 366208 3018 366217
rect 2962 366143 3018 366152
rect 2964 337612 3016 337618
rect 2964 337554 3016 337560
rect 2976 337521 3004 337554
rect 2962 337512 3018 337521
rect 2962 337447 3018 337456
rect 2964 323128 3016 323134
rect 2962 323096 2964 323105
rect 3016 323096 3018 323105
rect 2962 323031 3018 323040
rect 3068 308825 3096 686258
rect 3514 686216 3570 686225
rect 3240 686180 3292 686186
rect 3514 686151 3570 686160
rect 3240 686122 3292 686128
rect 3148 683392 3200 683398
rect 3148 683334 3200 683340
rect 3054 308816 3110 308825
rect 3054 308751 3110 308760
rect 3056 295316 3108 295322
rect 3056 295258 3108 295264
rect 3068 294409 3096 295258
rect 3054 294400 3110 294409
rect 3054 294335 3110 294344
rect 3160 280129 3188 683334
rect 3146 280120 3202 280129
rect 3146 280055 3202 280064
rect 3252 265713 3280 686122
rect 3332 686112 3384 686118
rect 3332 686054 3384 686060
rect 3238 265704 3294 265713
rect 3238 265639 3294 265648
rect 3148 251320 3200 251326
rect 3146 251288 3148 251297
rect 3200 251288 3202 251297
rect 3146 251223 3202 251232
rect 3344 237017 3372 686054
rect 3422 683768 3478 683777
rect 3422 683703 3478 683712
rect 3330 237008 3386 237017
rect 3330 236943 3386 236952
rect 3332 223576 3384 223582
rect 3332 223518 3384 223524
rect 3344 222601 3372 223518
rect 3330 222592 3386 222601
rect 3330 222527 3386 222536
rect 2780 208208 2832 208214
rect 2778 208176 2780 208185
rect 2832 208176 2834 208185
rect 2778 208111 2834 208120
rect 2780 179512 2832 179518
rect 2778 179480 2780 179489
rect 2832 179480 2834 179489
rect 2778 179415 2834 179424
rect 3148 165572 3200 165578
rect 3148 165514 3200 165520
rect 3160 165073 3188 165514
rect 3146 165064 3202 165073
rect 3146 164999 3202 165008
rect 3332 136604 3384 136610
rect 3332 136546 3384 136552
rect 3344 136377 3372 136546
rect 3330 136368 3386 136377
rect 3330 136303 3386 136312
rect 3332 122800 3384 122806
rect 3332 122742 3384 122748
rect 3344 122097 3372 122742
rect 3330 122088 3386 122097
rect 3330 122023 3386 122032
rect 3332 80028 3384 80034
rect 3332 79970 3384 79976
rect 3344 78985 3372 79970
rect 3330 78976 3386 78985
rect 3330 78911 3386 78920
rect 3436 7177 3464 683703
rect 3528 35873 3556 686151
rect 3606 683496 3662 683505
rect 3606 683431 3662 683440
rect 3620 50153 3648 683431
rect 3712 93265 3740 686831
rect 3882 686624 3938 686633
rect 3882 686559 3938 686568
rect 3790 683360 3846 683369
rect 3790 683295 3846 683304
rect 3698 93256 3754 93265
rect 3698 93191 3754 93200
rect 3804 64569 3832 683295
rect 3896 107681 3924 686559
rect 4068 685976 4120 685982
rect 4068 685918 4120 685924
rect 3974 683632 4030 683641
rect 3974 683567 4030 683576
rect 3988 150793 4016 683567
rect 4080 193905 4108 685918
rect 4066 193896 4122 193905
rect 4066 193831 4122 193840
rect 4816 179518 4844 687103
rect 111800 687074 111852 687080
rect 84198 687032 84254 687041
rect 63868 686996 63920 687002
rect 84198 686967 84254 686976
rect 63868 686938 63920 686944
rect 4988 686588 5040 686594
rect 4988 686530 5040 686536
rect 4896 683324 4948 683330
rect 4896 683266 4948 683272
rect 4908 208214 4936 683266
rect 5000 438734 5028 686530
rect 7564 686384 7616 686390
rect 7564 686326 7616 686332
rect 57978 686352 58034 686361
rect 5540 685636 5592 685642
rect 5540 685578 5592 685584
rect 5080 683868 5132 683874
rect 5080 683810 5132 683816
rect 5092 610502 5120 683810
rect 5552 682310 5580 685578
rect 6736 685432 6788 685438
rect 6736 685374 6788 685380
rect 6644 685228 6696 685234
rect 6644 685170 6696 685176
rect 6182 685128 6238 685137
rect 6182 685063 6238 685072
rect 5540 682304 5592 682310
rect 5540 682246 5592 682252
rect 5080 610496 5132 610502
rect 5080 610438 5132 610444
rect 4988 438728 5040 438734
rect 4988 438670 5040 438676
rect 6196 251326 6224 685063
rect 6552 685024 6604 685030
rect 6552 684966 6604 684972
rect 6460 684820 6512 684826
rect 6460 684762 6512 684768
rect 6368 684752 6420 684758
rect 6368 684694 6420 684700
rect 6276 684548 6328 684554
rect 6276 684490 6328 684496
rect 6288 337618 6316 684490
rect 6380 395078 6408 684694
rect 6472 452470 6500 684762
rect 6564 509998 6592 684966
rect 6656 567390 6684 685170
rect 6748 624918 6776 685374
rect 6826 683768 6882 683777
rect 6826 683703 6882 683712
rect 6840 683233 6868 683703
rect 6826 683224 6882 683233
rect 6826 683159 6882 683168
rect 6736 624912 6788 624918
rect 6736 624854 6788 624860
rect 6644 567384 6696 567390
rect 6644 567326 6696 567332
rect 6552 509992 6604 509998
rect 6552 509934 6604 509940
rect 6460 452464 6512 452470
rect 6460 452406 6512 452412
rect 6368 395072 6420 395078
rect 6368 395014 6420 395020
rect 6276 337612 6328 337618
rect 6276 337554 6328 337560
rect 7576 323134 7604 686326
rect 57978 686287 58034 686296
rect 45558 686080 45614 686089
rect 45558 686015 45614 686024
rect 41418 685944 41474 685953
rect 39856 685908 39908 685914
rect 41418 685879 41474 685888
rect 39856 685850 39908 685856
rect 39394 685264 39450 685273
rect 39394 685199 39450 685208
rect 25596 685092 25648 685098
rect 25596 685034 25648 685040
rect 24122 684720 24178 684729
rect 24122 684655 24178 684664
rect 22742 683904 22798 683913
rect 22742 683839 22798 683848
rect 16578 683768 16634 683777
rect 16578 683703 16634 683712
rect 16592 683233 16620 683703
rect 16578 683224 16634 683233
rect 16578 683159 16634 683168
rect 7564 323128 7616 323134
rect 7564 323070 7616 323076
rect 6184 251320 6236 251326
rect 6184 251262 6236 251268
rect 4896 208208 4948 208214
rect 4896 208150 4948 208156
rect 4804 179512 4856 179518
rect 4804 179454 4856 179460
rect 3974 150784 4030 150793
rect 3974 150719 4030 150728
rect 22756 136610 22784 683839
rect 22744 136604 22796 136610
rect 22744 136546 22796 136552
rect 24136 122806 24164 684655
rect 25504 684616 25556 684622
rect 25504 684558 25556 684564
rect 25516 295322 25544 684558
rect 25608 425066 25636 685034
rect 38108 684412 38160 684418
rect 38108 684354 38160 684360
rect 33784 684344 33836 684350
rect 33784 684286 33836 684292
rect 32404 683800 32456 683806
rect 32404 683742 32456 683748
rect 29644 683460 29696 683466
rect 29644 683402 29696 683408
rect 25596 425060 25648 425066
rect 25596 425002 25648 425008
rect 25504 295316 25556 295322
rect 25504 295258 25556 295264
rect 29656 223582 29684 683402
rect 32416 367062 32444 683742
rect 33796 669322 33824 684286
rect 38016 684208 38068 684214
rect 38016 684150 38068 684156
rect 37924 683936 37976 683942
rect 37924 683878 37976 683884
rect 35806 683768 35862 683777
rect 35806 683703 35862 683712
rect 35820 683233 35848 683703
rect 35806 683224 35862 683233
rect 35806 683159 35862 683168
rect 33784 669316 33836 669322
rect 33784 669258 33836 669264
rect 37936 481642 37964 683878
rect 38028 596154 38056 684150
rect 38120 654090 38148 684354
rect 39302 683768 39358 683777
rect 39302 683703 39358 683712
rect 38108 654084 38160 654090
rect 38108 654026 38160 654032
rect 38016 596148 38068 596154
rect 38016 596090 38068 596096
rect 37924 481636 37976 481642
rect 37924 481578 37976 481584
rect 32404 367056 32456 367062
rect 32404 366998 32456 367004
rect 29644 223576 29696 223582
rect 29644 223518 29696 223524
rect 24124 122800 24176 122806
rect 24124 122742 24176 122748
rect 3882 107672 3938 107681
rect 3882 107607 3938 107616
rect 39316 80034 39344 683703
rect 39408 165578 39436 685199
rect 39488 684072 39540 684078
rect 39488 684014 39540 684020
rect 39500 539578 39528 684014
rect 39580 684004 39632 684010
rect 39580 683946 39632 683952
rect 39592 553382 39620 683946
rect 39580 553376 39632 553382
rect 39580 553318 39632 553324
rect 39488 539572 39540 539578
rect 39488 539514 39540 539520
rect 39396 165572 39448 165578
rect 39396 165514 39448 165520
rect 39304 80028 39356 80034
rect 39304 79970 39356 79976
rect 3790 64560 3846 64569
rect 3790 64495 3846 64504
rect 26148 62076 26200 62082
rect 26148 62018 26200 62024
rect 24768 62008 24820 62014
rect 24768 61950 24820 61956
rect 19248 61940 19300 61946
rect 19248 61882 19300 61888
rect 15108 61804 15160 61810
rect 15108 61746 15160 61752
rect 10968 61736 11020 61742
rect 10968 61678 11020 61684
rect 9588 61600 9640 61606
rect 9588 61542 9640 61548
rect 6828 61464 6880 61470
rect 6828 61406 6880 61412
rect 4068 61396 4120 61402
rect 4068 61338 4120 61344
rect 3606 50144 3662 50153
rect 3606 50079 3662 50088
rect 3514 35864 3570 35873
rect 3514 35799 3570 35808
rect 3516 22092 3568 22098
rect 3516 22034 3568 22040
rect 3528 21457 3556 22034
rect 3514 21448 3570 21457
rect 3514 21383 3570 21392
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3470
rect 2884 480 2912 3538
rect 4080 480 4108 61338
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5276 480 5304 3606
rect 6840 626 6868 61406
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 6472 598 6868 626
rect 6472 480 6500 598
rect 7668 480 7696 4762
rect 9600 3398 9628 61542
rect 10980 3398 11008 61678
rect 13636 61532 13688 61538
rect 13636 61474 13688 61480
rect 12440 4956 12492 4962
rect 12440 4898 12492 4904
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 8864 480 8892 3334
rect 10060 480 10088 3334
rect 11256 480 11284 3674
rect 12452 480 12480 4898
rect 13648 480 13676 61474
rect 15120 3482 15148 61746
rect 16488 61668 16540 61674
rect 16488 61610 16540 61616
rect 14844 3454 15148 3482
rect 14844 480 14872 3454
rect 16500 3398 16528 61610
rect 17224 4888 17276 4894
rect 17224 4830 17276 4836
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16040 480 16068 3334
rect 17236 480 17264 4830
rect 19260 3058 19288 61882
rect 23388 61872 23440 61878
rect 23388 61814 23440 61820
rect 21916 5024 21968 5030
rect 21916 4966 21968 4972
rect 20720 4004 20772 4010
rect 20720 3946 20772 3952
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 18340 480 18368 2994
rect 19536 480 19564 3878
rect 20732 480 20760 3946
rect 21928 480 21956 4966
rect 23400 3482 23428 61814
rect 23124 3454 23428 3482
rect 23124 480 23152 3454
rect 24780 3398 24808 61950
rect 26160 3398 26188 62018
rect 31668 61328 31720 61334
rect 31668 61270 31720 61276
rect 28908 61260 28960 61266
rect 28908 61202 28960 61208
rect 26700 5092 26752 5098
rect 26700 5034 26752 5040
rect 24308 3392 24360 3398
rect 24308 3334 24360 3340
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 25504 3392 25556 3398
rect 25504 3334 25556 3340
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 24320 480 24348 3334
rect 25516 480 25544 3334
rect 26712 480 26740 5034
rect 28920 3398 28948 61202
rect 30288 5160 30340 5166
rect 30288 5102 30340 5108
rect 29092 3800 29144 3806
rect 29092 3742 29144 3748
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 27908 480 27936 3334
rect 29104 480 29132 3742
rect 30300 480 30328 5102
rect 31680 3482 31708 61270
rect 33048 61192 33100 61198
rect 33048 61134 33100 61140
rect 33060 3482 33088 61134
rect 38476 61056 38528 61062
rect 38476 60998 38528 61004
rect 35808 60988 35860 60994
rect 35808 60930 35860 60936
rect 33876 5296 33928 5302
rect 33876 5238 33928 5244
rect 31496 3454 31708 3482
rect 32692 3454 33088 3482
rect 31496 480 31524 3454
rect 32692 480 32720 3454
rect 33888 480 33916 5238
rect 35820 3398 35848 60930
rect 37372 5364 37424 5370
rect 37372 5306 37424 5312
rect 36176 3868 36228 3874
rect 36176 3810 36228 3816
rect 34980 3392 35032 3398
rect 34980 3334 35032 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 34992 480 35020 3334
rect 36188 480 36216 3810
rect 37384 480 37412 5306
rect 38488 626 38516 60998
rect 39868 30326 39896 685850
rect 41432 683890 41460 685879
rect 45572 683890 45600 686015
rect 49700 685908 49752 685914
rect 49700 685850 49752 685856
rect 49712 684570 49740 685850
rect 55126 684584 55182 684593
rect 49712 684542 50016 684570
rect 49988 683890 50016 684542
rect 55126 684519 55182 684528
rect 55140 683890 55168 684519
rect 57992 684162 58020 686287
rect 57992 684134 58756 684162
rect 41432 683862 41676 683890
rect 45572 683862 46000 683890
rect 49988 683862 50416 683890
rect 54832 683862 55168 683890
rect 58728 683890 58756 684134
rect 63880 683890 63908 686938
rect 75918 686760 75974 686769
rect 75918 686695 75974 686704
rect 71778 686488 71834 686497
rect 71778 686423 71834 686432
rect 68282 684856 68338 684865
rect 68282 684791 68338 684800
rect 68296 683890 68324 684791
rect 58728 683862 59156 683890
rect 63572 683862 63908 683890
rect 67988 683862 68324 683890
rect 71792 683890 71820 686423
rect 75932 684570 75960 686695
rect 81346 684992 81402 685001
rect 81346 684927 81402 684936
rect 75932 684542 76328 684570
rect 76300 683890 76328 684542
rect 81360 683890 81388 684927
rect 84212 684570 84240 686967
rect 102140 686452 102192 686458
rect 102140 686394 102192 686400
rect 93860 685908 93912 685914
rect 93860 685850 93912 685856
rect 84212 684542 85068 684570
rect 71792 683862 72312 683890
rect 76300 683862 76728 683890
rect 81144 683862 81388 683890
rect 85040 683890 85068 684542
rect 93872 683890 93900 685850
rect 102152 684570 102180 686394
rect 106280 686044 106332 686050
rect 106280 685986 106332 685992
rect 102152 684542 102640 684570
rect 102612 683890 102640 684542
rect 106292 684162 106320 685986
rect 106292 684134 107056 684162
rect 107028 683890 107056 684134
rect 111812 683890 111840 687074
rect 115940 686520 115992 686526
rect 115940 686462 115992 686468
rect 85040 683862 85468 683890
rect 93872 683862 94300 683890
rect 102612 683862 103040 683890
rect 107028 683862 107456 683890
rect 111780 683862 111840 683890
rect 115952 683890 115980 686462
rect 120906 685400 120962 685409
rect 120906 685335 120962 685344
rect 120920 683890 120948 685335
rect 124232 684570 124260 687142
rect 150440 687064 150492 687070
rect 150440 687006 150492 687012
rect 128360 686656 128412 686662
rect 128360 686598 128412 686604
rect 128372 684570 128400 686598
rect 132500 686248 132552 686254
rect 132500 686190 132552 686196
rect 132512 684570 132540 686190
rect 147220 684956 147272 684962
rect 147220 684898 147272 684904
rect 124232 684542 124536 684570
rect 128372 684542 128952 684570
rect 132512 684542 133368 684570
rect 115952 683862 116196 683890
rect 120612 683862 120948 683890
rect 124508 683890 124536 684542
rect 128924 683890 128952 684542
rect 133340 683890 133368 684542
rect 147232 683890 147260 684898
rect 150452 684570 150480 687006
rect 229020 687002 229048 687210
rect 229112 687002 229140 690678
rect 235920 688362 235948 699654
rect 244200 690742 244228 700538
rect 248328 700528 248380 700534
rect 248328 700470 248380 700476
rect 248340 690742 248368 700470
rect 256620 690742 256648 700810
rect 262128 700800 262180 700806
rect 262128 700742 262180 700748
rect 262140 690742 262168 700742
rect 267660 699854 267688 703520
rect 274548 700256 274600 700262
rect 274548 700198 274600 700204
rect 270408 700188 270460 700194
rect 270408 700130 270460 700136
rect 267648 699848 267700 699854
rect 267648 699790 267700 699796
rect 270420 690742 270448 700130
rect 274560 690742 274588 700198
rect 283852 699786 283880 703520
rect 300136 703474 300164 703520
rect 300136 703446 300256 703474
rect 288348 699984 288400 699990
rect 288348 699926 288400 699932
rect 284208 699916 284260 699922
rect 284208 699858 284260 699864
rect 283840 699780 283892 699786
rect 283840 699722 283892 699728
rect 242900 690736 242952 690742
rect 242900 690678 242952 690684
rect 244188 690736 244240 690742
rect 244188 690678 244240 690684
rect 247040 690736 247092 690742
rect 247040 690678 247092 690684
rect 248328 690736 248380 690742
rect 248328 690678 248380 690684
rect 255320 690736 255372 690742
rect 255320 690678 255372 690684
rect 256608 690736 256660 690742
rect 256608 690678 256660 690684
rect 260840 690736 260892 690742
rect 260840 690678 260892 690684
rect 262128 690736 262180 690742
rect 262128 690678 262180 690684
rect 269120 690736 269172 690742
rect 269120 690678 269172 690684
rect 270408 690736 270460 690742
rect 270408 690678 270460 690684
rect 273260 690736 273312 690742
rect 273260 690678 273312 690684
rect 274548 690736 274600 690742
rect 274548 690678 274600 690684
rect 235908 688356 235960 688362
rect 235908 688298 235960 688304
rect 238760 687948 238812 687954
rect 238760 687890 238812 687896
rect 230020 687268 230072 687274
rect 230020 687210 230072 687216
rect 230032 687002 230060 687210
rect 229008 686996 229060 687002
rect 229008 686938 229060 686944
rect 229100 686996 229152 687002
rect 229100 686938 229152 686944
rect 229928 686996 229980 687002
rect 229928 686938 229980 686944
rect 230020 686996 230072 687002
rect 230020 686938 230072 686944
rect 233240 686996 233292 687002
rect 233240 686938 233292 686944
rect 234620 686996 234672 687002
rect 234620 686938 234672 686944
rect 168380 686928 168432 686934
rect 168380 686870 168432 686876
rect 164240 686860 164292 686866
rect 164240 686802 164292 686808
rect 154580 686792 154632 686798
rect 154580 686734 154632 686740
rect 150452 684542 150848 684570
rect 124508 683862 124936 683890
rect 128924 683862 129352 683890
rect 133340 683862 133768 683890
rect 146924 683862 147260 683890
rect 150820 683890 150848 684542
rect 154592 684026 154620 686734
rect 160376 684684 160428 684690
rect 160376 684626 160428 684632
rect 154592 683998 155264 684026
rect 155236 683890 155264 683998
rect 160388 683890 160416 684626
rect 150820 683862 151248 683890
rect 155236 683862 155664 683890
rect 160080 683862 160416 683890
rect 164252 683890 164280 686802
rect 168392 683890 168420 686870
rect 226156 685840 226208 685846
rect 226156 685782 226208 685788
rect 213000 685772 213052 685778
rect 213000 685714 213052 685720
rect 199844 685704 199896 685710
rect 199844 685646 199896 685652
rect 186688 685568 186740 685574
rect 186688 685510 186740 685516
rect 173532 685364 173584 685370
rect 173532 685306 173584 685312
rect 173544 683890 173572 685306
rect 177856 684888 177908 684894
rect 177856 684830 177908 684836
rect 177868 683890 177896 684830
rect 186700 683890 186728 685510
rect 191012 685160 191064 685166
rect 191012 685102 191064 685108
rect 191024 683890 191052 685102
rect 195106 684140 195158 684146
rect 195106 684082 195158 684088
rect 164252 683862 164404 683890
rect 168392 683862 168820 683890
rect 173236 683862 173572 683890
rect 177560 683862 177896 683890
rect 186392 683862 186728 683890
rect 190716 683862 191052 683890
rect 195118 683876 195146 684082
rect 199856 683890 199884 685646
rect 204168 685296 204220 685302
rect 204168 685238 204220 685244
rect 204180 683890 204208 685238
rect 208308 684276 208360 684282
rect 208308 684218 208360 684224
rect 208320 683890 208348 684218
rect 213012 683890 213040 685714
rect 217416 685500 217468 685506
rect 217416 685442 217468 685448
rect 217428 683890 217456 685442
rect 221740 684480 221792 684486
rect 221740 684422 221792 684428
rect 221752 683890 221780 684422
rect 226168 683890 226196 685782
rect 199548 683862 199884 683890
rect 203872 683862 204208 683890
rect 208288 683862 208348 683890
rect 212704 683862 213040 683890
rect 217120 683862 217456 683890
rect 221444 683862 221780 683890
rect 225860 683862 226196 683890
rect 229940 683890 229968 686938
rect 233252 685545 233280 686938
rect 233238 685536 233294 685545
rect 233238 685471 233294 685480
rect 234632 683890 234660 686938
rect 229940 683862 230276 683890
rect 234600 683862 234660 683890
rect 238772 683890 238800 687890
rect 242912 683890 242940 690678
rect 247052 684570 247080 690678
rect 251180 688016 251232 688022
rect 251180 687958 251232 687964
rect 247052 684542 247356 684570
rect 247328 683890 247356 684542
rect 251192 684026 251220 687958
rect 255332 684026 255360 690678
rect 260852 684162 260880 690678
rect 264980 688152 265032 688158
rect 264980 688094 265032 688100
rect 260852 684134 260926 684162
rect 251192 683998 251772 684026
rect 255332 683998 256096 684026
rect 251744 683890 251772 683998
rect 238772 683862 239016 683890
rect 242912 683862 243432 683890
rect 247328 683862 247756 683890
rect 251744 683862 252172 683890
rect 256068 683754 256096 683998
rect 260898 683876 260926 684134
rect 264992 683890 265020 688094
rect 269132 684570 269160 690678
rect 269132 684542 269344 684570
rect 269316 683890 269344 684542
rect 264992 683862 265328 683890
rect 269316 683862 269744 683890
rect 273272 683754 273300 690678
rect 278688 688288 278740 688294
rect 278688 688230 278740 688236
rect 277306 684312 277362 684321
rect 277306 684247 277362 684256
rect 276938 684040 276994 684049
rect 276938 683975 276994 683984
rect 142508 683738 142844 683754
rect 142508 683732 142856 683738
rect 142508 683726 142804 683732
rect 256068 683726 256588 683754
rect 273272 683726 274068 683754
rect 142804 683674 142856 683680
rect 182088 683664 182140 683670
rect 138092 683602 138428 683618
rect 181976 683612 182088 683618
rect 181976 683606 182140 683612
rect 138092 683596 138440 683602
rect 138092 683590 138388 683596
rect 181976 683590 182128 683606
rect 138388 683538 138440 683544
rect 276952 683369 276980 683975
rect 277320 683369 277348 684247
rect 278700 683890 278728 688230
rect 284220 687274 284248 699858
rect 283196 687268 283248 687274
rect 283196 687210 283248 687216
rect 284208 687268 284260 687274
rect 284208 687210 284260 687216
rect 280618 684040 280674 684049
rect 280618 683975 280674 683984
rect 278484 683862 278728 683890
rect 280632 683369 280660 683975
rect 283208 683890 283236 687210
rect 288360 684026 288388 699926
rect 295340 699848 295392 699854
rect 295340 699790 295392 699796
rect 291936 688424 291988 688430
rect 291936 688366 291988 688372
rect 282900 683862 283236 683890
rect 287716 683998 288388 684026
rect 287716 683754 287744 683998
rect 291948 683890 291976 688366
rect 291640 683862 291976 683890
rect 287224 683726 287744 683754
rect 295352 683754 295380 699790
rect 299480 699780 299532 699786
rect 299480 699722 299532 699728
rect 298190 684312 298246 684321
rect 298190 684247 298246 684256
rect 298098 684176 298154 684185
rect 298098 684111 298154 684120
rect 298112 684026 298140 684111
rect 298204 684026 298232 684247
rect 298112 683998 298232 684026
rect 299492 684026 299520 699722
rect 300228 692850 300256 703446
rect 325700 701004 325752 701010
rect 325700 700946 325752 700952
rect 321560 700936 321612 700942
rect 321560 700878 321612 700884
rect 309140 700120 309192 700126
rect 309140 700062 309192 700068
rect 299572 692844 299624 692850
rect 299572 692786 299624 692792
rect 300216 692844 300268 692850
rect 300216 692786 300268 692792
rect 299584 688430 299612 692786
rect 299572 688424 299624 688430
rect 299572 688366 299624 688372
rect 304448 688356 304500 688362
rect 304448 688298 304500 688304
rect 302146 684312 302202 684321
rect 302202 684270 302280 684298
rect 302146 684247 302202 684256
rect 302252 684185 302280 684270
rect 302238 684176 302294 684185
rect 302238 684111 302294 684120
rect 299492 683998 299980 684026
rect 299952 683890 299980 683998
rect 304460 683890 304488 688298
rect 309152 684162 309180 700062
rect 313280 700052 313332 700058
rect 313280 699994 313332 700000
rect 312450 684176 312506 684185
rect 309152 684134 309226 684162
rect 299952 683862 300380 683890
rect 304460 683862 304796 683890
rect 309198 683876 309226 684134
rect 312450 684111 312506 684120
rect 311162 684040 311218 684049
rect 311162 683975 311218 683984
rect 295352 683726 296056 683754
rect 311176 683369 311204 683975
rect 312464 683369 312492 684111
rect 313002 684040 313058 684049
rect 313002 683975 313058 683984
rect 313016 683369 313044 683975
rect 313292 683890 313320 699994
rect 317604 688220 317656 688226
rect 317604 688162 317656 688168
rect 317616 683890 317644 688162
rect 318798 684176 318854 684185
rect 318798 684111 318854 684120
rect 313292 683862 313536 683890
rect 317616 683862 317952 683890
rect 318812 683369 318840 684111
rect 321572 684026 321600 700878
rect 321572 683998 321876 684026
rect 321848 683754 321876 683998
rect 325712 683754 325740 700946
rect 332520 699922 332548 703520
rect 339500 700732 339552 700738
rect 339500 700674 339552 700680
rect 335360 700664 335412 700670
rect 335360 700606 335412 700612
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 330760 688084 330812 688090
rect 330760 688026 330812 688032
rect 328366 684176 328422 684185
rect 328366 684111 328422 684120
rect 321848 683726 322368 683754
rect 325712 683726 326692 683754
rect 328380 683482 328408 684111
rect 328458 684040 328514 684049
rect 328458 683975 328514 683984
rect 328472 683482 328500 683975
rect 330772 683890 330800 688026
rect 333242 684176 333298 684185
rect 333242 684111 333298 684120
rect 330772 683862 331108 683890
rect 331218 683768 331274 683777
rect 331402 683768 331458 683777
rect 331274 683726 331402 683754
rect 331218 683703 331274 683712
rect 331402 683703 331458 683712
rect 331218 683632 331274 683641
rect 331402 683632 331458 683641
rect 331274 683590 331402 683618
rect 331218 683567 331274 683576
rect 331402 683567 331458 683576
rect 328380 683454 328500 683482
rect 331218 683496 331274 683505
rect 331402 683496 331458 683505
rect 331274 683454 331402 683482
rect 331218 683431 331274 683440
rect 331402 683431 331458 683440
rect 333256 683369 333284 684111
rect 333426 684040 333482 684049
rect 333426 683975 333482 683984
rect 333440 683369 333468 683975
rect 335372 683890 335400 700606
rect 339512 683890 339540 700674
rect 343640 700460 343692 700466
rect 343640 700402 343692 700408
rect 335372 683862 335524 683890
rect 339512 683862 339848 683890
rect 343652 683754 343680 700402
rect 347780 700324 347832 700330
rect 347780 700266 347832 700272
rect 347792 683754 347820 700266
rect 348804 699990 348832 703520
rect 364996 703474 365024 703520
rect 364996 703446 365116 703474
rect 351920 700392 351972 700398
rect 351920 700334 351972 700340
rect 348792 699984 348844 699990
rect 348792 699926 348844 699932
rect 351932 684026 351960 700334
rect 365088 692850 365116 703446
rect 397472 700194 397500 703520
rect 413664 700262 413692 703520
rect 429856 703474 429884 703520
rect 429856 703446 429976 703474
rect 413652 700256 413704 700262
rect 413652 700198 413704 700204
rect 397460 700188 397512 700194
rect 397460 700130 397512 700136
rect 429948 692850 429976 703446
rect 462332 700874 462360 703520
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 478524 700806 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 494900 692850 494928 703446
rect 527192 700602 527220 703520
rect 527180 700596 527232 700602
rect 527180 700538 527232 700544
rect 543476 700534 543504 703520
rect 559668 703474 559696 703520
rect 559668 703446 559788 703474
rect 543464 700528 543516 700534
rect 543464 700470 543516 700476
rect 559760 692850 559788 703446
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 364340 692844 364392 692850
rect 364340 692786 364392 692792
rect 365076 692844 365128 692850
rect 365076 692786 365128 692792
rect 429200 692844 429252 692850
rect 429200 692786 429252 692792
rect 429936 692844 429988 692850
rect 429936 692786 429988 692792
rect 494060 692844 494112 692850
rect 494060 692786 494112 692792
rect 494888 692844 494940 692850
rect 494888 692786 494940 692792
rect 558920 692844 558972 692850
rect 558920 692786 558972 692792
rect 559748 692844 559800 692850
rect 559748 692786 559800 692792
rect 364352 688294 364380 692786
rect 364340 688288 364392 688294
rect 364340 688230 364392 688236
rect 429212 688158 429240 692786
rect 429200 688152 429252 688158
rect 429200 688094 429252 688100
rect 494072 688022 494100 692786
rect 494060 688016 494112 688022
rect 494060 687958 494112 687964
rect 558932 687954 558960 692786
rect 558920 687948 558972 687954
rect 558920 687890 558972 687896
rect 379428 687200 379480 687206
rect 379428 687142 379480 687148
rect 480258 687168 480314 687177
rect 365904 687132 365956 687138
rect 365904 687074 365956 687080
rect 357440 685636 357492 685642
rect 357440 685578 357492 685584
rect 356624 685086 357388 685114
rect 356624 685001 356652 685086
rect 357360 685001 357388 685086
rect 356610 684992 356666 685001
rect 356610 684927 356666 684936
rect 357346 684992 357402 685001
rect 357346 684927 357402 684936
rect 356978 684856 357034 684865
rect 357346 684856 357402 684865
rect 357034 684814 357346 684842
rect 356978 684791 357034 684800
rect 357346 684791 357402 684800
rect 357162 684720 357218 684729
rect 357346 684720 357402 684729
rect 357218 684678 357346 684706
rect 357162 684655 357218 684664
rect 357346 684655 357402 684664
rect 357346 684448 357402 684457
rect 357346 684383 357402 684392
rect 357360 684185 357388 684383
rect 357346 684176 357402 684185
rect 357346 684111 357402 684120
rect 351932 683998 352512 684026
rect 352484 683754 352512 683998
rect 357452 683890 357480 685578
rect 361580 684412 361632 684418
rect 361580 684354 361632 684360
rect 360106 684312 360162 684321
rect 360106 684247 360162 684256
rect 360120 684049 360148 684247
rect 360106 684040 360162 684049
rect 360106 683975 360162 683984
rect 357420 683862 357480 683890
rect 361592 683890 361620 684354
rect 365916 684350 365944 687074
rect 370228 685432 370280 685438
rect 370228 685374 370280 685380
rect 365812 684344 365864 684350
rect 365812 684286 365864 684292
rect 365904 684344 365956 684350
rect 365904 684286 365956 684292
rect 367006 684312 367062 684321
rect 365824 683890 365852 684286
rect 367006 684247 367062 684256
rect 367020 684049 367048 684247
rect 367006 684040 367062 684049
rect 367006 683975 367062 683984
rect 370240 683890 370268 685374
rect 379334 684312 379390 684321
rect 379334 684247 379390 684256
rect 379348 684214 379376 684247
rect 374644 684208 374696 684214
rect 374644 684150 374696 684156
rect 379336 684208 379388 684214
rect 379336 684150 379388 684156
rect 379440 684162 379468 687142
rect 480258 687103 480314 687112
rect 411168 687064 411220 687070
rect 411168 687006 411220 687012
rect 405740 686724 405792 686730
rect 405740 686666 405792 686672
rect 383752 685228 383804 685234
rect 383752 685170 383804 685176
rect 374656 683890 374684 684150
rect 379440 684134 379560 684162
rect 361592 683862 361836 683890
rect 365824 683862 366160 683890
rect 370240 683862 370576 683890
rect 374656 683862 374992 683890
rect 379072 683874 379408 683890
rect 379532 683874 379560 684134
rect 383764 683890 383792 685170
rect 396540 685024 396592 685030
rect 396540 684966 396592 684972
rect 386326 684312 386382 684321
rect 386326 684247 386382 684256
rect 386340 684214 386368 684247
rect 386328 684208 386380 684214
rect 386328 684150 386380 684156
rect 387800 684072 387852 684078
rect 387800 684014 387852 684020
rect 379060 683868 379408 683874
rect 379112 683862 379408 683868
rect 379520 683868 379572 683874
rect 379060 683810 379112 683816
rect 383732 683862 383792 683890
rect 387812 683890 387840 684014
rect 392216 684004 392268 684010
rect 392216 683946 392268 683952
rect 392228 683890 392256 683946
rect 396552 683890 396580 684966
rect 398748 684412 398800 684418
rect 398748 684354 398800 684360
rect 405648 684412 405700 684418
rect 405648 684354 405700 684360
rect 398760 684321 398788 684354
rect 405660 684321 405688 684354
rect 398746 684312 398802 684321
rect 398746 684247 398802 684256
rect 405646 684312 405702 684321
rect 405646 684247 405702 684256
rect 400956 683936 401008 683942
rect 387812 683862 388148 683890
rect 392228 683862 392564 683890
rect 396552 683862 396888 683890
rect 405752 683890 405780 686666
rect 411180 685234 411208 687006
rect 418528 686588 418580 686594
rect 418528 686530 418580 686536
rect 411168 685228 411220 685234
rect 411168 685170 411220 685176
rect 414112 685092 414164 685098
rect 414112 685034 414164 685040
rect 409880 684820 409932 684826
rect 409880 684762 409932 684768
rect 401008 683884 401304 683890
rect 400956 683878 401304 683884
rect 400968 683862 401304 683878
rect 405720 683862 405780 683890
rect 409892 683890 409920 684762
rect 414124 683890 414152 685034
rect 418068 684412 418120 684418
rect 418068 684354 418120 684360
rect 418080 684321 418108 684354
rect 418066 684312 418122 684321
rect 418066 684247 418122 684256
rect 418540 683890 418568 686530
rect 444840 686384 444892 686390
rect 444840 686326 444892 686332
rect 440424 686316 440476 686322
rect 440424 686258 440476 686264
rect 422852 684752 422904 684758
rect 422852 684694 422904 684700
rect 422864 683890 422892 684694
rect 436100 684548 436152 684554
rect 436100 684490 436152 684496
rect 424968 684412 425020 684418
rect 424968 684354 425020 684360
rect 424980 684321 425008 684354
rect 424966 684312 425022 684321
rect 424966 684247 425022 684256
rect 436112 683890 436140 684490
rect 437388 684412 437440 684418
rect 437388 684354 437440 684360
rect 437400 684321 437428 684354
rect 437386 684312 437442 684321
rect 437386 684247 437442 684256
rect 440436 683890 440464 686258
rect 444288 684412 444340 684418
rect 444288 684354 444340 684360
rect 444300 684321 444328 684354
rect 444286 684312 444342 684321
rect 444286 684247 444342 684256
rect 444852 683890 444880 686326
rect 453580 686180 453632 686186
rect 453580 686122 453632 686128
rect 449164 684616 449216 684622
rect 449164 684558 449216 684564
rect 449176 683890 449204 684558
rect 453592 683890 453620 686122
rect 471152 686112 471204 686118
rect 471152 686054 471204 686060
rect 462318 685128 462374 685137
rect 462318 685063 462374 685072
rect 456708 684412 456760 684418
rect 456708 684354 456760 684360
rect 456720 684321 456748 684354
rect 456706 684312 456762 684321
rect 456706 684247 456762 684256
rect 462332 683890 462360 685063
rect 463608 684412 463660 684418
rect 463608 684354 463660 684360
rect 463620 684321 463648 684354
rect 463606 684312 463662 684321
rect 463606 684247 463662 684256
rect 471164 683890 471192 686054
rect 476026 684312 476082 684321
rect 476026 684247 476082 684256
rect 476040 684214 476068 684247
rect 476028 684208 476080 684214
rect 476028 684150 476080 684156
rect 480272 683890 480300 687103
rect 580078 687032 580134 687041
rect 580078 686967 580134 686976
rect 580172 686996 580224 687002
rect 539324 686928 539376 686934
rect 506570 686896 506626 686905
rect 539324 686870 539376 686876
rect 506570 686831 506626 686840
rect 484400 685976 484452 685982
rect 484400 685918 484452 685924
rect 482926 684312 482982 684321
rect 482926 684247 482982 684256
rect 482940 684214 482968 684247
rect 482928 684208 482980 684214
rect 482928 684150 482980 684156
rect 409892 683862 410044 683890
rect 414124 683862 414460 683890
rect 418540 683862 418876 683890
rect 422864 683862 423200 683890
rect 436112 683862 436356 683890
rect 440436 683862 440772 683890
rect 444852 683862 445188 683890
rect 449176 683862 449512 683890
rect 453592 683862 453928 683890
rect 462332 683862 462668 683890
rect 471164 683862 471500 683890
rect 480240 683862 480300 683890
rect 484412 683890 484440 685918
rect 488630 685264 488686 685273
rect 488630 685199 488686 685208
rect 488644 683890 488672 685199
rect 501786 684720 501842 684729
rect 501786 684655 501842 684664
rect 495346 684312 495402 684321
rect 495346 684247 495402 684256
rect 495360 684078 495388 684247
rect 495348 684072 495400 684078
rect 495348 684014 495400 684020
rect 497924 684072 497976 684078
rect 497924 684014 497976 684020
rect 493046 683904 493102 683913
rect 484412 683862 484656 683890
rect 488644 683862 488980 683890
rect 493102 683862 493396 683890
rect 493046 683839 493102 683848
rect 379520 683810 379572 683816
rect 427268 683800 427320 683806
rect 343652 683726 344264 683754
rect 347792 683726 348680 683754
rect 352484 683726 353004 683754
rect 427320 683748 427616 683754
rect 427268 683742 427616 683748
rect 427280 683726 427616 683742
rect 497936 683641 497964 684014
rect 501800 683890 501828 684655
rect 506584 683890 506612 686831
rect 539048 686656 539100 686662
rect 510618 686624 510674 686633
rect 539048 686598 539100 686604
rect 510618 686559 510674 686568
rect 501800 683862 502136 683890
rect 506552 683862 506612 683890
rect 509238 683904 509294 683913
rect 510632 683890 510660 686559
rect 538956 686520 539008 686526
rect 538956 686462 539008 686468
rect 538864 686452 538916 686458
rect 538864 686394 538916 686400
rect 528098 686216 528154 686225
rect 528098 686151 528154 686160
rect 528112 683890 528140 686151
rect 510632 683862 510968 683890
rect 528112 683862 528448 683890
rect 509238 683839 509294 683848
rect 509252 683641 509280 683839
rect 514942 683768 514998 683777
rect 514998 683726 515292 683754
rect 514942 683703 514998 683712
rect 497462 683632 497518 683641
rect 497922 683632 497978 683641
rect 497518 683590 497812 683618
rect 497462 683567 497518 683576
rect 497922 683567 497978 683576
rect 509238 683632 509294 683641
rect 509238 683567 509294 683576
rect 532698 683632 532754 683641
rect 532754 683590 532864 683618
rect 532698 683567 532754 683576
rect 431868 683528 431920 683534
rect 519358 683496 519414 683505
rect 431920 683476 432032 683482
rect 431868 683470 432032 683476
rect 431880 683454 432032 683470
rect 466748 683466 467084 683482
rect 466736 683460 467084 683466
rect 466788 683454 467084 683460
rect 519414 683454 519708 683482
rect 519358 683431 519414 683440
rect 466736 683402 466788 683408
rect 458180 683392 458232 683398
rect 276938 683360 276994 683369
rect 89870 683262 89898 683332
rect 98610 683262 98638 683332
rect 276938 683295 276994 683304
rect 277306 683360 277362 683369
rect 277306 683295 277362 683304
rect 280618 683360 280674 683369
rect 280618 683295 280674 683304
rect 311162 683360 311218 683369
rect 311162 683295 311218 683304
rect 312450 683360 312506 683369
rect 312450 683295 312506 683304
rect 313002 683360 313058 683369
rect 313002 683295 313058 683304
rect 318798 683360 318854 683369
rect 318798 683295 318854 683304
rect 333242 683360 333298 683369
rect 333242 683295 333298 683304
rect 333426 683360 333482 683369
rect 521658 683360 521714 683369
rect 458232 683340 458344 683346
rect 458180 683334 458344 683340
rect 458192 683318 458344 683334
rect 475488 683330 475824 683346
rect 475476 683324 475824 683330
rect 333426 683295 333482 683304
rect 475528 683318 475824 683324
rect 523788 683330 524124 683346
rect 521658 683295 521660 683304
rect 475476 683266 475528 683272
rect 521712 683295 521714 683304
rect 523776 683324 524124 683330
rect 521660 683266 521712 683272
rect 523828 683318 524124 683324
rect 537280 683318 538260 683346
rect 523776 683266 523828 683272
rect 89858 683256 89910 683262
rect 89858 683198 89910 683204
rect 98598 683256 98650 683262
rect 98598 683198 98650 683204
rect 113560 64246 114448 64274
rect 40020 64110 40264 64138
rect 39948 61124 40000 61130
rect 39948 61066 40000 61072
rect 39856 30320 39908 30326
rect 39856 30262 39908 30268
rect 39960 626 39988 61066
rect 40132 59696 40184 59702
rect 40132 59638 40184 59644
rect 40144 3534 40172 59638
rect 40132 3528 40184 3534
rect 40132 3470 40184 3476
rect 40236 3466 40264 64110
rect 40696 64110 41032 64138
rect 41432 64110 42044 64138
rect 42812 64110 43056 64138
rect 43456 64110 44068 64138
rect 44744 64110 45080 64138
rect 45572 64110 46092 64138
rect 46952 64110 47104 64138
rect 47780 64110 48116 64138
rect 48792 64110 49128 64138
rect 49712 64110 50140 64138
rect 51092 64110 51244 64138
rect 51920 64110 52256 64138
rect 52932 64110 53268 64138
rect 53852 64110 54280 64138
rect 55292 64110 55352 64138
rect 40696 59702 40724 64110
rect 40776 60852 40828 60858
rect 40776 60794 40828 60800
rect 40684 59696 40736 59702
rect 40684 59638 40736 59644
rect 40788 58018 40816 60794
rect 40696 57990 40816 58018
rect 40696 3942 40724 57990
rect 40960 5228 41012 5234
rect 40960 5170 41012 5176
rect 40684 3936 40736 3942
rect 40684 3878 40736 3884
rect 40224 3460 40276 3466
rect 40224 3402 40276 3408
rect 38488 598 38608 626
rect 38580 480 38608 598
rect 39776 598 39988 626
rect 39776 480 39804 598
rect 40972 480 41000 5170
rect 41432 3602 41460 64110
rect 42812 61402 42840 64110
rect 43456 61554 43484 64110
rect 42904 61526 43484 61554
rect 42800 61396 42852 61402
rect 42800 61338 42852 61344
rect 42708 60920 42760 60926
rect 42708 60862 42760 60868
rect 42720 4146 42748 60862
rect 42904 60722 42932 61526
rect 44744 61470 44772 64110
rect 44732 61464 44784 61470
rect 44732 61406 44784 61412
rect 43444 61396 43496 61402
rect 43444 61338 43496 61344
rect 42892 60716 42944 60722
rect 42892 60658 42944 60664
rect 43076 60716 43128 60722
rect 43076 60658 43128 60664
rect 43088 57934 43116 60658
rect 42800 57928 42852 57934
rect 42800 57870 42852 57876
rect 43076 57928 43128 57934
rect 43076 57870 43128 57876
rect 42812 48346 42840 57870
rect 42800 48340 42852 48346
rect 42800 48282 42852 48288
rect 42984 48340 43036 48346
rect 42984 48282 43036 48288
rect 42996 41478 43024 48282
rect 42984 41472 43036 41478
rect 42984 41414 43036 41420
rect 42984 41336 43036 41342
rect 42984 41278 43036 41284
rect 42996 38690 43024 41278
rect 42892 38684 42944 38690
rect 42892 38626 42944 38632
rect 42984 38684 43036 38690
rect 42984 38626 43036 38632
rect 42904 33998 42932 38626
rect 42892 33992 42944 33998
rect 42892 33934 42944 33940
rect 43260 33992 43312 33998
rect 43260 33934 43312 33940
rect 43272 29034 43300 33934
rect 43076 29028 43128 29034
rect 43076 28970 43128 28976
rect 43260 29028 43312 29034
rect 43260 28970 43312 28976
rect 43088 22250 43116 28970
rect 42996 22222 43116 22250
rect 42996 19378 43024 22222
rect 42892 19372 42944 19378
rect 42892 19314 42944 19320
rect 42984 19372 43036 19378
rect 42984 19314 43036 19320
rect 42904 12458 42932 19314
rect 42904 12430 43024 12458
rect 42156 4140 42208 4146
rect 42156 4082 42208 4088
rect 42708 4140 42760 4146
rect 42708 4082 42760 4088
rect 41420 3596 41472 3602
rect 41420 3538 41472 3544
rect 42168 480 42196 4082
rect 42996 3670 43024 12430
rect 43456 3738 43484 61338
rect 45572 4826 45600 64110
rect 46952 61606 46980 64110
rect 47780 61742 47808 64110
rect 47768 61736 47820 61742
rect 47768 61678 47820 61684
rect 46940 61600 46992 61606
rect 46940 61542 46992 61548
rect 46848 61464 46900 61470
rect 46848 61406 46900 61412
rect 45560 4820 45612 4826
rect 45560 4762 45612 4768
rect 43444 3732 43496 3738
rect 43444 3674 43496 3680
rect 44548 3732 44600 3738
rect 44548 3674 44600 3680
rect 42984 3664 43036 3670
rect 42984 3606 43036 3612
rect 43352 3460 43404 3466
rect 43352 3402 43404 3408
rect 43364 480 43392 3402
rect 44560 480 44588 3674
rect 46860 3534 46888 61406
rect 48792 61402 48820 64110
rect 49608 61600 49660 61606
rect 49608 61542 49660 61548
rect 48780 61396 48832 61402
rect 48780 61338 48832 61344
rect 47584 60784 47636 60790
rect 47584 60726 47636 60732
rect 47400 4820 47452 4826
rect 47400 4762 47452 4768
rect 46940 3936 46992 3942
rect 46940 3878 46992 3884
rect 45744 3528 45796 3534
rect 45744 3470 45796 3476
rect 46848 3528 46900 3534
rect 46848 3470 46900 3476
rect 45756 480 45784 3470
rect 46952 480 46980 3878
rect 47412 3738 47440 4762
rect 47596 4010 47624 60726
rect 47584 4004 47636 4010
rect 47584 3946 47636 3952
rect 47400 3732 47452 3738
rect 47400 3674 47452 3680
rect 48136 3392 48188 3398
rect 48136 3334 48188 3340
rect 48148 480 48176 3334
rect 49620 626 49648 61542
rect 49712 4962 49740 64110
rect 51092 61538 51120 64110
rect 51920 61810 51948 64110
rect 51908 61804 51960 61810
rect 51908 61746 51960 61752
rect 52932 61674 52960 64110
rect 53748 61736 53800 61742
rect 53748 61678 53800 61684
rect 52920 61668 52972 61674
rect 52920 61610 52972 61616
rect 51080 61532 51132 61538
rect 51080 61474 51132 61480
rect 50988 61396 51040 61402
rect 50988 61338 51040 61344
rect 49700 4956 49752 4962
rect 49700 4898 49752 4904
rect 51000 4146 51028 61338
rect 50528 4140 50580 4146
rect 50528 4082 50580 4088
rect 50988 4140 51040 4146
rect 50988 4082 51040 4088
rect 49344 598 49648 626
rect 49344 480 49372 598
rect 50540 480 50568 4082
rect 51632 3664 51684 3670
rect 51632 3606 51684 3612
rect 51644 480 51672 3606
rect 53760 3466 53788 61678
rect 53852 4894 53880 64110
rect 55324 61946 55352 64110
rect 55968 64110 56304 64138
rect 56980 64110 57316 64138
rect 57992 64110 58328 64138
rect 59340 64110 59400 64138
rect 55312 61940 55364 61946
rect 55312 61882 55364 61888
rect 55128 61532 55180 61538
rect 55128 61474 55180 61480
rect 53840 4888 53892 4894
rect 53840 4830 53892 4836
rect 55140 3602 55168 61474
rect 55968 60858 55996 64110
rect 56508 61804 56560 61810
rect 56508 61746 56560 61752
rect 55956 60852 56008 60858
rect 55956 60794 56008 60800
rect 54024 3596 54076 3602
rect 54024 3538 54076 3544
rect 55128 3596 55180 3602
rect 55128 3538 55180 3544
rect 52828 3460 52880 3466
rect 52828 3402 52880 3408
rect 53748 3460 53800 3466
rect 53748 3402 53800 3408
rect 52840 480 52868 3402
rect 54036 480 54064 3538
rect 56520 3482 56548 61746
rect 56980 60790 57008 64110
rect 57888 61668 57940 61674
rect 57888 61610 57940 61616
rect 56968 60784 57020 60790
rect 56968 60726 57020 60732
rect 56428 3454 56548 3482
rect 55220 3392 55272 3398
rect 55220 3334 55272 3340
rect 55232 480 55260 3334
rect 56428 480 56456 3454
rect 57900 626 57928 61610
rect 57992 5030 58020 64110
rect 59372 61878 59400 64110
rect 60016 64110 60352 64138
rect 61028 64110 61364 64138
rect 62132 64110 62468 64138
rect 63480 64110 63540 64138
rect 60016 62014 60044 64110
rect 61028 62082 61056 64110
rect 61016 62076 61068 62082
rect 61016 62018 61068 62024
rect 60004 62008 60056 62014
rect 60004 61950 60056 61956
rect 60648 62008 60700 62014
rect 60648 61950 60700 61956
rect 59912 61940 59964 61946
rect 59912 61882 59964 61888
rect 59360 61872 59412 61878
rect 59360 61814 59412 61820
rect 59924 61198 59952 61882
rect 59912 61192 59964 61198
rect 59912 61134 59964 61140
rect 60004 60784 60056 60790
rect 60004 60726 60056 60732
rect 57980 5024 58032 5030
rect 57980 4966 58032 4972
rect 60016 3806 60044 60726
rect 60004 3800 60056 3806
rect 60004 3742 60056 3748
rect 58808 3732 58860 3738
rect 58808 3674 58860 3680
rect 57624 598 57928 626
rect 57624 480 57652 598
rect 58820 480 58848 3674
rect 60660 3602 60688 61950
rect 62028 61872 62080 61878
rect 62028 61814 62080 61820
rect 62040 3602 62068 61814
rect 62132 5098 62160 64110
rect 63512 61266 63540 64110
rect 64248 64110 64492 64138
rect 64892 64110 65504 64138
rect 66272 64110 66516 64138
rect 67192 64110 67528 64138
rect 67652 64110 68540 64138
rect 69216 64110 69552 64138
rect 70412 64110 70564 64138
rect 70688 64110 71576 64138
rect 72252 64110 72588 64138
rect 73356 64110 73692 64138
rect 74704 64110 74856 64138
rect 63500 61260 63552 61266
rect 63500 61202 63552 61208
rect 64144 61260 64196 61266
rect 64144 61202 64196 61208
rect 62120 5092 62172 5098
rect 62120 5034 62172 5040
rect 64156 3874 64184 61202
rect 64248 60790 64276 64110
rect 64788 62076 64840 62082
rect 64788 62018 64840 62024
rect 64236 60784 64288 60790
rect 64236 60726 64288 60732
rect 64696 4004 64748 4010
rect 64696 3946 64748 3952
rect 64144 3868 64196 3874
rect 64144 3810 64196 3816
rect 62396 3800 62448 3806
rect 62396 3742 62448 3748
rect 60004 3596 60056 3602
rect 60004 3538 60056 3544
rect 60648 3596 60700 3602
rect 60648 3538 60700 3544
rect 61200 3596 61252 3602
rect 61200 3538 61252 3544
rect 62028 3596 62080 3602
rect 62028 3538 62080 3544
rect 62120 3596 62172 3602
rect 62120 3538 62172 3544
rect 60016 480 60044 3538
rect 61212 480 61240 3538
rect 62132 3398 62160 3538
rect 62120 3392 62172 3398
rect 62120 3334 62172 3340
rect 62408 480 62436 3742
rect 63592 3392 63644 3398
rect 63592 3334 63644 3340
rect 63604 480 63632 3334
rect 64708 1986 64736 3946
rect 64800 3398 64828 62018
rect 64892 5166 64920 64110
rect 66272 61334 66300 64110
rect 67192 61946 67220 64110
rect 67180 61940 67232 61946
rect 67180 61882 67232 61888
rect 66260 61328 66312 61334
rect 66260 61270 66312 61276
rect 67548 61328 67600 61334
rect 67548 61270 67600 61276
rect 64880 5160 64932 5166
rect 64880 5102 64932 5108
rect 65984 4888 66036 4894
rect 65984 4830 66036 4836
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 64708 1958 64828 1986
rect 64800 480 64828 1958
rect 65996 480 66024 4830
rect 67560 3380 67588 61270
rect 67652 5302 67680 64110
rect 68928 61940 68980 61946
rect 68928 61882 68980 61888
rect 68284 60852 68336 60858
rect 68284 60794 68336 60800
rect 67640 5296 67692 5302
rect 67640 5238 67692 5244
rect 68296 4010 68324 60794
rect 68284 4004 68336 4010
rect 68284 3946 68336 3952
rect 68940 3398 68968 61882
rect 69216 60994 69244 64110
rect 70412 61266 70440 64110
rect 70400 61260 70452 61266
rect 70400 61202 70452 61208
rect 69204 60988 69256 60994
rect 69204 60930 69256 60936
rect 70688 5370 70716 64110
rect 71596 61192 71648 61198
rect 71596 61134 71648 61140
rect 71608 60994 71636 61134
rect 72252 61062 72280 64110
rect 73068 61260 73120 61266
rect 73068 61202 73120 61208
rect 72240 61056 72292 61062
rect 72240 60998 72292 61004
rect 71596 60988 71648 60994
rect 71596 60930 71648 60936
rect 71688 60988 71740 60994
rect 71688 60930 71740 60936
rect 70676 5364 70728 5370
rect 70676 5306 70728 5312
rect 69480 4956 69532 4962
rect 69480 4898 69532 4904
rect 67192 3352 67588 3380
rect 68284 3392 68336 3398
rect 67192 480 67220 3352
rect 68284 3334 68336 3340
rect 68928 3392 68980 3398
rect 68928 3334 68980 3340
rect 68296 480 68324 3334
rect 69492 480 69520 4898
rect 71700 3466 71728 60930
rect 73080 4146 73108 61202
rect 73356 61130 73384 64110
rect 74540 61464 74592 61470
rect 74540 61406 74592 61412
rect 73344 61124 73396 61130
rect 73344 61066 73396 61072
rect 74552 60926 74580 61406
rect 74540 60920 74592 60926
rect 74540 60862 74592 60868
rect 74540 56704 74592 56710
rect 74540 56646 74592 56652
rect 74552 56574 74580 56646
rect 74828 56642 74856 64110
rect 75380 64110 75716 64138
rect 76392 64110 76728 64138
rect 77312 64110 77740 64138
rect 78752 64110 78812 64138
rect 75380 61198 75408 64110
rect 75368 61192 75420 61198
rect 75368 61134 75420 61140
rect 75828 61192 75880 61198
rect 75828 61134 75880 61140
rect 75184 61124 75236 61130
rect 75184 61066 75236 61072
rect 74632 56636 74684 56642
rect 74632 56578 74684 56584
rect 74816 56636 74868 56642
rect 74816 56578 74868 56584
rect 74264 56568 74316 56574
rect 74264 56510 74316 56516
rect 74540 56568 74592 56574
rect 74540 56510 74592 56516
rect 74276 46986 74304 56510
rect 74264 46980 74316 46986
rect 74264 46922 74316 46928
rect 74448 46980 74500 46986
rect 74448 46922 74500 46928
rect 74460 37330 74488 46922
rect 74356 37324 74408 37330
rect 74356 37266 74408 37272
rect 74448 37324 74500 37330
rect 74448 37266 74500 37272
rect 74368 37194 74396 37266
rect 74356 37188 74408 37194
rect 74356 37130 74408 37136
rect 74446 27704 74502 27713
rect 74446 27639 74502 27648
rect 74460 27606 74488 27639
rect 74264 27600 74316 27606
rect 74264 27542 74316 27548
rect 74448 27600 74500 27606
rect 74448 27542 74500 27548
rect 74276 18018 74304 27542
rect 74080 18012 74132 18018
rect 74080 17954 74132 17960
rect 74264 18012 74316 18018
rect 74264 17954 74316 17960
rect 74092 9722 74120 17954
rect 74080 9716 74132 9722
rect 74080 9658 74132 9664
rect 74264 9716 74316 9722
rect 74264 9658 74316 9664
rect 71872 4140 71924 4146
rect 71872 4082 71924 4088
rect 73068 4140 73120 4146
rect 73068 4082 73120 4088
rect 70676 3460 70728 3466
rect 70676 3402 70728 3408
rect 71688 3460 71740 3466
rect 71688 3402 71740 3408
rect 70688 480 70716 3402
rect 71884 480 71912 4082
rect 72976 3868 73028 3874
rect 72976 3810 73028 3816
rect 72988 1986 73016 3810
rect 72988 1958 73108 1986
rect 73080 480 73108 1958
rect 74276 480 74304 9658
rect 74644 5234 74672 56578
rect 74724 37188 74776 37194
rect 74724 37130 74776 37136
rect 74736 27713 74764 37130
rect 74722 27704 74778 27713
rect 74722 27639 74778 27648
rect 74632 5228 74684 5234
rect 74632 5170 74684 5176
rect 75196 4026 75224 61066
rect 75276 61056 75328 61062
rect 75276 60998 75328 61004
rect 75288 56710 75316 60998
rect 75276 56704 75328 56710
rect 75276 56646 75328 56652
rect 75104 3998 75224 4026
rect 75104 3534 75132 3998
rect 75184 3936 75236 3942
rect 75184 3878 75236 3884
rect 75196 3670 75224 3878
rect 75184 3664 75236 3670
rect 75184 3606 75236 3612
rect 75092 3528 75144 3534
rect 75092 3470 75144 3476
rect 75840 626 75868 61134
rect 76392 61130 76420 64110
rect 76564 61464 76616 61470
rect 76564 61406 76616 61412
rect 76380 61124 76432 61130
rect 76380 61066 76432 61072
rect 76576 60722 76604 61406
rect 76564 60716 76616 60722
rect 76564 60658 76616 60664
rect 76748 60716 76800 60722
rect 76748 60658 76800 60664
rect 76760 57934 76788 60658
rect 76472 57928 76524 57934
rect 76472 57870 76524 57876
rect 76748 57928 76800 57934
rect 76748 57870 76800 57876
rect 76484 48346 76512 57870
rect 76472 48340 76524 48346
rect 76472 48282 76524 48288
rect 76656 48340 76708 48346
rect 76656 48282 76708 48288
rect 76668 41614 76696 48282
rect 76656 41608 76708 41614
rect 76656 41550 76708 41556
rect 76656 41472 76708 41478
rect 76656 41414 76708 41420
rect 76668 38826 76696 41414
rect 76656 38820 76708 38826
rect 76656 38762 76708 38768
rect 76564 38684 76616 38690
rect 76564 38626 76616 38632
rect 76576 31634 76604 38626
rect 76576 31606 76788 31634
rect 76760 22114 76788 31606
rect 76576 22086 76788 22114
rect 76576 12458 76604 22086
rect 76576 12430 76696 12458
rect 76668 4010 76696 12430
rect 77312 4826 77340 64110
rect 78588 61124 78640 61130
rect 78588 61066 78640 61072
rect 77300 4820 77352 4826
rect 77300 4762 77352 4768
rect 78600 4146 78628 61066
rect 78784 60926 78812 64110
rect 79428 64110 79764 64138
rect 80072 64110 80776 64138
rect 81452 64110 81788 64138
rect 82800 64110 82860 64138
rect 79428 61470 79456 64110
rect 79416 61464 79468 61470
rect 79416 61406 79468 61412
rect 78772 60920 78824 60926
rect 78772 60862 78824 60868
rect 79968 60920 80020 60926
rect 79968 60862 80020 60868
rect 79980 4146 80008 60862
rect 77852 4140 77904 4146
rect 77852 4082 77904 4088
rect 78588 4140 78640 4146
rect 78588 4082 78640 4088
rect 79048 4140 79100 4146
rect 79048 4082 79100 4088
rect 79968 4140 80020 4146
rect 79968 4082 80020 4088
rect 76656 4004 76708 4010
rect 76656 3946 76708 3952
rect 76656 3460 76708 3466
rect 76656 3402 76708 3408
rect 75472 598 75868 626
rect 75472 480 75500 598
rect 76668 480 76696 3402
rect 77864 480 77892 4082
rect 79060 480 79088 4082
rect 80072 3330 80100 64110
rect 81452 61606 81480 64110
rect 81440 61600 81492 61606
rect 81440 61542 81492 61548
rect 82636 61600 82688 61606
rect 82636 61542 82688 61548
rect 82648 3670 82676 61542
rect 82728 61464 82780 61470
rect 82728 61406 82780 61412
rect 81440 3664 81492 3670
rect 81440 3606 81492 3612
rect 82636 3664 82688 3670
rect 82636 3606 82688 3612
rect 80244 3460 80296 3466
rect 80244 3402 80296 3408
rect 80060 3324 80112 3330
rect 80060 3266 80112 3272
rect 80256 480 80284 3402
rect 81452 480 81480 3606
rect 82740 3482 82768 61406
rect 82832 61402 82860 64110
rect 83016 64110 83812 64138
rect 84580 64110 84916 64138
rect 85592 64110 85928 64138
rect 86940 64110 87000 64138
rect 82820 61396 82872 61402
rect 82820 61338 82872 61344
rect 83016 3942 83044 64110
rect 84580 61742 84608 64110
rect 84568 61736 84620 61742
rect 84568 61678 84620 61684
rect 85488 61736 85540 61742
rect 85488 61678 85540 61684
rect 83832 4072 83884 4078
rect 83832 4014 83884 4020
rect 83004 3936 83056 3942
rect 83004 3878 83056 3884
rect 82648 3454 82768 3482
rect 82648 480 82676 3454
rect 83844 480 83872 4014
rect 84844 3936 84896 3942
rect 84844 3878 84896 3884
rect 84856 3602 84884 3878
rect 85500 3602 85528 61678
rect 85592 61538 85620 64110
rect 85580 61532 85632 61538
rect 85580 61474 85632 61480
rect 86868 61396 86920 61402
rect 86868 61338 86920 61344
rect 86880 3602 86908 61338
rect 86972 3942 87000 64110
rect 87616 64110 87952 64138
rect 88628 64110 88964 64138
rect 89824 64110 89976 64138
rect 90652 64110 90988 64138
rect 91664 64110 92000 64138
rect 92492 64110 93012 64138
rect 93872 64110 94024 64138
rect 94700 64110 95036 64138
rect 95252 64110 96140 64138
rect 96816 64110 97152 64138
rect 98012 64110 98164 64138
rect 98288 64110 99176 64138
rect 99852 64110 100188 64138
rect 100864 64110 101200 64138
rect 87616 61810 87644 64110
rect 87604 61804 87656 61810
rect 87604 61746 87656 61752
rect 88628 61674 88656 64110
rect 88616 61668 88668 61674
rect 88616 61610 88668 61616
rect 89628 60784 89680 60790
rect 89628 60726 89680 60732
rect 86960 3936 87012 3942
rect 86960 3878 87012 3884
rect 87328 3936 87380 3942
rect 87328 3878 87380 3884
rect 84844 3596 84896 3602
rect 84844 3538 84896 3544
rect 84936 3596 84988 3602
rect 84936 3538 84988 3544
rect 85488 3596 85540 3602
rect 85488 3538 85540 3544
rect 86132 3596 86184 3602
rect 86132 3538 86184 3544
rect 86868 3596 86920 3602
rect 86868 3538 86920 3544
rect 84948 480 84976 3538
rect 86144 480 86172 3538
rect 87340 480 87368 3878
rect 89640 3602 89668 60726
rect 89824 3738 89852 64110
rect 90652 62014 90680 64110
rect 90640 62008 90692 62014
rect 90640 61950 90692 61956
rect 91664 61878 91692 64110
rect 91652 61872 91704 61878
rect 91652 61814 91704 61820
rect 92388 61872 92440 61878
rect 92388 61814 92440 61820
rect 91008 61668 91060 61674
rect 91008 61610 91060 61616
rect 89812 3732 89864 3738
rect 89812 3674 89864 3680
rect 90916 3732 90968 3738
rect 90916 3674 90968 3680
rect 88524 3596 88576 3602
rect 88524 3538 88576 3544
rect 89628 3596 89680 3602
rect 89628 3538 89680 3544
rect 89720 3596 89772 3602
rect 89720 3538 89772 3544
rect 88536 480 88564 3538
rect 89732 480 89760 3538
rect 90928 480 90956 3674
rect 91020 3602 91048 61610
rect 91008 3596 91060 3602
rect 91008 3538 91060 3544
rect 92400 3346 92428 61814
rect 92492 3806 92520 64110
rect 93872 62082 93900 64110
rect 93860 62076 93912 62082
rect 93860 62018 93912 62024
rect 93768 61532 93820 61538
rect 93768 61474 93820 61480
rect 92480 3800 92532 3806
rect 92480 3742 92532 3748
rect 93780 3398 93808 61474
rect 94700 60858 94728 64110
rect 94688 60852 94740 60858
rect 94688 60794 94740 60800
rect 95252 4894 95280 64110
rect 96528 62008 96580 62014
rect 96528 61950 96580 61956
rect 95240 4888 95292 4894
rect 95240 4830 95292 4836
rect 94504 3732 94556 3738
rect 94504 3674 94556 3680
rect 92124 3318 92428 3346
rect 93308 3392 93360 3398
rect 93308 3334 93360 3340
rect 93768 3392 93820 3398
rect 93768 3334 93820 3340
rect 92124 480 92152 3318
rect 93320 480 93348 3334
rect 94516 480 94544 3674
rect 96540 3398 96568 61950
rect 96816 61334 96844 64110
rect 98012 61946 98040 64110
rect 98000 61940 98052 61946
rect 98000 61882 98052 61888
rect 96804 61328 96856 61334
rect 96804 61270 96856 61276
rect 97908 61328 97960 61334
rect 97908 61270 97960 61276
rect 97920 3398 97948 61270
rect 98288 4962 98316 64110
rect 99288 61940 99340 61946
rect 99288 61882 99340 61888
rect 98276 4956 98328 4962
rect 98276 4898 98328 4904
rect 98092 4004 98144 4010
rect 98092 3946 98144 3952
rect 95700 3392 95752 3398
rect 95700 3334 95752 3340
rect 96528 3392 96580 3398
rect 96528 3334 96580 3340
rect 96896 3392 96948 3398
rect 96896 3334 96948 3340
rect 97908 3392 97960 3398
rect 97908 3334 97960 3340
rect 95712 480 95740 3334
rect 96908 480 96936 3334
rect 98104 480 98132 3946
rect 99300 480 99328 61882
rect 99852 60994 99880 64110
rect 100668 61804 100720 61810
rect 100668 61746 100720 61752
rect 99840 60988 99892 60994
rect 99840 60930 99892 60936
rect 100680 3346 100708 61746
rect 100864 61266 100892 64110
rect 102198 63866 102226 64124
rect 102152 63838 102226 63866
rect 102888 64110 103224 64138
rect 103900 64110 104236 64138
rect 104912 64110 105248 64138
rect 106260 64110 106320 64138
rect 100852 61260 100904 61266
rect 100852 61202 100904 61208
rect 102152 3874 102180 63838
rect 102888 61062 102916 64110
rect 103900 61198 103928 64110
rect 104808 61260 104860 61266
rect 104808 61202 104860 61208
rect 103888 61192 103940 61198
rect 103888 61134 103940 61140
rect 102876 61056 102928 61062
rect 102876 60998 102928 61004
rect 103428 61056 103480 61062
rect 103428 60998 103480 61004
rect 102140 3868 102192 3874
rect 102140 3810 102192 3816
rect 101588 3800 101640 3806
rect 101588 3742 101640 3748
rect 100496 3318 100708 3346
rect 100496 480 100524 3318
rect 101600 480 101628 3742
rect 103440 3398 103468 60998
rect 104820 3534 104848 61202
rect 103980 3528 104032 3534
rect 103980 3470 104032 3476
rect 104808 3528 104860 3534
rect 104808 3470 104860 3476
rect 102784 3392 102836 3398
rect 102784 3334 102836 3340
rect 103428 3392 103480 3398
rect 103428 3334 103480 3340
rect 102796 480 102824 3334
rect 103992 480 104020 3470
rect 104912 3466 104940 64110
rect 106292 61130 106320 64110
rect 107028 64110 107364 64138
rect 107672 64110 108376 64138
rect 109144 64110 109388 64138
rect 110400 64110 110460 64138
rect 106280 61124 106332 61130
rect 106280 61066 106332 61072
rect 107028 60926 107056 64110
rect 107476 62076 107528 62082
rect 107476 62018 107528 62024
rect 107016 60920 107068 60926
rect 107016 60862 107068 60868
rect 106372 3664 106424 3670
rect 106372 3606 106424 3612
rect 104900 3460 104952 3466
rect 104900 3402 104952 3408
rect 105176 3392 105228 3398
rect 105176 3334 105228 3340
rect 105188 480 105216 3334
rect 106384 480 106412 3606
rect 107488 3482 107516 62018
rect 107568 61192 107620 61198
rect 107568 61134 107620 61140
rect 107580 3670 107608 61134
rect 107568 3664 107620 3670
rect 107568 3606 107620 3612
rect 107488 3454 107608 3482
rect 107672 3466 107700 64110
rect 109144 61606 109172 64110
rect 109132 61600 109184 61606
rect 109132 61542 109184 61548
rect 110328 61600 110380 61606
rect 110328 61542 110380 61548
rect 107580 480 107608 3454
rect 107660 3460 107712 3466
rect 107660 3402 107712 3408
rect 108764 3324 108816 3330
rect 108764 3266 108816 3272
rect 108776 480 108804 3266
rect 110340 610 110368 61542
rect 110432 61470 110460 64110
rect 110524 64110 111412 64138
rect 112088 64110 112424 64138
rect 113192 64110 113436 64138
rect 110420 61464 110472 61470
rect 110420 61406 110472 61412
rect 110524 4078 110552 64110
rect 112088 61742 112116 64110
rect 112076 61736 112128 61742
rect 112076 61678 112128 61684
rect 113088 61736 113140 61742
rect 113088 61678 113140 61684
rect 111708 61464 111760 61470
rect 111708 61406 111760 61412
rect 111720 4146 111748 61406
rect 113100 4146 113128 61678
rect 113192 61402 113220 64110
rect 113560 62370 113588 64246
rect 113468 62342 113588 62370
rect 115124 64110 115460 64138
rect 116136 64110 116472 64138
rect 113180 61396 113232 61402
rect 113180 61338 113232 61344
rect 113468 51202 113496 62342
rect 114468 61124 114520 61130
rect 114468 61066 114520 61072
rect 113456 51196 113508 51202
rect 113456 51138 113508 51144
rect 113456 51060 113508 51066
rect 113456 51002 113508 51008
rect 113468 48346 113496 51002
rect 113272 48340 113324 48346
rect 113272 48282 113324 48288
rect 113456 48340 113508 48346
rect 113456 48282 113508 48288
rect 113284 41478 113312 48282
rect 113272 41472 113324 41478
rect 113272 41414 113324 41420
rect 113364 41404 113416 41410
rect 113364 41346 113416 41352
rect 113376 38622 113404 41346
rect 113180 38616 113232 38622
rect 113180 38558 113232 38564
rect 113364 38616 113416 38622
rect 113364 38558 113416 38564
rect 113192 29034 113220 38558
rect 113180 29028 113232 29034
rect 113180 28970 113232 28976
rect 113456 29028 113508 29034
rect 113456 28970 113508 28976
rect 113468 24154 113496 28970
rect 113376 24126 113496 24154
rect 111156 4140 111208 4146
rect 111156 4082 111208 4088
rect 111708 4140 111760 4146
rect 111708 4082 111760 4088
rect 112352 4140 112404 4146
rect 112352 4082 112404 4088
rect 113088 4140 113140 4146
rect 113088 4082 113140 4088
rect 110512 4072 110564 4078
rect 110512 4014 110564 4020
rect 109960 604 110012 610
rect 109960 546 110012 552
rect 110328 604 110380 610
rect 110328 546 110380 552
rect 109972 480 110000 546
rect 111168 480 111196 4082
rect 112364 480 112392 4082
rect 113376 3942 113404 24126
rect 114480 4146 114508 61066
rect 115124 60790 115152 64110
rect 116136 61674 116164 64110
rect 117470 63866 117498 64124
rect 117424 63838 117498 63866
rect 118252 64110 118588 64138
rect 119264 64110 119600 64138
rect 120092 64110 120612 64138
rect 121472 64110 121624 64138
rect 122300 64110 122636 64138
rect 122852 64110 123648 64138
rect 124324 64110 124660 64138
rect 125672 64110 125732 64138
rect 116124 61668 116176 61674
rect 116124 61610 116176 61616
rect 117228 61668 117280 61674
rect 117228 61610 117280 61616
rect 117136 60988 117188 60994
rect 117136 60930 117188 60936
rect 115848 60920 115900 60926
rect 115848 60862 115900 60868
rect 115112 60784 115164 60790
rect 115112 60726 115164 60732
rect 113548 4140 113600 4146
rect 113548 4082 113600 4088
rect 114468 4140 114520 4146
rect 114468 4082 114520 4088
rect 113364 3936 113416 3942
rect 113364 3878 113416 3884
rect 113560 480 113588 4082
rect 115860 3534 115888 60862
rect 117148 4146 117176 60930
rect 115940 4140 115992 4146
rect 115940 4082 115992 4088
rect 117136 4140 117188 4146
rect 117136 4082 117188 4088
rect 114744 3528 114796 3534
rect 114744 3470 114796 3476
rect 115848 3528 115900 3534
rect 115848 3470 115900 3476
rect 114756 480 114784 3470
rect 115952 480 115980 4082
rect 117240 4026 117268 61610
rect 117148 3998 117268 4026
rect 117148 480 117176 3998
rect 117424 3602 117452 63838
rect 118252 61878 118280 64110
rect 118240 61872 118292 61878
rect 118240 61814 118292 61820
rect 119264 61538 119292 64110
rect 119252 61532 119304 61538
rect 119252 61474 119304 61480
rect 118608 61396 118660 61402
rect 118608 61338 118660 61344
rect 117412 3596 117464 3602
rect 117412 3538 117464 3544
rect 118620 2854 118648 61338
rect 119988 60852 120040 60858
rect 119988 60794 120040 60800
rect 120000 3602 120028 60794
rect 120092 3738 120120 64110
rect 121472 62014 121500 64110
rect 121460 62008 121512 62014
rect 121460 61950 121512 61956
rect 122300 61334 122328 64110
rect 122748 61872 122800 61878
rect 122748 61814 122800 61820
rect 122288 61328 122340 61334
rect 122288 61270 122340 61276
rect 121368 60784 121420 60790
rect 121368 60726 121420 60732
rect 120080 3732 120132 3738
rect 120080 3674 120132 3680
rect 121380 3602 121408 60726
rect 122760 3602 122788 61814
rect 122852 4010 122880 64110
rect 124128 62008 124180 62014
rect 124128 61950 124180 61956
rect 122840 4004 122892 4010
rect 122840 3946 122892 3952
rect 119436 3596 119488 3602
rect 119436 3538 119488 3544
rect 119988 3596 120040 3602
rect 119988 3538 120040 3544
rect 120632 3596 120684 3602
rect 120632 3538 120684 3544
rect 121368 3596 121420 3602
rect 121368 3538 121420 3544
rect 121828 3596 121880 3602
rect 121828 3538 121880 3544
rect 122748 3596 122800 3602
rect 122748 3538 122800 3544
rect 118240 2848 118292 2854
rect 118240 2790 118292 2796
rect 118608 2848 118660 2854
rect 118608 2790 118660 2796
rect 118252 480 118280 2790
rect 119448 480 119476 3538
rect 120644 480 120672 3538
rect 121840 480 121868 3538
rect 124140 3534 124168 61950
rect 124324 61946 124352 64110
rect 124312 61940 124364 61946
rect 124312 61882 124364 61888
rect 125704 61810 125732 64110
rect 125796 64110 126684 64138
rect 127360 64110 127696 64138
rect 128372 64110 128708 64138
rect 125692 61804 125744 61810
rect 125692 61746 125744 61752
rect 125416 61532 125468 61538
rect 125416 61474 125468 61480
rect 123024 3528 123076 3534
rect 123024 3470 123076 3476
rect 124128 3528 124180 3534
rect 124128 3470 124180 3476
rect 123036 480 123064 3470
rect 124220 3324 124272 3330
rect 124220 3266 124272 3272
rect 124232 480 124260 3266
rect 125428 480 125456 61474
rect 125508 61328 125560 61334
rect 125508 61270 125560 61276
rect 125520 3330 125548 61270
rect 125796 3806 125824 64110
rect 127360 61062 127388 64110
rect 128372 61266 128400 64110
rect 129798 63866 129826 64124
rect 129752 63838 129826 63866
rect 130488 64110 130824 64138
rect 131500 64110 131836 64138
rect 132696 64110 132848 64138
rect 133860 64110 133920 64138
rect 128360 61260 128412 61266
rect 128360 61202 128412 61208
rect 129648 61260 129700 61266
rect 129648 61202 129700 61208
rect 127348 61056 127400 61062
rect 127348 60998 127400 61004
rect 125784 3800 125836 3806
rect 125784 3742 125836 3748
rect 126612 3664 126664 3670
rect 126612 3606 126664 3612
rect 125508 3324 125560 3330
rect 125508 3266 125560 3272
rect 126624 480 126652 3606
rect 127808 3596 127860 3602
rect 127808 3538 127860 3544
rect 127820 480 127848 3538
rect 129660 3534 129688 61202
rect 129752 3738 129780 63838
rect 130488 61198 130516 64110
rect 131500 62082 131528 64110
rect 131488 62076 131540 62082
rect 131488 62018 131540 62024
rect 132408 62076 132460 62082
rect 132408 62018 132460 62024
rect 130476 61192 130528 61198
rect 130476 61134 130528 61140
rect 129740 3732 129792 3738
rect 129740 3674 129792 3680
rect 129004 3528 129056 3534
rect 129004 3470 129056 3476
rect 129648 3528 129700 3534
rect 129648 3470 129700 3476
rect 130200 3528 130252 3534
rect 130200 3470 130252 3476
rect 129016 480 129044 3470
rect 130212 480 130240 3470
rect 132420 3398 132448 62018
rect 132592 3460 132644 3466
rect 132592 3402 132644 3408
rect 131396 3392 131448 3398
rect 131396 3334 131448 3340
rect 132408 3392 132460 3398
rect 132408 3334 132460 3340
rect 131408 480 131436 3334
rect 132604 480 132632 3402
rect 132696 3330 132724 64110
rect 133788 61940 133840 61946
rect 133788 61882 133840 61888
rect 133696 61804 133748 61810
rect 133696 61746 133748 61752
rect 133708 3466 133736 61746
rect 133696 3460 133748 3466
rect 133696 3402 133748 3408
rect 132684 3324 132736 3330
rect 132684 3266 132736 3272
rect 133800 480 133828 61882
rect 133892 61606 133920 64110
rect 134536 64110 134872 64138
rect 135548 64110 135884 64138
rect 136652 64110 136896 64138
rect 137572 64110 137908 64138
rect 138584 64110 138920 64138
rect 139688 64110 140024 64138
rect 140792 64110 141036 64138
rect 141712 64110 142048 64138
rect 142724 64110 143060 64138
rect 143736 64110 144072 64138
rect 144932 64110 145084 64138
rect 145760 64110 146096 64138
rect 146772 64110 147108 64138
rect 147692 64110 148120 64138
rect 133880 61600 133932 61606
rect 133880 61542 133932 61548
rect 134536 61470 134564 64110
rect 135548 61742 135576 64110
rect 135536 61736 135588 61742
rect 135536 61678 135588 61684
rect 136548 61736 136600 61742
rect 136548 61678 136600 61684
rect 135168 61600 135220 61606
rect 135168 61542 135220 61548
rect 134524 61464 134576 61470
rect 134524 61406 134576 61412
rect 135180 3482 135208 61542
rect 134904 3454 135208 3482
rect 136560 3466 136588 61678
rect 136652 61130 136680 64110
rect 136640 61124 136692 61130
rect 136640 61066 136692 61072
rect 137572 60926 137600 64110
rect 137928 61464 137980 61470
rect 137928 61406 137980 61412
rect 137560 60920 137612 60926
rect 137560 60862 137612 60868
rect 137940 3466 137968 61406
rect 138584 60994 138612 64110
rect 139688 61674 139716 64110
rect 139676 61668 139728 61674
rect 139676 61610 139728 61616
rect 140792 61402 140820 64110
rect 140780 61396 140832 61402
rect 140780 61338 140832 61344
rect 139308 61192 139360 61198
rect 139308 61134 139360 61140
rect 138572 60988 138624 60994
rect 138572 60930 138624 60936
rect 139320 3466 139348 61134
rect 140688 61056 140740 61062
rect 140688 60998 140740 61004
rect 140700 3466 140728 60998
rect 141712 60858 141740 64110
rect 142068 61668 142120 61674
rect 142068 61610 142120 61616
rect 141976 61396 142028 61402
rect 141976 61338 142028 61344
rect 141700 60852 141752 60858
rect 141700 60794 141752 60800
rect 136088 3460 136140 3466
rect 134904 480 134932 3454
rect 136088 3402 136140 3408
rect 136548 3460 136600 3466
rect 136548 3402 136600 3408
rect 137284 3460 137336 3466
rect 137284 3402 137336 3408
rect 137928 3460 137980 3466
rect 137928 3402 137980 3408
rect 138480 3460 138532 3466
rect 138480 3402 138532 3408
rect 139308 3460 139360 3466
rect 139308 3402 139360 3408
rect 139676 3460 139728 3466
rect 139676 3402 139728 3408
rect 140688 3460 140740 3466
rect 140688 3402 140740 3408
rect 136100 480 136128 3402
rect 137296 480 137324 3402
rect 138492 480 138520 3402
rect 139688 480 139716 3402
rect 140872 3052 140924 3058
rect 140872 2994 140924 3000
rect 140884 480 140912 2994
rect 141988 1578 142016 61338
rect 142080 3058 142108 61610
rect 142724 60790 142752 64110
rect 143736 61878 143764 64110
rect 144932 62014 144960 64110
rect 144920 62008 144972 62014
rect 144920 61950 144972 61956
rect 143724 61872 143776 61878
rect 143724 61814 143776 61820
rect 144828 61872 144880 61878
rect 144828 61814 144880 61820
rect 143448 61124 143500 61130
rect 143448 61066 143500 61072
rect 142712 60784 142764 60790
rect 142712 60726 142764 60732
rect 143460 3346 143488 61066
rect 144840 3346 144868 61814
rect 145760 61334 145788 64110
rect 146208 62008 146260 62014
rect 146208 61950 146260 61956
rect 145748 61328 145800 61334
rect 145748 61270 145800 61276
rect 146220 3534 146248 61950
rect 146772 61538 146800 64110
rect 146760 61532 146812 61538
rect 146760 61474 146812 61480
rect 147588 60920 147640 60926
rect 147588 60862 147640 60868
rect 147600 3534 147628 60862
rect 147692 3670 147720 64110
rect 149118 63866 149146 64124
rect 149072 63838 149146 63866
rect 149808 64110 150144 64138
rect 150636 64110 151248 64138
rect 151924 64110 152260 64138
rect 153272 64110 153332 64138
rect 148968 61328 149020 61334
rect 148968 61270 149020 61276
rect 147680 3664 147732 3670
rect 147680 3606 147732 3612
rect 148980 3534 149008 61270
rect 149072 3602 149100 63838
rect 149808 61266 149836 64110
rect 149796 61260 149848 61266
rect 149796 61202 149848 61208
rect 150348 61260 150400 61266
rect 150348 61202 150400 61208
rect 149060 3596 149112 3602
rect 149060 3538 149112 3544
rect 145656 3528 145708 3534
rect 145656 3470 145708 3476
rect 146208 3528 146260 3534
rect 146208 3470 146260 3476
rect 146852 3528 146904 3534
rect 146852 3470 146904 3476
rect 147588 3528 147640 3534
rect 147588 3470 147640 3476
rect 148048 3528 148100 3534
rect 148048 3470 148100 3476
rect 148968 3528 149020 3534
rect 148968 3470 149020 3476
rect 143276 3318 143488 3346
rect 144472 3318 144868 3346
rect 142068 3052 142120 3058
rect 142068 2994 142120 3000
rect 141988 1550 142108 1578
rect 142080 480 142108 1550
rect 143276 480 143304 3318
rect 144472 480 144500 3318
rect 145668 480 145696 3470
rect 146864 480 146892 3470
rect 148060 480 148088 3470
rect 150360 3330 150388 61202
rect 150440 3528 150492 3534
rect 150440 3470 150492 3476
rect 149244 3324 149296 3330
rect 149244 3266 149296 3272
rect 150348 3324 150400 3330
rect 150348 3266 150400 3272
rect 149256 480 149284 3266
rect 150452 480 150480 3470
rect 150636 3398 150664 64110
rect 151924 62082 151952 64110
rect 151912 62076 151964 62082
rect 151912 62018 151964 62024
rect 153108 62076 153160 62082
rect 153108 62018 153160 62024
rect 151636 61532 151688 61538
rect 151636 61474 151688 61480
rect 151648 3482 151676 61474
rect 151728 60988 151780 60994
rect 151728 60930 151780 60936
rect 151740 3534 151768 60930
rect 151556 3454 151676 3482
rect 151728 3528 151780 3534
rect 153120 3482 153148 62018
rect 153304 61810 153332 64110
rect 153948 64110 154284 64138
rect 154960 64110 155296 64138
rect 155972 64110 156308 64138
rect 157320 64110 157380 64138
rect 153948 61946 153976 64110
rect 153936 61940 153988 61946
rect 153936 61882 153988 61888
rect 153292 61804 153344 61810
rect 153292 61746 153344 61752
rect 154488 61804 154540 61810
rect 154488 61746 154540 61752
rect 154500 3534 154528 61746
rect 154960 61606 154988 64110
rect 155972 61742 156000 64110
rect 155960 61736 156012 61742
rect 155960 61678 156012 61684
rect 154948 61600 155000 61606
rect 154948 61542 155000 61548
rect 155868 61600 155920 61606
rect 155868 61542 155920 61548
rect 155880 3534 155908 61542
rect 157352 61470 157380 64110
rect 157996 64110 158332 64138
rect 159008 64110 159344 64138
rect 160112 64110 160356 64138
rect 161032 64110 161368 64138
rect 162136 64110 162472 64138
rect 163148 64110 163484 64138
rect 164252 64110 164496 64138
rect 165172 64110 165508 64138
rect 166184 64110 166520 64138
rect 167196 64110 167532 64138
rect 168392 64110 168544 64138
rect 169220 64110 169556 64138
rect 170232 64110 170568 64138
rect 171336 64110 171580 64138
rect 172592 64110 172652 64138
rect 157340 61464 157392 61470
rect 157340 61406 157392 61412
rect 157996 61198 158024 64110
rect 158628 61940 158680 61946
rect 158628 61882 158680 61888
rect 157984 61192 158036 61198
rect 157984 61134 158036 61140
rect 157248 60852 157300 60858
rect 157248 60794 157300 60800
rect 157260 3534 157288 60794
rect 151728 3470 151780 3476
rect 152752 3454 153148 3482
rect 153936 3528 153988 3534
rect 153936 3470 153988 3476
rect 154488 3528 154540 3534
rect 154488 3470 154540 3476
rect 155132 3528 155184 3534
rect 155132 3470 155184 3476
rect 155868 3528 155920 3534
rect 155868 3470 155920 3476
rect 156328 3528 156380 3534
rect 156328 3470 156380 3476
rect 157248 3528 157300 3534
rect 157248 3470 157300 3476
rect 150624 3392 150676 3398
rect 150624 3334 150676 3340
rect 151556 480 151584 3454
rect 152752 480 152780 3454
rect 153948 480 153976 3470
rect 155144 480 155172 3470
rect 156340 480 156368 3470
rect 158640 3330 158668 61882
rect 159008 61062 159036 64110
rect 159916 61736 159968 61742
rect 159916 61678 159968 61684
rect 158996 61056 159048 61062
rect 158996 60998 159048 61004
rect 159928 3602 159956 61678
rect 160112 61674 160140 64110
rect 160100 61668 160152 61674
rect 160100 61610 160152 61616
rect 160008 61464 160060 61470
rect 160008 61406 160060 61412
rect 158720 3596 158772 3602
rect 158720 3538 158772 3544
rect 159916 3596 159968 3602
rect 159916 3538 159968 3544
rect 157524 3324 157576 3330
rect 157524 3266 157576 3272
rect 158628 3324 158680 3330
rect 158628 3266 158680 3272
rect 157536 480 157564 3266
rect 158732 480 158760 3538
rect 160020 3482 160048 61406
rect 161032 61402 161060 64110
rect 161020 61396 161072 61402
rect 161020 61338 161072 61344
rect 161388 61192 161440 61198
rect 161388 61134 161440 61140
rect 161400 3482 161428 61134
rect 162136 61130 162164 64110
rect 163148 61878 163176 64110
rect 164252 62014 164280 64110
rect 164240 62008 164292 62014
rect 164240 61950 164292 61956
rect 163136 61872 163188 61878
rect 163136 61814 163188 61820
rect 164148 61668 164200 61674
rect 164148 61610 164200 61616
rect 162768 61396 162820 61402
rect 162768 61338 162820 61344
rect 162124 61124 162176 61130
rect 162124 61066 162176 61072
rect 162780 3534 162808 61338
rect 164160 3534 164188 61610
rect 165172 60926 165200 64110
rect 165528 61872 165580 61878
rect 165528 61814 165580 61820
rect 165160 60920 165212 60926
rect 165160 60862 165212 60868
rect 159928 3454 160048 3482
rect 161124 3454 161428 3482
rect 162308 3528 162360 3534
rect 162308 3470 162360 3476
rect 162768 3528 162820 3534
rect 162768 3470 162820 3476
rect 163504 3528 163556 3534
rect 163504 3470 163556 3476
rect 164148 3528 164200 3534
rect 164148 3470 164200 3476
rect 159928 480 159956 3454
rect 161124 480 161152 3454
rect 162320 480 162348 3470
rect 163516 480 163544 3470
rect 165540 3466 165568 61814
rect 166184 61334 166212 64110
rect 166172 61328 166224 61334
rect 166172 61270 166224 61276
rect 167196 61266 167224 64110
rect 168288 62008 168340 62014
rect 168288 61950 168340 61956
rect 168196 61328 168248 61334
rect 168196 61270 168248 61276
rect 167184 61260 167236 61266
rect 167184 61202 167236 61208
rect 166908 61124 166960 61130
rect 166908 61066 166960 61072
rect 166920 3534 166948 61066
rect 168208 3602 168236 61270
rect 167092 3596 167144 3602
rect 167092 3538 167144 3544
rect 168196 3596 168248 3602
rect 168196 3538 168248 3544
rect 165896 3528 165948 3534
rect 165896 3470 165948 3476
rect 166908 3528 166960 3534
rect 166908 3470 166960 3476
rect 164700 3460 164752 3466
rect 164700 3402 164752 3408
rect 165528 3460 165580 3466
rect 165528 3402 165580 3408
rect 164712 480 164740 3402
rect 165908 480 165936 3470
rect 167104 480 167132 3538
rect 168300 3482 168328 61950
rect 168392 60994 168420 64110
rect 169220 61538 169248 64110
rect 170232 62082 170260 64110
rect 170220 62076 170272 62082
rect 170220 62018 170272 62024
rect 171048 62076 171100 62082
rect 171048 62018 171100 62024
rect 169208 61532 169260 61538
rect 169208 61474 169260 61480
rect 169668 61532 169720 61538
rect 169668 61474 169720 61480
rect 168380 60988 168432 60994
rect 168380 60930 168432 60936
rect 169680 3482 169708 61474
rect 168208 3454 168328 3482
rect 169404 3454 169708 3482
rect 168208 480 168236 3454
rect 169404 480 169432 3454
rect 171060 3398 171088 62018
rect 171336 61810 171364 64110
rect 171324 61804 171376 61810
rect 171324 61746 171376 61752
rect 172624 61606 172652 64110
rect 173360 64110 173696 64138
rect 174372 64110 174708 64138
rect 175384 64110 175720 64138
rect 176732 64110 176792 64138
rect 172612 61600 172664 61606
rect 172612 61542 172664 61548
rect 172428 61260 172480 61266
rect 172428 61202 172480 61208
rect 172440 3534 172468 61202
rect 173360 60858 173388 64110
rect 174372 61946 174400 64110
rect 174360 61940 174412 61946
rect 174360 61882 174412 61888
rect 175188 61940 175240 61946
rect 175188 61882 175240 61888
rect 173808 61804 173860 61810
rect 173808 61746 173860 61752
rect 173348 60852 173400 60858
rect 173348 60794 173400 60800
rect 173820 3534 173848 61746
rect 171784 3528 171836 3534
rect 171784 3470 171836 3476
rect 172428 3528 172480 3534
rect 172428 3470 172480 3476
rect 172980 3528 173032 3534
rect 172980 3470 173032 3476
rect 173808 3528 173860 3534
rect 173808 3470 173860 3476
rect 170588 3392 170640 3398
rect 170588 3334 170640 3340
rect 171048 3392 171100 3398
rect 171048 3334 171100 3340
rect 170600 480 170628 3334
rect 171796 480 171824 3470
rect 172992 480 173020 3470
rect 175200 3330 175228 61882
rect 175384 61742 175412 64110
rect 175372 61736 175424 61742
rect 175372 61678 175424 61684
rect 176476 61736 176528 61742
rect 176476 61678 176528 61684
rect 174176 3324 174228 3330
rect 174176 3266 174228 3272
rect 175188 3324 175240 3330
rect 175188 3266 175240 3272
rect 174188 480 174216 3266
rect 176488 3058 176516 61678
rect 176568 61600 176620 61606
rect 176568 61542 176620 61548
rect 175372 3052 175424 3058
rect 175372 2994 175424 3000
rect 176476 3052 176528 3058
rect 176476 2994 176528 3000
rect 175384 480 175412 2994
rect 176580 480 176608 61542
rect 176764 61470 176792 64110
rect 177408 64110 177744 64138
rect 178420 64110 178756 64138
rect 179432 64110 179768 64138
rect 180780 64110 180840 64138
rect 176752 61464 176804 61470
rect 176752 61406 176804 61412
rect 177408 61198 177436 64110
rect 177948 61464 178000 61470
rect 177948 61406 178000 61412
rect 177396 61192 177448 61198
rect 177396 61134 177448 61140
rect 177960 3482 177988 61406
rect 178420 61402 178448 64110
rect 179432 61674 179460 64110
rect 180812 61878 180840 64110
rect 181456 64110 181792 64138
rect 182468 64110 182804 64138
rect 183572 64110 183816 64138
rect 184920 64110 184980 64138
rect 180800 61872 180852 61878
rect 180800 61814 180852 61820
rect 179420 61668 179472 61674
rect 179420 61610 179472 61616
rect 178408 61396 178460 61402
rect 178408 61338 178460 61344
rect 180708 61396 180760 61402
rect 180708 61338 180760 61344
rect 179328 61192 179380 61198
rect 179328 61134 179380 61140
rect 179340 3482 179368 61134
rect 180720 3534 180748 61338
rect 181456 61130 181484 64110
rect 182088 61668 182140 61674
rect 182088 61610 182140 61616
rect 181444 61124 181496 61130
rect 181444 61066 181496 61072
rect 177776 3454 177988 3482
rect 178972 3454 179368 3482
rect 180156 3528 180208 3534
rect 180156 3470 180208 3476
rect 180708 3528 180760 3534
rect 180708 3470 180760 3476
rect 177776 480 177804 3454
rect 178972 480 179000 3454
rect 180168 480 180196 3470
rect 182100 3126 182128 61610
rect 182468 61334 182496 64110
rect 183572 62014 183600 64110
rect 183560 62008 183612 62014
rect 183560 61950 183612 61956
rect 184848 61872 184900 61878
rect 184848 61814 184900 61820
rect 182456 61328 182508 61334
rect 182456 61270 182508 61276
rect 183468 61328 183520 61334
rect 183468 61270 183520 61276
rect 183480 3534 183508 61270
rect 184756 61124 184808 61130
rect 184756 61066 184808 61072
rect 184768 3534 184796 61066
rect 182548 3528 182600 3534
rect 182548 3470 182600 3476
rect 183468 3528 183520 3534
rect 183468 3470 183520 3476
rect 183744 3528 183796 3534
rect 183744 3470 183796 3476
rect 184756 3528 184808 3534
rect 184756 3470 184808 3476
rect 181352 3120 181404 3126
rect 181352 3062 181404 3068
rect 182088 3120 182140 3126
rect 182088 3062 182140 3068
rect 181364 480 181392 3062
rect 182560 480 182588 3470
rect 183756 480 183784 3470
rect 184860 480 184888 61814
rect 184952 61538 184980 64110
rect 185596 64110 185932 64138
rect 186608 64110 186944 64138
rect 187712 64110 187956 64138
rect 188632 64110 188968 64138
rect 189644 64110 189980 64138
rect 190748 64110 190992 64138
rect 191852 64110 192004 64138
rect 192680 64110 193016 64138
rect 193692 64110 194028 64138
rect 194704 64110 195040 64138
rect 195992 64110 196144 64138
rect 196820 64110 197156 64138
rect 197832 64110 198168 64138
rect 198844 64110 199180 64138
rect 200192 64110 200252 64138
rect 185596 62082 185624 64110
rect 185584 62076 185636 62082
rect 185584 62018 185636 62024
rect 186228 62008 186280 62014
rect 186228 61950 186280 61956
rect 184940 61532 184992 61538
rect 184940 61474 184992 61480
rect 186240 3482 186268 61950
rect 186608 61266 186636 64110
rect 187712 61810 187740 64110
rect 188632 61946 188660 64110
rect 188620 61940 188672 61946
rect 188620 61882 188672 61888
rect 187700 61804 187752 61810
rect 187700 61746 187752 61752
rect 188988 61804 189040 61810
rect 188988 61746 189040 61752
rect 187608 61532 187660 61538
rect 187608 61474 187660 61480
rect 186596 61260 186648 61266
rect 186596 61202 186648 61208
rect 187620 3482 187648 61474
rect 189000 3534 189028 61746
rect 189644 61742 189672 64110
rect 189632 61736 189684 61742
rect 189632 61678 189684 61684
rect 190368 61736 190420 61742
rect 190368 61678 190420 61684
rect 190380 3534 190408 61678
rect 190748 61606 190776 64110
rect 190736 61600 190788 61606
rect 190736 61542 190788 61548
rect 191748 61600 191800 61606
rect 191748 61542 191800 61548
rect 186056 3454 186268 3482
rect 187252 3454 187648 3482
rect 188436 3528 188488 3534
rect 188436 3470 188488 3476
rect 188988 3528 189040 3534
rect 188988 3470 189040 3476
rect 189632 3528 189684 3534
rect 189632 3470 189684 3476
rect 190368 3528 190420 3534
rect 190368 3470 190420 3476
rect 186056 480 186084 3454
rect 187252 480 187280 3454
rect 188448 480 188476 3470
rect 189644 480 189672 3470
rect 191760 3058 191788 61542
rect 191852 61470 191880 64110
rect 191840 61464 191892 61470
rect 191840 61406 191892 61412
rect 192680 61198 192708 64110
rect 193128 61464 193180 61470
rect 193128 61406 193180 61412
rect 192668 61192 192720 61198
rect 192668 61134 192720 61140
rect 193140 3534 193168 61406
rect 193692 61402 193720 64110
rect 194704 61674 194732 64110
rect 194692 61668 194744 61674
rect 194692 61610 194744 61616
rect 195888 61668 195940 61674
rect 195888 61610 195940 61616
rect 193680 61396 193732 61402
rect 193680 61338 193732 61344
rect 194416 61396 194468 61402
rect 194416 61338 194468 61344
rect 192024 3528 192076 3534
rect 192024 3470 192076 3476
rect 193128 3528 193180 3534
rect 193128 3470 193180 3476
rect 193220 3528 193272 3534
rect 193220 3470 193272 3476
rect 190828 3052 190880 3058
rect 190828 2994 190880 3000
rect 191748 3052 191800 3058
rect 191748 2994 191800 3000
rect 190840 480 190868 2994
rect 192036 480 192064 3470
rect 193232 480 193260 3470
rect 194428 480 194456 61338
rect 194508 61260 194560 61266
rect 194508 61202 194560 61208
rect 194520 3534 194548 61202
rect 194508 3528 194560 3534
rect 195900 3482 195928 61610
rect 195992 61334 196020 64110
rect 195980 61328 196032 61334
rect 195980 61270 196032 61276
rect 196820 61130 196848 64110
rect 197268 61940 197320 61946
rect 197268 61882 197320 61888
rect 196808 61124 196860 61130
rect 196808 61066 196860 61072
rect 197280 3534 197308 61882
rect 197832 61878 197860 64110
rect 198648 62076 198700 62082
rect 198648 62018 198700 62024
rect 197820 61872 197872 61878
rect 197820 61814 197872 61820
rect 198660 3534 198688 62018
rect 198844 62014 198872 64110
rect 198832 62008 198884 62014
rect 198832 61950 198884 61956
rect 200028 61872 200080 61878
rect 200028 61814 200080 61820
rect 200040 3534 200068 61814
rect 200224 61538 200252 64110
rect 200868 64110 201204 64138
rect 201880 64110 202216 64138
rect 202892 64110 203228 64138
rect 204240 64110 204300 64138
rect 200868 61810 200896 64110
rect 200856 61804 200908 61810
rect 200856 61746 200908 61752
rect 201408 61804 201460 61810
rect 201408 61746 201460 61752
rect 200212 61532 200264 61538
rect 200212 61474 200264 61480
rect 201420 3534 201448 61746
rect 201880 61742 201908 64110
rect 202696 62008 202748 62014
rect 202696 61950 202748 61956
rect 201868 61736 201920 61742
rect 201868 61678 201920 61684
rect 202708 3602 202736 61950
rect 202892 61606 202920 64110
rect 202880 61600 202932 61606
rect 202880 61542 202932 61548
rect 204168 61600 204220 61606
rect 204168 61542 204220 61548
rect 202788 61532 202840 61538
rect 202788 61474 202840 61480
rect 201500 3596 201552 3602
rect 201500 3538 201552 3544
rect 202696 3596 202748 3602
rect 202696 3538 202748 3544
rect 194508 3470 194560 3476
rect 195624 3454 195928 3482
rect 196808 3528 196860 3534
rect 196808 3470 196860 3476
rect 197268 3528 197320 3534
rect 197268 3470 197320 3476
rect 198004 3528 198056 3534
rect 198004 3470 198056 3476
rect 198648 3528 198700 3534
rect 198648 3470 198700 3476
rect 199200 3528 199252 3534
rect 199200 3470 199252 3476
rect 200028 3528 200080 3534
rect 200028 3470 200080 3476
rect 200396 3528 200448 3534
rect 200396 3470 200448 3476
rect 201408 3528 201460 3534
rect 201408 3470 201460 3476
rect 195624 480 195652 3454
rect 196820 480 196848 3470
rect 198016 480 198044 3470
rect 199212 480 199240 3470
rect 200408 480 200436 3470
rect 201512 480 201540 3538
rect 202800 3482 202828 61474
rect 204180 3482 204208 61542
rect 204272 61470 204300 64110
rect 204916 64110 205252 64138
rect 205928 64110 206264 64138
rect 207032 64110 207368 64138
rect 208380 64110 208440 64138
rect 204260 61464 204312 61470
rect 204260 61406 204312 61412
rect 204916 61266 204944 64110
rect 205548 61464 205600 61470
rect 205548 61406 205600 61412
rect 204904 61260 204956 61266
rect 204904 61202 204956 61208
rect 205560 3534 205588 61406
rect 205928 61402 205956 64110
rect 207032 61674 207060 64110
rect 208412 61946 208440 64110
rect 209056 64110 209392 64138
rect 210068 64110 210404 64138
rect 211172 64110 211416 64138
rect 212092 64110 212428 64138
rect 213104 64110 213440 64138
rect 214116 64110 214452 64138
rect 215312 64110 215464 64138
rect 216140 64110 216476 64138
rect 217152 64110 217488 64138
rect 218256 64110 218592 64138
rect 219452 64110 219604 64138
rect 220280 64110 220616 64138
rect 221292 64110 221628 64138
rect 222304 64110 222640 64138
rect 223652 64110 223712 64138
rect 209056 62082 209084 64110
rect 209044 62076 209096 62082
rect 209044 62018 209096 62024
rect 208400 61940 208452 61946
rect 208400 61882 208452 61888
rect 209688 61940 209740 61946
rect 209688 61882 209740 61888
rect 207020 61668 207072 61674
rect 207020 61610 207072 61616
rect 208308 61668 208360 61674
rect 208308 61610 208360 61616
rect 205916 61396 205968 61402
rect 205916 61338 205968 61344
rect 206928 61328 206980 61334
rect 206928 61270 206980 61276
rect 202708 3454 202828 3482
rect 203904 3454 204208 3482
rect 205088 3528 205140 3534
rect 205088 3470 205140 3476
rect 205548 3528 205600 3534
rect 205548 3470 205600 3476
rect 202708 480 202736 3454
rect 203904 480 203932 3454
rect 205100 480 205128 3470
rect 206940 3058 206968 61270
rect 208320 3534 208348 61610
rect 209700 3534 209728 61882
rect 210068 61878 210096 64110
rect 210056 61872 210108 61878
rect 210056 61814 210108 61820
rect 211172 61810 211200 64110
rect 212092 62014 212120 64110
rect 212080 62008 212132 62014
rect 212080 61950 212132 61956
rect 211160 61804 211212 61810
rect 211160 61746 211212 61752
rect 212448 61804 212500 61810
rect 212448 61746 212500 61752
rect 211068 61736 211120 61742
rect 211068 61678 211120 61684
rect 210976 61396 211028 61402
rect 210976 61338 211028 61344
rect 207480 3528 207532 3534
rect 207480 3470 207532 3476
rect 208308 3528 208360 3534
rect 208308 3470 208360 3476
rect 208676 3528 208728 3534
rect 208676 3470 208728 3476
rect 209688 3528 209740 3534
rect 209688 3470 209740 3476
rect 209872 3528 209924 3534
rect 209872 3470 209924 3476
rect 206284 3052 206336 3058
rect 206284 2994 206336 3000
rect 206928 3052 206980 3058
rect 206928 2994 206980 3000
rect 206296 480 206324 2994
rect 207492 480 207520 3470
rect 208688 480 208716 3470
rect 209884 480 209912 3470
rect 210988 1578 211016 61338
rect 211080 3534 211108 61678
rect 211068 3528 211120 3534
rect 212460 3482 212488 61746
rect 213104 61538 213132 64110
rect 214116 61606 214144 64110
rect 214104 61600 214156 61606
rect 214104 61542 214156 61548
rect 215208 61600 215260 61606
rect 215208 61542 215260 61548
rect 213092 61532 213144 61538
rect 213092 61474 213144 61480
rect 213828 61532 213880 61538
rect 213828 61474 213880 61480
rect 213840 3482 213868 61474
rect 215220 3534 215248 61542
rect 215312 61470 215340 64110
rect 215300 61464 215352 61470
rect 215300 61406 215352 61412
rect 216140 61334 216168 64110
rect 216588 62008 216640 62014
rect 216588 61950 216640 61956
rect 216128 61328 216180 61334
rect 216128 61270 216180 61276
rect 216600 3534 216628 61950
rect 217152 61674 217180 64110
rect 218256 61946 218284 64110
rect 218244 61940 218296 61946
rect 218244 61882 218296 61888
rect 217968 61872 218020 61878
rect 217968 61814 218020 61820
rect 217140 61668 217192 61674
rect 217140 61610 217192 61616
rect 217980 3534 218008 61814
rect 219452 61742 219480 64110
rect 219440 61736 219492 61742
rect 219440 61678 219492 61684
rect 219256 61668 219308 61674
rect 219256 61610 219308 61616
rect 219268 3534 219296 61610
rect 219348 61464 219400 61470
rect 219348 61406 219400 61412
rect 211068 3470 211120 3476
rect 212276 3454 212488 3482
rect 213472 3454 213868 3482
rect 214656 3528 214708 3534
rect 214656 3470 214708 3476
rect 215208 3528 215260 3534
rect 215208 3470 215260 3476
rect 215852 3528 215904 3534
rect 215852 3470 215904 3476
rect 216588 3528 216640 3534
rect 216588 3470 216640 3476
rect 217048 3528 217100 3534
rect 217048 3470 217100 3476
rect 217968 3528 218020 3534
rect 217968 3470 218020 3476
rect 218152 3528 218204 3534
rect 218152 3470 218204 3476
rect 219256 3528 219308 3534
rect 219256 3470 219308 3476
rect 210988 1550 211108 1578
rect 211080 480 211108 1550
rect 212276 480 212304 3454
rect 213472 480 213500 3454
rect 214668 480 214696 3470
rect 215864 480 215892 3470
rect 217060 480 217088 3470
rect 218164 480 218192 3470
rect 219360 480 219388 61406
rect 220280 61402 220308 64110
rect 221292 61810 221320 64110
rect 221280 61804 221332 61810
rect 221280 61746 221332 61752
rect 222108 61804 222160 61810
rect 222108 61746 222160 61752
rect 220268 61396 220320 61402
rect 220268 61338 220320 61344
rect 220728 60784 220780 60790
rect 220728 60726 220780 60732
rect 220740 3482 220768 60726
rect 222120 3482 222148 61746
rect 222304 61538 222332 64110
rect 223684 61606 223712 64110
rect 224328 64110 224664 64138
rect 225340 64110 225676 64138
rect 226352 64110 226688 64138
rect 227700 64110 227760 64138
rect 224328 62014 224356 64110
rect 224316 62008 224368 62014
rect 224316 61950 224368 61956
rect 225340 61878 225368 64110
rect 225328 61872 225380 61878
rect 225328 61814 225380 61820
rect 226248 61872 226300 61878
rect 226248 61814 226300 61820
rect 223672 61600 223724 61606
rect 223672 61542 223724 61548
rect 222292 61532 222344 61538
rect 222292 61474 222344 61480
rect 224868 61532 224920 61538
rect 224868 61474 224920 61480
rect 223488 61056 223540 61062
rect 223488 60998 223540 61004
rect 223500 3534 223528 60998
rect 224880 3534 224908 61474
rect 226260 3534 226288 61814
rect 226352 61674 226380 64110
rect 226340 61668 226392 61674
rect 226340 61610 226392 61616
rect 227628 61668 227680 61674
rect 227628 61610 227680 61616
rect 227640 3534 227668 61610
rect 227732 61470 227760 64110
rect 228376 64110 228712 64138
rect 229480 64110 229816 64138
rect 230492 64110 230828 64138
rect 231840 64110 231900 64138
rect 227720 61464 227772 61470
rect 227720 61406 227772 61412
rect 228376 60790 228404 64110
rect 229008 61940 229060 61946
rect 229008 61882 229060 61888
rect 228916 61464 228968 61470
rect 228916 61406 228968 61412
rect 228364 60784 228416 60790
rect 228364 60726 228416 60732
rect 228928 3602 228956 61406
rect 227720 3596 227772 3602
rect 227720 3538 227772 3544
rect 228916 3596 228968 3602
rect 228916 3538 228968 3544
rect 220556 3454 220768 3482
rect 221752 3454 222148 3482
rect 222936 3528 222988 3534
rect 222936 3470 222988 3476
rect 223488 3528 223540 3534
rect 223488 3470 223540 3476
rect 224132 3528 224184 3534
rect 224132 3470 224184 3476
rect 224868 3528 224920 3534
rect 224868 3470 224920 3476
rect 225328 3528 225380 3534
rect 225328 3470 225380 3476
rect 226248 3528 226300 3534
rect 226248 3470 226300 3476
rect 226524 3528 226576 3534
rect 226524 3470 226576 3476
rect 227628 3528 227680 3534
rect 227628 3470 227680 3476
rect 220556 480 220584 3454
rect 221752 480 221780 3454
rect 222948 480 222976 3470
rect 224144 480 224172 3470
rect 225340 480 225368 3470
rect 226536 480 226564 3470
rect 227732 480 227760 3538
rect 229020 3482 229048 61882
rect 229480 61810 229508 64110
rect 229468 61804 229520 61810
rect 229468 61746 229520 61752
rect 230492 61062 230520 64110
rect 231872 61538 231900 64110
rect 232516 64110 232852 64138
rect 233528 64110 233864 64138
rect 234632 64110 234876 64138
rect 235552 64110 235888 64138
rect 236564 64110 236900 64138
rect 237576 64110 237912 64138
rect 238772 64110 238924 64138
rect 239692 64110 240028 64138
rect 240704 64110 241040 64138
rect 241716 64110 242052 64138
rect 242912 64110 243064 64138
rect 243740 64110 244076 64138
rect 244752 64110 245088 64138
rect 245764 64110 246100 64138
rect 247112 64110 247172 64138
rect 232516 61878 232544 64110
rect 232504 61872 232556 61878
rect 232504 61814 232556 61820
rect 233528 61674 233556 64110
rect 233516 61668 233568 61674
rect 233516 61610 233568 61616
rect 231860 61532 231912 61538
rect 231860 61474 231912 61480
rect 234632 61470 234660 64110
rect 235552 61946 235580 64110
rect 235540 61940 235592 61946
rect 235540 61882 235592 61888
rect 234620 61464 234672 61470
rect 234620 61406 234672 61412
rect 233148 61124 233200 61130
rect 233148 61066 233200 61072
rect 230480 61056 230532 61062
rect 230480 60998 230532 61004
rect 231768 60852 231820 60858
rect 231768 60794 231820 60800
rect 230388 60784 230440 60790
rect 230388 60726 230440 60732
rect 230400 3482 230428 60726
rect 231780 3534 231808 60794
rect 233160 3534 233188 61066
rect 234528 61056 234580 61062
rect 234528 60998 234580 61004
rect 234540 3534 234568 60998
rect 235908 60988 235960 60994
rect 235908 60930 235960 60936
rect 228928 3454 229048 3482
rect 230124 3454 230428 3482
rect 231308 3528 231360 3534
rect 231308 3470 231360 3476
rect 231768 3528 231820 3534
rect 231768 3470 231820 3476
rect 232504 3528 232556 3534
rect 232504 3470 232556 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 233700 3528 233752 3534
rect 233700 3470 233752 3476
rect 234528 3528 234580 3534
rect 234528 3470 234580 3476
rect 228928 480 228956 3454
rect 230124 480 230152 3454
rect 231320 480 231348 3470
rect 232516 480 232544 3470
rect 233712 480 233740 3470
rect 235920 3330 235948 60930
rect 236564 60790 236592 64110
rect 237288 61464 237340 61470
rect 237288 61406 237340 61412
rect 237196 61396 237248 61402
rect 237196 61338 237248 61344
rect 236552 60784 236604 60790
rect 236552 60726 236604 60732
rect 234804 3324 234856 3330
rect 234804 3266 234856 3272
rect 235908 3324 235960 3330
rect 235908 3266 235960 3272
rect 234816 480 234844 3266
rect 236000 3256 236052 3262
rect 236000 3198 236052 3204
rect 236012 480 236040 3198
rect 237208 480 237236 61338
rect 237300 3262 237328 61406
rect 237576 60858 237604 64110
rect 238668 61600 238720 61606
rect 238668 61542 238720 61548
rect 237564 60852 237616 60858
rect 237564 60794 237616 60800
rect 238680 3482 238708 61542
rect 238772 61130 238800 64110
rect 238760 61124 238812 61130
rect 238760 61066 238812 61072
rect 239692 61062 239720 64110
rect 239680 61056 239732 61062
rect 239680 60998 239732 61004
rect 240704 60994 240732 64110
rect 241716 61470 241744 64110
rect 241704 61464 241756 61470
rect 241704 61406 241756 61412
rect 242912 61402 242940 64110
rect 243740 61606 243768 64110
rect 243728 61600 243780 61606
rect 243728 61542 243780 61548
rect 242900 61396 242952 61402
rect 242900 61338 242952 61344
rect 241428 61056 241480 61062
rect 241428 60998 241480 61004
rect 240692 60988 240744 60994
rect 240692 60930 240744 60936
rect 240048 60852 240100 60858
rect 240048 60794 240100 60800
rect 240060 3534 240088 60794
rect 241440 3534 241468 60998
rect 242808 60920 242860 60926
rect 242808 60862 242860 60868
rect 238404 3454 238708 3482
rect 239588 3528 239640 3534
rect 239588 3470 239640 3476
rect 240048 3528 240100 3534
rect 240048 3470 240100 3476
rect 240784 3528 240836 3534
rect 240784 3470 240836 3476
rect 241428 3528 241480 3534
rect 241428 3470 241480 3476
rect 237288 3256 237340 3262
rect 237288 3198 237340 3204
rect 238404 480 238432 3454
rect 239600 480 239628 3470
rect 240796 480 240824 3470
rect 242820 3466 242848 60862
rect 244752 60858 244780 64110
rect 245476 61124 245528 61130
rect 245476 61066 245528 61072
rect 244740 60852 244792 60858
rect 244740 60794 244792 60800
rect 244188 60784 244240 60790
rect 244188 60726 244240 60732
rect 244200 3534 244228 60726
rect 244372 3596 244424 3602
rect 244372 3538 244424 3544
rect 243176 3528 243228 3534
rect 243176 3470 243228 3476
rect 244188 3528 244240 3534
rect 244188 3470 244240 3476
rect 241980 3460 242032 3466
rect 241980 3402 242032 3408
rect 242808 3460 242860 3466
rect 242808 3402 242860 3408
rect 241992 480 242020 3402
rect 243188 480 243216 3470
rect 244384 480 244412 3538
rect 245488 3482 245516 61066
rect 245764 61062 245792 64110
rect 246948 61532 247000 61538
rect 246948 61474 247000 61480
rect 245752 61056 245804 61062
rect 245752 60998 245804 61004
rect 245568 60988 245620 60994
rect 245568 60930 245620 60936
rect 245580 3602 245608 60930
rect 245568 3596 245620 3602
rect 245568 3538 245620 3544
rect 246960 3482 246988 61474
rect 247144 60926 247172 64110
rect 247788 64110 248124 64138
rect 248800 64110 249136 64138
rect 249812 64110 250148 64138
rect 251252 64110 251312 64138
rect 247132 60920 247184 60926
rect 247132 60862 247184 60868
rect 247788 60790 247816 64110
rect 248800 60994 248828 64110
rect 249812 61130 249840 64110
rect 251284 61538 251312 64110
rect 251928 64110 252264 64138
rect 252940 64110 253276 64138
rect 253952 64110 254288 64138
rect 255300 64110 255360 64138
rect 251272 61532 251324 61538
rect 251272 61474 251324 61480
rect 249800 61124 249852 61130
rect 249800 61066 249852 61072
rect 248788 60988 248840 60994
rect 248788 60930 248840 60936
rect 251088 60988 251140 60994
rect 251088 60930 251140 60936
rect 249708 60920 249760 60926
rect 249708 60862 249760 60868
rect 247776 60784 247828 60790
rect 247776 60726 247828 60732
rect 249064 60784 249116 60790
rect 249064 60726 249116 60732
rect 245488 3454 245608 3482
rect 245580 480 245608 3454
rect 246776 3454 246988 3482
rect 246776 480 246804 3454
rect 249076 3398 249104 60726
rect 249720 3534 249748 60862
rect 249156 3528 249208 3534
rect 249156 3470 249208 3476
rect 249708 3528 249760 3534
rect 249708 3470 249760 3476
rect 247960 3392 248012 3398
rect 247960 3334 248012 3340
rect 249064 3392 249116 3398
rect 249064 3334 249116 3340
rect 247972 480 248000 3334
rect 249168 480 249196 3470
rect 251100 3466 251128 60930
rect 251928 60790 251956 64110
rect 252940 60926 252968 64110
rect 253952 60994 253980 64110
rect 253940 60988 253992 60994
rect 253940 60930 253992 60936
rect 255228 60988 255280 60994
rect 255228 60930 255280 60936
rect 252928 60920 252980 60926
rect 252928 60862 252980 60868
rect 253756 60920 253808 60926
rect 253756 60862 253808 60868
rect 252468 60852 252520 60858
rect 252468 60794 252520 60800
rect 251916 60784 251968 60790
rect 251916 60726 251968 60732
rect 252480 3534 252508 60794
rect 252652 3596 252704 3602
rect 252652 3538 252704 3544
rect 251456 3528 251508 3534
rect 251456 3470 251508 3476
rect 252468 3528 252520 3534
rect 252468 3470 252520 3476
rect 250352 3460 250404 3466
rect 250352 3402 250404 3408
rect 251088 3460 251140 3466
rect 251088 3402 251140 3408
rect 250364 480 250392 3402
rect 251468 480 251496 3470
rect 252664 480 252692 3538
rect 253768 3482 253796 60862
rect 253848 60784 253900 60790
rect 253848 60726 253900 60732
rect 253860 3602 253888 60726
rect 253848 3596 253900 3602
rect 253848 3538 253900 3544
rect 255240 3482 255268 60930
rect 255332 60858 255360 64110
rect 255976 64110 256312 64138
rect 256988 64110 257324 64138
rect 258184 64110 258336 64138
rect 259012 64110 259348 64138
rect 260024 64110 260360 64138
rect 261036 64110 261372 64138
rect 262232 64110 262476 64138
rect 263152 64110 263488 64138
rect 263704 64110 264500 64138
rect 265176 64110 265512 64138
rect 266372 64110 266524 64138
rect 267200 64110 267536 64138
rect 267844 64110 268548 64138
rect 269132 64110 269560 64138
rect 255320 60852 255372 60858
rect 255320 60794 255372 60800
rect 255976 60790 256004 64110
rect 256608 61124 256660 61130
rect 256608 61066 256660 61072
rect 255964 60784 256016 60790
rect 255964 60726 256016 60732
rect 256620 3482 256648 61066
rect 256988 60926 257016 64110
rect 257988 61056 258040 61062
rect 257988 60998 258040 61004
rect 256976 60920 257028 60926
rect 256976 60862 257028 60868
rect 258000 3534 258028 60998
rect 258184 60994 258212 64110
rect 259012 61130 259040 64110
rect 259000 61124 259052 61130
rect 259000 61066 259052 61072
rect 260024 61062 260052 64110
rect 260012 61056 260064 61062
rect 260012 60998 260064 61004
rect 258172 60988 258224 60994
rect 258172 60930 258224 60936
rect 260748 60852 260800 60858
rect 260748 60794 260800 60800
rect 259368 60784 259420 60790
rect 259368 60726 259420 60732
rect 259380 3534 259408 60726
rect 253768 3454 253888 3482
rect 253860 480 253888 3454
rect 255056 3454 255268 3482
rect 256252 3454 256648 3482
rect 257436 3528 257488 3534
rect 257436 3470 257488 3476
rect 257988 3528 258040 3534
rect 257988 3470 258040 3476
rect 258632 3528 258684 3534
rect 258632 3470 258684 3476
rect 259368 3528 259420 3534
rect 259368 3470 259420 3476
rect 255056 480 255084 3454
rect 256252 480 256280 3454
rect 257448 480 257476 3470
rect 258644 480 258672 3470
rect 260760 3058 260788 60794
rect 261036 60790 261064 64110
rect 262232 60858 262260 64110
rect 262220 60852 262272 60858
rect 262220 60794 262272 60800
rect 263152 60790 263180 64110
rect 261024 60784 261076 60790
rect 261024 60726 261076 60732
rect 262128 60784 262180 60790
rect 262128 60726 262180 60732
rect 263140 60784 263192 60790
rect 263140 60726 263192 60732
rect 263508 60784 263560 60790
rect 263508 60726 263560 60732
rect 262140 3058 262168 60726
rect 262220 3528 262272 3534
rect 263520 3482 263548 60726
rect 263704 3534 263732 64110
rect 264888 60852 264940 60858
rect 264888 60794 264940 60800
rect 262220 3470 262272 3476
rect 259828 3052 259880 3058
rect 259828 2994 259880 3000
rect 260748 3052 260800 3058
rect 260748 2994 260800 3000
rect 261024 3052 261076 3058
rect 261024 2994 261076 3000
rect 262128 3052 262180 3058
rect 262128 2994 262180 3000
rect 259840 480 259868 2994
rect 261036 480 261064 2994
rect 262232 480 262260 3470
rect 263428 3454 263548 3482
rect 263692 3528 263744 3534
rect 264900 3482 264928 60794
rect 265176 60790 265204 64110
rect 266372 60858 266400 64110
rect 266360 60852 266412 60858
rect 266360 60794 266412 60800
rect 267200 60790 267228 64110
rect 265164 60784 265216 60790
rect 265164 60726 265216 60732
rect 266268 60784 266320 60790
rect 266268 60726 266320 60732
rect 267188 60784 267240 60790
rect 267188 60726 267240 60732
rect 266280 3534 266308 60726
rect 263692 3470 263744 3476
rect 264624 3454 264928 3482
rect 265808 3528 265860 3534
rect 265808 3470 265860 3476
rect 266268 3528 266320 3534
rect 266268 3470 266320 3476
rect 263428 480 263456 3454
rect 264624 480 264652 3454
rect 265820 480 265848 3470
rect 267844 3262 267872 64110
rect 269132 60738 269160 64110
rect 270558 63866 270586 64124
rect 270512 63838 270586 63866
rect 270696 64110 271584 64138
rect 271892 64110 272596 64138
rect 273364 64110 273700 64138
rect 270512 60738 270540 63838
rect 269040 60710 269160 60738
rect 270420 60710 270540 60738
rect 269040 3534 269068 60710
rect 270420 3534 270448 60710
rect 268108 3528 268160 3534
rect 268108 3470 268160 3476
rect 269028 3528 269080 3534
rect 269028 3470 269080 3476
rect 269304 3528 269356 3534
rect 269304 3470 269356 3476
rect 270408 3528 270460 3534
rect 270696 3482 270724 64110
rect 271892 3482 271920 64110
rect 273364 3534 273392 64110
rect 274698 63866 274726 64124
rect 274652 63838 274726 63866
rect 274836 64110 275724 64138
rect 276032 64110 276736 64138
rect 277412 64110 277748 64138
rect 278760 64110 278820 64138
rect 274652 60738 274680 63838
rect 274560 60710 274680 60738
rect 270408 3470 270460 3476
rect 267004 3256 267056 3262
rect 267004 3198 267056 3204
rect 267832 3256 267884 3262
rect 267832 3198 267884 3204
rect 267016 480 267044 3198
rect 268120 480 268148 3470
rect 269316 480 269344 3470
rect 270512 3454 270724 3482
rect 271708 3454 271920 3482
rect 272892 3528 272944 3534
rect 272892 3470 272944 3476
rect 273352 3528 273404 3534
rect 273352 3470 273404 3476
rect 270512 480 270540 3454
rect 271708 480 271736 3454
rect 272904 480 272932 3470
rect 274560 2922 274588 60710
rect 274836 3262 274864 64110
rect 276032 3534 276060 64110
rect 276020 3528 276072 3534
rect 276020 3470 276072 3476
rect 276480 3528 276532 3534
rect 276480 3470 276532 3476
rect 277412 3482 277440 64110
rect 278792 3482 278820 64110
rect 278884 64110 279772 64138
rect 280172 64110 280784 64138
rect 281552 64110 281796 64138
rect 282808 64110 282868 64138
rect 283820 64110 284248 64138
rect 284924 64110 285628 64138
rect 285936 64110 286272 64138
rect 286948 64110 287008 64138
rect 287960 64110 288388 64138
rect 288972 64110 289308 64138
rect 289984 64110 290320 64138
rect 290996 64110 291056 64138
rect 292008 64110 292528 64138
rect 293020 64110 293356 64138
rect 294032 64110 294368 64138
rect 295044 64110 295288 64138
rect 296148 64110 296668 64138
rect 297160 64110 297496 64138
rect 298172 64110 298508 64138
rect 299184 64110 299336 64138
rect 300196 64110 300808 64138
rect 301208 64110 301544 64138
rect 302220 64110 302556 64138
rect 303232 64110 303476 64138
rect 304244 64110 304948 64138
rect 305256 64110 305592 64138
rect 278884 3602 278912 64110
rect 278872 3596 278924 3602
rect 278872 3538 278924 3544
rect 280068 3596 280120 3602
rect 280068 3538 280120 3544
rect 274824 3256 274876 3262
rect 274824 3198 274876 3204
rect 275284 3256 275336 3262
rect 275284 3198 275336 3204
rect 274088 2916 274140 2922
rect 274088 2858 274140 2864
rect 274548 2916 274600 2922
rect 274548 2858 274600 2864
rect 274100 480 274128 2858
rect 275296 480 275324 3198
rect 276492 480 276520 3470
rect 277412 3454 277716 3482
rect 278792 3454 278912 3482
rect 277688 480 277716 3454
rect 278884 480 278912 3454
rect 280080 480 280108 3538
rect 280172 3330 280200 64110
rect 281552 3534 281580 64110
rect 282840 60738 282868 64110
rect 284220 60738 284248 64110
rect 282840 60710 282960 60738
rect 284220 60710 284432 60738
rect 281540 3528 281592 3534
rect 281540 3470 281592 3476
rect 282460 3528 282512 3534
rect 282460 3470 282512 3476
rect 282932 3482 282960 60710
rect 284404 3482 284432 60710
rect 285600 3482 285628 64110
rect 286244 60790 286272 64110
rect 286980 61010 287008 64110
rect 286980 60982 287100 61010
rect 286232 60784 286284 60790
rect 286232 60726 286284 60732
rect 286968 60784 287020 60790
rect 286968 60726 287020 60732
rect 286980 4128 287008 60726
rect 287072 59106 287100 60982
rect 288360 60738 288388 64110
rect 289280 60790 289308 64110
rect 290292 60790 290320 64110
rect 289268 60784 289320 60790
rect 288360 60710 288480 60738
rect 289268 60726 289320 60732
rect 290004 60784 290056 60790
rect 290004 60726 290056 60732
rect 290280 60784 290332 60790
rect 290280 60726 290332 60732
rect 287072 59078 287284 59106
rect 286980 4100 287192 4128
rect 280160 3324 280212 3330
rect 280160 3266 280212 3272
rect 281264 3324 281316 3330
rect 281264 3266 281316 3272
rect 281276 480 281304 3266
rect 282472 480 282500 3470
rect 282932 3454 283696 3482
rect 284404 3454 284800 3482
rect 285600 3454 285996 3482
rect 283668 480 283696 3454
rect 284772 480 284800 3454
rect 285968 480 285996 3454
rect 287164 480 287192 4100
rect 287256 3482 287284 59078
rect 288452 3482 288480 60710
rect 290016 3482 290044 60726
rect 287256 3454 288388 3482
rect 288452 3454 289584 3482
rect 290016 3454 290780 3482
rect 288360 480 288388 3454
rect 289556 480 289584 3454
rect 290752 480 290780 3454
rect 291028 2990 291056 64110
rect 291108 60784 291160 60790
rect 291108 60726 291160 60732
rect 291120 3534 291148 60726
rect 292500 3534 292528 64110
rect 293328 60790 293356 64110
rect 294340 60790 294368 64110
rect 293316 60784 293368 60790
rect 293316 60726 293368 60732
rect 293868 60784 293920 60790
rect 293868 60726 293920 60732
rect 294328 60784 294380 60790
rect 294328 60726 294380 60732
rect 295156 60784 295208 60790
rect 295156 60726 295208 60732
rect 293880 3602 293908 60726
rect 295168 4078 295196 60726
rect 295156 4072 295208 4078
rect 295156 4014 295208 4020
rect 293868 3596 293920 3602
rect 293868 3538 293920 3544
rect 291108 3528 291160 3534
rect 291108 3470 291160 3476
rect 291936 3528 291988 3534
rect 291936 3470 291988 3476
rect 292488 3528 292540 3534
rect 292488 3470 292540 3476
rect 294328 3528 294380 3534
rect 294328 3470 294380 3476
rect 291016 2984 291068 2990
rect 291016 2926 291068 2932
rect 291948 480 291976 3470
rect 293132 2984 293184 2990
rect 293132 2926 293184 2932
rect 293144 480 293172 2926
rect 294340 480 294368 3470
rect 295260 3466 295288 64110
rect 296640 4146 296668 64110
rect 297468 60790 297496 64110
rect 298480 60790 298508 64110
rect 297456 60784 297508 60790
rect 297456 60726 297508 60732
rect 298008 60784 298060 60790
rect 298008 60726 298060 60732
rect 298468 60784 298520 60790
rect 298468 60726 298520 60732
rect 296628 4140 296680 4146
rect 296628 4082 296680 4088
rect 296720 4072 296772 4078
rect 296720 4014 296772 4020
rect 295524 3596 295576 3602
rect 295524 3538 295576 3544
rect 295248 3460 295300 3466
rect 295248 3402 295300 3408
rect 295536 480 295564 3538
rect 296732 480 296760 4014
rect 298020 3534 298048 60726
rect 299112 4140 299164 4146
rect 299112 4082 299164 4088
rect 298008 3528 298060 3534
rect 298008 3470 298060 3476
rect 297916 3460 297968 3466
rect 297916 3402 297968 3408
rect 297928 480 297956 3402
rect 299124 480 299152 4082
rect 299308 2990 299336 64110
rect 299388 60784 299440 60790
rect 299388 60726 299440 60732
rect 299400 3058 299428 60726
rect 300308 3528 300360 3534
rect 300308 3470 300360 3476
rect 299388 3052 299440 3058
rect 299388 2994 299440 3000
rect 299296 2984 299348 2990
rect 299296 2926 299348 2932
rect 300320 480 300348 3470
rect 300780 3466 300808 64110
rect 301516 60790 301544 64110
rect 302528 60790 302556 64110
rect 301504 60784 301556 60790
rect 301504 60726 301556 60732
rect 302148 60784 302200 60790
rect 302148 60726 302200 60732
rect 302516 60784 302568 60790
rect 302516 60726 302568 60732
rect 302160 3534 302188 60726
rect 303448 3602 303476 64110
rect 303528 60784 303580 60790
rect 303528 60726 303580 60732
rect 303436 3596 303488 3602
rect 303436 3538 303488 3544
rect 302148 3528 302200 3534
rect 302148 3470 302200 3476
rect 300768 3460 300820 3466
rect 300768 3402 300820 3408
rect 303540 3194 303568 60726
rect 304920 4146 304948 64110
rect 305564 60790 305592 64110
rect 306254 63866 306282 64124
rect 307372 64110 307708 64138
rect 308384 64110 309088 64138
rect 309396 64110 309732 64138
rect 306208 63838 306282 63866
rect 305552 60784 305604 60790
rect 305552 60726 305604 60732
rect 304908 4140 304960 4146
rect 304908 4082 304960 4088
rect 305000 3528 305052 3534
rect 305000 3470 305052 3476
rect 303804 3460 303856 3466
rect 303804 3402 303856 3408
rect 303528 3188 303580 3194
rect 303528 3130 303580 3136
rect 301412 3052 301464 3058
rect 301412 2994 301464 3000
rect 301424 480 301452 2994
rect 302608 2984 302660 2990
rect 302608 2926 302660 2932
rect 302620 480 302648 2926
rect 303816 480 303844 3402
rect 305012 480 305040 3470
rect 306208 3466 306236 63838
rect 306288 60784 306340 60790
rect 306288 60726 306340 60732
rect 306300 3738 306328 60726
rect 306288 3732 306340 3738
rect 306288 3674 306340 3680
rect 307392 3596 307444 3602
rect 307392 3538 307444 3544
rect 306196 3460 306248 3466
rect 306196 3402 306248 3408
rect 306196 3188 306248 3194
rect 306196 3130 306248 3136
rect 306208 480 306236 3130
rect 307404 480 307432 3538
rect 307680 3262 307708 64110
rect 308588 4140 308640 4146
rect 308588 4082 308640 4088
rect 307668 3256 307720 3262
rect 307668 3198 307720 3204
rect 308600 480 308628 4082
rect 309060 3534 309088 64110
rect 309704 60790 309732 64110
rect 310394 63866 310422 64124
rect 311420 64110 311848 64138
rect 312432 64110 312768 64138
rect 313444 64110 313780 64138
rect 314456 64110 314608 64138
rect 315468 64110 315988 64138
rect 316480 64110 316816 64138
rect 317492 64110 317828 64138
rect 318596 64110 318656 64138
rect 319608 64110 320128 64138
rect 320620 64110 320956 64138
rect 321632 64110 321968 64138
rect 322644 64110 322796 64138
rect 323656 64110 324268 64138
rect 324668 64110 325004 64138
rect 325680 64110 326016 64138
rect 326692 64110 327028 64138
rect 327704 64110 328408 64138
rect 328716 64110 329052 64138
rect 329820 64110 330156 64138
rect 330832 64110 331076 64138
rect 331844 64110 332548 64138
rect 332856 64110 333192 64138
rect 310348 63838 310422 63866
rect 309692 60784 309744 60790
rect 309692 60726 309744 60732
rect 309784 3732 309836 3738
rect 309784 3674 309836 3680
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 309796 480 309824 3674
rect 310348 3398 310376 63838
rect 310428 60784 310480 60790
rect 310428 60726 310480 60732
rect 310336 3392 310388 3398
rect 310336 3334 310388 3340
rect 310440 3330 310468 60726
rect 310980 3460 311032 3466
rect 310980 3402 311032 3408
rect 310428 3324 310480 3330
rect 310428 3266 310480 3272
rect 310992 480 311020 3402
rect 311820 3058 311848 64110
rect 312740 60790 312768 64110
rect 313752 60790 313780 64110
rect 312728 60784 312780 60790
rect 312728 60726 312780 60732
rect 313188 60784 313240 60790
rect 313188 60726 313240 60732
rect 313740 60784 313792 60790
rect 313740 60726 313792 60732
rect 314476 60784 314528 60790
rect 314476 60726 314528 60732
rect 313200 3874 313228 60726
rect 313188 3868 313240 3874
rect 313188 3810 313240 3816
rect 314488 3670 314516 60726
rect 314476 3664 314528 3670
rect 314476 3606 314528 3612
rect 314580 3602 314608 64110
rect 314568 3596 314620 3602
rect 314568 3538 314620 3544
rect 313372 3528 313424 3534
rect 313372 3470 313424 3476
rect 312176 3256 312228 3262
rect 312176 3198 312228 3204
rect 311808 3052 311860 3058
rect 311808 2994 311860 3000
rect 312188 480 312216 3198
rect 313384 480 313412 3470
rect 315960 3466 315988 64110
rect 316788 60790 316816 64110
rect 317800 60790 317828 64110
rect 316776 60784 316828 60790
rect 316776 60726 316828 60732
rect 317328 60784 317380 60790
rect 317328 60726 317380 60732
rect 317788 60784 317840 60790
rect 317788 60726 317840 60732
rect 317340 3534 317368 60726
rect 318064 3868 318116 3874
rect 318064 3810 318116 3816
rect 317328 3528 317380 3534
rect 317328 3470 317380 3476
rect 315948 3460 316000 3466
rect 315948 3402 316000 3408
rect 315764 3392 315816 3398
rect 315764 3334 315816 3340
rect 314568 3324 314620 3330
rect 314568 3266 314620 3272
rect 314580 480 314608 3266
rect 315776 480 315804 3334
rect 316960 3052 317012 3058
rect 316960 2994 317012 3000
rect 316972 480 317000 2994
rect 318076 480 318104 3810
rect 318628 3398 318656 64110
rect 318708 60784 318760 60790
rect 318708 60726 318760 60732
rect 318616 3392 318668 3398
rect 318616 3334 318668 3340
rect 318720 2922 318748 60726
rect 320100 4146 320128 64110
rect 320928 60790 320956 64110
rect 321940 60790 321968 64110
rect 320916 60784 320968 60790
rect 320916 60726 320968 60732
rect 321468 60784 321520 60790
rect 321468 60726 321520 60732
rect 321928 60784 321980 60790
rect 321928 60726 321980 60732
rect 320088 4140 320140 4146
rect 320088 4082 320140 4088
rect 319260 3664 319312 3670
rect 319260 3606 319312 3612
rect 318708 2916 318760 2922
rect 318708 2858 318760 2864
rect 319272 480 319300 3606
rect 320456 3596 320508 3602
rect 320456 3538 320508 3544
rect 320468 480 320496 3538
rect 321480 3058 321508 60726
rect 322768 3466 322796 64110
rect 322848 60784 322900 60790
rect 322848 60726 322900 60732
rect 322860 3670 322888 60726
rect 322848 3664 322900 3670
rect 322848 3606 322900 3612
rect 324240 3602 324268 64110
rect 324976 60790 325004 64110
rect 325988 60790 326016 64110
rect 324964 60784 325016 60790
rect 324964 60726 325016 60732
rect 325608 60784 325660 60790
rect 325608 60726 325660 60732
rect 325976 60784 326028 60790
rect 325976 60726 326028 60732
rect 326896 60784 326948 60790
rect 326896 60726 326948 60732
rect 325620 3942 325648 60726
rect 326436 4140 326488 4146
rect 326436 4082 326488 4088
rect 325608 3936 325660 3942
rect 325608 3878 325660 3884
rect 324228 3596 324280 3602
rect 324228 3538 324280 3544
rect 322848 3528 322900 3534
rect 322848 3470 322900 3476
rect 321652 3460 321704 3466
rect 321652 3402 321704 3408
rect 322756 3460 322808 3466
rect 322756 3402 322808 3408
rect 321468 3052 321520 3058
rect 321468 2994 321520 3000
rect 321664 480 321692 3402
rect 322860 480 322888 3470
rect 325240 3392 325292 3398
rect 325240 3334 325292 3340
rect 324044 2916 324096 2922
rect 324044 2858 324096 2864
rect 324056 480 324084 2858
rect 325252 480 325280 3334
rect 326448 480 326476 4082
rect 326908 3398 326936 60726
rect 326896 3392 326948 3398
rect 326896 3334 326948 3340
rect 327000 2922 327028 64110
rect 328380 3806 328408 64110
rect 329024 60790 329052 64110
rect 330128 60790 330156 64110
rect 329012 60784 329064 60790
rect 329012 60726 329064 60732
rect 329748 60784 329800 60790
rect 329748 60726 329800 60732
rect 330116 60784 330168 60790
rect 330116 60726 330168 60732
rect 328368 3800 328420 3806
rect 328368 3742 328420 3748
rect 328828 3664 328880 3670
rect 328828 3606 328880 3612
rect 327632 3052 327684 3058
rect 327632 2994 327684 3000
rect 326988 2916 327040 2922
rect 326988 2858 327040 2864
rect 327644 480 327672 2994
rect 328840 480 328868 3606
rect 329760 2990 329788 60726
rect 331048 3534 331076 64110
rect 331128 60784 331180 60790
rect 331128 60726 331180 60732
rect 331140 3670 331168 60726
rect 332520 4010 332548 64110
rect 333164 60790 333192 64110
rect 333854 63866 333882 64124
rect 334880 64110 335308 64138
rect 335892 64110 336228 64138
rect 336904 64110 337240 64138
rect 337916 64110 338068 64138
rect 338928 64110 339448 64138
rect 340032 64110 340368 64138
rect 341044 64110 341380 64138
rect 342056 64110 342208 64138
rect 343068 64110 343588 64138
rect 344080 64110 344416 64138
rect 345092 64110 345428 64138
rect 346104 64110 346256 64138
rect 347116 64110 347728 64138
rect 348128 64110 348464 64138
rect 349140 64110 349476 64138
rect 350152 64110 350488 64138
rect 351256 64110 351868 64138
rect 352268 64110 352604 64138
rect 353280 64110 353616 64138
rect 354292 64110 354536 64138
rect 355304 64110 356008 64138
rect 356316 64110 356652 64138
rect 357328 64110 357388 64138
rect 358340 64110 358768 64138
rect 359352 64110 359688 64138
rect 360364 64110 360700 64138
rect 361376 64110 361436 64138
rect 362480 64110 362908 64138
rect 363492 64110 363828 64138
rect 364504 64110 364840 64138
rect 365516 64110 365668 64138
rect 366528 64110 367048 64138
rect 367540 64110 367876 64138
rect 368552 64110 368888 64138
rect 369564 64110 369808 64138
rect 370576 64110 371188 64138
rect 371588 64110 371924 64138
rect 372600 64110 372936 64138
rect 373704 64110 373856 64138
rect 374716 64110 375328 64138
rect 375728 64110 376064 64138
rect 376740 64110 377076 64138
rect 377752 64110 378088 64138
rect 378764 64110 379468 64138
rect 379776 64110 380112 64138
rect 333808 63838 333882 63866
rect 333152 60784 333204 60790
rect 333152 60726 333204 60732
rect 332508 4004 332560 4010
rect 332508 3946 332560 3952
rect 332416 3936 332468 3942
rect 332416 3878 332468 3884
rect 331128 3664 331180 3670
rect 331128 3606 331180 3612
rect 331220 3596 331272 3602
rect 331220 3538 331272 3544
rect 331036 3528 331088 3534
rect 331036 3470 331088 3476
rect 330024 3460 330076 3466
rect 330024 3402 330076 3408
rect 329748 2984 329800 2990
rect 329748 2926 329800 2932
rect 330036 480 330064 3402
rect 331232 480 331260 3538
rect 332428 480 332456 3878
rect 333808 3602 333836 63838
rect 333888 60784 333940 60790
rect 333888 60726 333940 60732
rect 333900 3874 333928 60726
rect 335280 3942 335308 64110
rect 336200 60790 336228 64110
rect 337212 60790 337240 64110
rect 336188 60784 336240 60790
rect 336188 60726 336240 60732
rect 336648 60784 336700 60790
rect 336648 60726 336700 60732
rect 337200 60784 337252 60790
rect 337200 60726 337252 60732
rect 337936 60784 337988 60790
rect 337936 60726 337988 60732
rect 335268 3936 335320 3942
rect 335268 3878 335320 3884
rect 333888 3868 333940 3874
rect 333888 3810 333940 3816
rect 336660 3806 336688 60726
rect 335912 3800 335964 3806
rect 335912 3742 335964 3748
rect 336648 3800 336700 3806
rect 336648 3742 336700 3748
rect 333796 3596 333848 3602
rect 333796 3538 333848 3544
rect 333612 3392 333664 3398
rect 333612 3334 333664 3340
rect 333624 480 333652 3334
rect 334716 2916 334768 2922
rect 334716 2858 334768 2864
rect 334728 480 334756 2858
rect 335924 480 335952 3742
rect 337948 3738 337976 60726
rect 337936 3732 337988 3738
rect 337936 3674 337988 3680
rect 338040 3466 338068 64110
rect 339420 4146 339448 64110
rect 340340 60790 340368 64110
rect 341352 60790 341380 64110
rect 340328 60784 340380 60790
rect 340328 60726 340380 60732
rect 340788 60784 340840 60790
rect 340788 60726 340840 60732
rect 341340 60784 341392 60790
rect 341340 60726 341392 60732
rect 342076 60784 342128 60790
rect 342076 60726 342128 60732
rect 339408 4140 339460 4146
rect 339408 4082 339460 4088
rect 340800 4078 340828 60726
rect 340788 4072 340840 4078
rect 340788 4014 340840 4020
rect 342088 4010 342116 60726
rect 340696 4004 340748 4010
rect 340696 3946 340748 3952
rect 342076 4004 342128 4010
rect 342076 3946 342128 3952
rect 338304 3664 338356 3670
rect 338304 3606 338356 3612
rect 338028 3460 338080 3466
rect 338028 3402 338080 3408
rect 337108 2984 337160 2990
rect 337108 2926 337160 2932
rect 337120 480 337148 2926
rect 338316 480 338344 3606
rect 339500 3528 339552 3534
rect 339500 3470 339552 3476
rect 339512 480 339540 3470
rect 340708 480 340736 3946
rect 342180 3874 342208 64110
rect 341892 3868 341944 3874
rect 341892 3810 341944 3816
rect 342168 3868 342220 3874
rect 342168 3810 342220 3816
rect 341904 480 341932 3810
rect 343560 3670 343588 64110
rect 344388 60790 344416 64110
rect 345400 60790 345428 64110
rect 344376 60784 344428 60790
rect 344376 60726 344428 60732
rect 344928 60784 344980 60790
rect 344928 60726 344980 60732
rect 345388 60784 345440 60790
rect 345388 60726 345440 60732
rect 344284 3936 344336 3942
rect 344284 3878 344336 3884
rect 343548 3664 343600 3670
rect 343548 3606 343600 3612
rect 343088 3596 343140 3602
rect 343088 3538 343140 3544
rect 343100 480 343128 3538
rect 344296 480 344324 3878
rect 344940 3602 344968 60726
rect 345480 3800 345532 3806
rect 345480 3742 345532 3748
rect 344928 3596 344980 3602
rect 344928 3538 344980 3544
rect 345492 480 345520 3742
rect 346228 3534 346256 64110
rect 346308 60784 346360 60790
rect 346308 60726 346360 60732
rect 346320 3806 346348 60726
rect 347700 3942 347728 64110
rect 348436 60790 348464 64110
rect 349448 60790 349476 64110
rect 348424 60784 348476 60790
rect 348424 60726 348476 60732
rect 349068 60784 349120 60790
rect 349068 60726 349120 60732
rect 349436 60784 349488 60790
rect 349436 60726 349488 60732
rect 350356 60784 350408 60790
rect 350356 60726 350408 60732
rect 349080 4146 349108 60726
rect 348976 4140 349028 4146
rect 348976 4082 349028 4088
rect 349068 4140 349120 4146
rect 349068 4082 349120 4088
rect 348988 4026 349016 4082
rect 350264 4072 350316 4078
rect 348988 3998 349108 4026
rect 350264 4014 350316 4020
rect 347688 3936 347740 3942
rect 347688 3878 347740 3884
rect 346308 3800 346360 3806
rect 346308 3742 346360 3748
rect 346676 3732 346728 3738
rect 346676 3674 346728 3680
rect 346216 3528 346268 3534
rect 346216 3470 346268 3476
rect 346688 480 346716 3674
rect 347872 3460 347924 3466
rect 347872 3402 347924 3408
rect 347884 480 347912 3402
rect 349080 480 349108 3998
rect 350276 480 350304 4014
rect 350368 3738 350396 60726
rect 350356 3732 350408 3738
rect 350356 3674 350408 3680
rect 350460 3466 350488 64110
rect 351840 4078 351868 64110
rect 352576 60790 352604 64110
rect 353588 60790 353616 64110
rect 352564 60784 352616 60790
rect 352564 60726 352616 60732
rect 353208 60784 353260 60790
rect 353208 60726 353260 60732
rect 353576 60784 353628 60790
rect 353576 60726 353628 60732
rect 351828 4072 351880 4078
rect 351828 4014 351880 4020
rect 351368 4004 351420 4010
rect 351368 3946 351420 3952
rect 350448 3460 350500 3466
rect 350448 3402 350500 3408
rect 351380 480 351408 3946
rect 353220 3874 353248 60726
rect 352564 3868 352616 3874
rect 352564 3810 352616 3816
rect 353208 3868 353260 3874
rect 353208 3810 353260 3816
rect 352576 480 352604 3810
rect 354508 3670 354536 64110
rect 354588 60784 354640 60790
rect 354588 60726 354640 60732
rect 354600 4010 354628 60726
rect 354588 4004 354640 4010
rect 354588 3946 354640 3952
rect 353760 3664 353812 3670
rect 353760 3606 353812 3612
rect 354496 3664 354548 3670
rect 354496 3606 354548 3612
rect 353772 480 353800 3606
rect 354956 3596 355008 3602
rect 354956 3538 355008 3544
rect 354968 480 354996 3538
rect 355980 3398 356008 64110
rect 356624 60790 356652 64110
rect 356612 60784 356664 60790
rect 356612 60726 356664 60732
rect 357256 60784 357308 60790
rect 357256 60726 357308 60732
rect 357268 3806 357296 60726
rect 356152 3800 356204 3806
rect 356152 3742 356204 3748
rect 357256 3800 357308 3806
rect 357256 3742 357308 3748
rect 355968 3392 356020 3398
rect 355968 3334 356020 3340
rect 356164 480 356192 3742
rect 357360 3618 357388 64110
rect 358544 3936 358596 3942
rect 358544 3878 358596 3884
rect 357268 3602 357388 3618
rect 357256 3596 357388 3602
rect 357308 3590 357388 3596
rect 357256 3538 357308 3544
rect 357348 3528 357400 3534
rect 357348 3470 357400 3476
rect 357360 480 357388 3470
rect 358556 480 358584 3878
rect 358740 3534 358768 64110
rect 359660 60790 359688 64110
rect 360672 60790 360700 64110
rect 359648 60784 359700 60790
rect 359648 60726 359700 60732
rect 360108 60784 360160 60790
rect 360108 60726 360160 60732
rect 360660 60784 360712 60790
rect 360660 60726 360712 60732
rect 359740 4140 359792 4146
rect 359740 4082 359792 4088
rect 358728 3528 358780 3534
rect 358728 3470 358780 3476
rect 359752 480 359780 4082
rect 360120 3942 360148 60726
rect 360108 3936 360160 3942
rect 360108 3878 360160 3884
rect 361408 3738 361436 64110
rect 361488 60784 361540 60790
rect 361488 60726 361540 60732
rect 360936 3732 360988 3738
rect 360936 3674 360988 3680
rect 361396 3732 361448 3738
rect 361396 3674 361448 3680
rect 360948 480 360976 3674
rect 361500 3194 361528 60726
rect 362880 4146 362908 64110
rect 363800 60790 363828 64110
rect 364812 60790 364840 64110
rect 363788 60784 363840 60790
rect 363788 60726 363840 60732
rect 364248 60784 364300 60790
rect 364248 60726 364300 60732
rect 364800 60784 364852 60790
rect 364800 60726 364852 60732
rect 365536 60784 365588 60790
rect 365536 60726 365588 60732
rect 362868 4140 362920 4146
rect 362868 4082 362920 4088
rect 363328 4072 363380 4078
rect 363328 4014 363380 4020
rect 362132 3460 362184 3466
rect 362132 3402 362184 3408
rect 361488 3188 361540 3194
rect 361488 3130 361540 3136
rect 362144 480 362172 3402
rect 363340 480 363368 4014
rect 364260 3262 364288 60726
rect 365548 3874 365576 60726
rect 364524 3868 364576 3874
rect 364524 3810 364576 3816
rect 365536 3868 365588 3874
rect 365536 3810 365588 3816
rect 364248 3256 364300 3262
rect 364248 3198 364300 3204
rect 364536 480 364564 3810
rect 365640 3466 365668 64110
rect 367020 4078 367048 64110
rect 367848 60790 367876 64110
rect 368860 60790 368888 64110
rect 367836 60784 367888 60790
rect 367836 60726 367888 60732
rect 368388 60784 368440 60790
rect 368388 60726 368440 60732
rect 368848 60784 368900 60790
rect 368848 60726 368900 60732
rect 369676 60784 369728 60790
rect 369676 60726 369728 60732
rect 367008 4072 367060 4078
rect 367008 4014 367060 4020
rect 365720 4004 365772 4010
rect 365720 3946 365772 3952
rect 365628 3460 365680 3466
rect 365628 3402 365680 3408
rect 365732 480 365760 3946
rect 368400 3670 368428 60726
rect 369216 3800 369268 3806
rect 369216 3742 369268 3748
rect 366916 3664 366968 3670
rect 366916 3606 366968 3612
rect 368388 3664 368440 3670
rect 368388 3606 368440 3612
rect 366928 480 366956 3606
rect 368020 3392 368072 3398
rect 368020 3334 368072 3340
rect 368032 480 368060 3334
rect 369228 480 369256 3742
rect 369688 3330 369716 60726
rect 369780 3398 369808 64110
rect 371160 3806 371188 64110
rect 371896 60790 371924 64110
rect 372908 60790 372936 64110
rect 371884 60784 371936 60790
rect 371884 60726 371936 60732
rect 372528 60784 372580 60790
rect 372528 60726 372580 60732
rect 372896 60784 372948 60790
rect 372896 60726 372948 60732
rect 371148 3800 371200 3806
rect 371148 3742 371200 3748
rect 372540 3602 372568 60726
rect 372804 3936 372856 3942
rect 372804 3878 372856 3884
rect 370412 3596 370464 3602
rect 370412 3538 370464 3544
rect 372528 3596 372580 3602
rect 372528 3538 372580 3544
rect 369768 3392 369820 3398
rect 369768 3334 369820 3340
rect 369676 3324 369728 3330
rect 369676 3266 369728 3272
rect 370424 480 370452 3538
rect 371608 3528 371660 3534
rect 371608 3470 371660 3476
rect 371620 480 371648 3470
rect 372816 480 372844 3878
rect 373828 3534 373856 64110
rect 373908 60784 373960 60790
rect 373908 60726 373960 60732
rect 373920 4010 373948 60726
rect 373908 4004 373960 4010
rect 373908 3946 373960 3952
rect 375300 3738 375328 64110
rect 376036 60790 376064 64110
rect 377048 60790 377076 64110
rect 376024 60784 376076 60790
rect 376024 60726 376076 60732
rect 376668 60784 376720 60790
rect 376668 60726 376720 60732
rect 377036 60784 377088 60790
rect 377036 60726 377088 60732
rect 377956 60784 378008 60790
rect 377956 60726 378008 60732
rect 376392 4140 376444 4146
rect 376392 4082 376444 4088
rect 375196 3732 375248 3738
rect 375196 3674 375248 3680
rect 375288 3732 375340 3738
rect 375288 3674 375340 3680
rect 373816 3528 373868 3534
rect 373816 3470 373868 3476
rect 374000 3188 374052 3194
rect 374000 3130 374052 3136
rect 374012 480 374040 3130
rect 375208 480 375236 3674
rect 376404 480 376432 4082
rect 376680 3126 376708 60726
rect 377968 4146 377996 60726
rect 377956 4140 378008 4146
rect 377956 4082 378008 4088
rect 378060 3942 378088 64110
rect 378048 3936 378100 3942
rect 378048 3878 378100 3884
rect 379440 3874 379468 64110
rect 380084 60790 380112 64110
rect 380774 63866 380802 64124
rect 381800 64110 382228 64138
rect 382812 64110 383148 64138
rect 383824 64110 384160 64138
rect 384928 64110 384988 64138
rect 385940 64110 386368 64138
rect 386952 64110 387288 64138
rect 387964 64110 388300 64138
rect 388976 64110 389036 64138
rect 389988 64110 390508 64138
rect 391000 64110 391336 64138
rect 392012 64110 392348 64138
rect 393024 64110 393176 64138
rect 394036 64110 394648 64138
rect 395048 64110 395384 64138
rect 396152 64110 396488 64138
rect 397164 64110 397408 64138
rect 398176 64110 398788 64138
rect 399188 64110 399524 64138
rect 400200 64110 400536 64138
rect 401212 64110 401548 64138
rect 402224 64110 402560 64138
rect 403236 64110 403572 64138
rect 380728 63838 380802 63866
rect 380072 60784 380124 60790
rect 380072 60726 380124 60732
rect 378784 3868 378836 3874
rect 378784 3810 378836 3816
rect 379428 3868 379480 3874
rect 379428 3810 379480 3816
rect 377588 3256 377640 3262
rect 377588 3198 377640 3204
rect 376668 3120 376720 3126
rect 376668 3062 376720 3068
rect 377600 480 377628 3198
rect 378796 480 378824 3810
rect 380728 3466 380756 63838
rect 380808 60784 380860 60790
rect 380808 60726 380860 60732
rect 379980 3460 380032 3466
rect 379980 3402 380032 3408
rect 380716 3460 380768 3466
rect 380716 3402 380768 3408
rect 379992 480 380020 3402
rect 380820 3194 380848 60726
rect 382200 4078 382228 64110
rect 383120 60790 383148 64110
rect 384132 60790 384160 64110
rect 383108 60784 383160 60790
rect 383108 60726 383160 60732
rect 383568 60784 383620 60790
rect 383568 60726 383620 60732
rect 384120 60784 384172 60790
rect 384120 60726 384172 60732
rect 384856 60784 384908 60790
rect 384856 60726 384908 60732
rect 381176 4072 381228 4078
rect 381176 4014 381228 4020
rect 382188 4072 382240 4078
rect 382188 4014 382240 4020
rect 380808 3188 380860 3194
rect 380808 3130 380860 3136
rect 381188 480 381216 4014
rect 383580 3670 383608 60726
rect 382372 3664 382424 3670
rect 382372 3606 382424 3612
rect 383568 3664 383620 3670
rect 383568 3606 383620 3612
rect 382384 480 382412 3606
rect 384672 3392 384724 3398
rect 384672 3334 384724 3340
rect 383568 3324 383620 3330
rect 383568 3266 383620 3272
rect 383580 480 383608 3266
rect 384684 480 384712 3334
rect 384868 2990 384896 60726
rect 384960 3058 384988 64110
rect 385868 3800 385920 3806
rect 385868 3742 385920 3748
rect 384948 3052 385000 3058
rect 384948 2994 385000 3000
rect 384856 2984 384908 2990
rect 384856 2926 384908 2932
rect 385880 480 385908 3742
rect 386340 3262 386368 64110
rect 387260 60790 387288 64110
rect 388272 60790 388300 64110
rect 387248 60784 387300 60790
rect 387248 60726 387300 60732
rect 387708 60784 387760 60790
rect 387708 60726 387760 60732
rect 388260 60784 388312 60790
rect 388260 60726 388312 60732
rect 387720 3806 387748 60726
rect 388260 4004 388312 4010
rect 388260 3946 388312 3952
rect 387708 3800 387760 3806
rect 387708 3742 387760 3748
rect 387064 3596 387116 3602
rect 387064 3538 387116 3544
rect 386328 3256 386380 3262
rect 386328 3198 386380 3204
rect 387076 480 387104 3538
rect 388272 480 388300 3946
rect 389008 3602 389036 64110
rect 389088 60784 389140 60790
rect 389088 60726 389140 60732
rect 388996 3596 389048 3602
rect 388996 3538 389048 3544
rect 389100 3330 389128 60726
rect 390480 4010 390508 64110
rect 391308 60790 391336 64110
rect 392320 60790 392348 64110
rect 391296 60784 391348 60790
rect 391296 60726 391348 60732
rect 391848 60784 391900 60790
rect 391848 60726 391900 60732
rect 392308 60784 392360 60790
rect 392308 60726 392360 60732
rect 390468 4004 390520 4010
rect 390468 3946 390520 3952
rect 390652 3732 390704 3738
rect 390652 3674 390704 3680
rect 389456 3528 389508 3534
rect 389456 3470 389508 3476
rect 389088 3324 389140 3330
rect 389088 3266 389140 3272
rect 389468 480 389496 3470
rect 390664 480 390692 3674
rect 391860 3398 391888 60726
rect 393044 4140 393096 4146
rect 393044 4082 393096 4088
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391848 3120 391900 3126
rect 391848 3062 391900 3068
rect 391860 480 391888 3062
rect 393056 480 393084 4082
rect 393148 3534 393176 64110
rect 393228 60784 393280 60790
rect 393228 60726 393280 60732
rect 393136 3528 393188 3534
rect 393136 3470 393188 3476
rect 393240 3126 393268 60726
rect 394240 3936 394292 3942
rect 394240 3878 394292 3884
rect 393228 3120 393280 3126
rect 393228 3062 393280 3068
rect 394252 480 394280 3878
rect 394620 3738 394648 64110
rect 395356 60790 395384 64110
rect 396460 60790 396488 64110
rect 395344 60784 395396 60790
rect 395344 60726 395396 60732
rect 395988 60784 396040 60790
rect 395988 60726 396040 60732
rect 396448 60784 396500 60790
rect 396448 60726 396500 60732
rect 397276 60784 397328 60790
rect 397276 60726 397328 60732
rect 396000 4146 396028 60726
rect 395988 4140 396040 4146
rect 395988 4082 396040 4088
rect 397288 3942 397316 60726
rect 397276 3936 397328 3942
rect 397276 3878 397328 3884
rect 397380 3874 397408 64110
rect 395436 3868 395488 3874
rect 395436 3810 395488 3816
rect 397368 3868 397420 3874
rect 397368 3810 397420 3816
rect 394608 3732 394660 3738
rect 394608 3674 394660 3680
rect 395448 480 395476 3810
rect 397828 3460 397880 3466
rect 397828 3402 397880 3408
rect 396632 3188 396684 3194
rect 396632 3130 396684 3136
rect 396644 480 396672 3130
rect 397840 480 397868 3402
rect 398760 3194 398788 64110
rect 399496 61742 399524 64110
rect 399484 61736 399536 61742
rect 399484 61678 399536 61684
rect 400508 60790 400536 64110
rect 400496 60784 400548 60790
rect 400496 60726 400548 60732
rect 401416 60784 401468 60790
rect 401416 60726 401468 60732
rect 401428 4078 401456 60726
rect 399024 4072 399076 4078
rect 399024 4014 399076 4020
rect 401416 4072 401468 4078
rect 401416 4014 401468 4020
rect 398748 3188 398800 3194
rect 398748 3130 398800 3136
rect 399036 480 399064 4014
rect 401520 3670 401548 64110
rect 402532 61606 402560 64110
rect 402520 61600 402572 61606
rect 402520 61542 402572 61548
rect 403544 60790 403572 64110
rect 404234 63866 404262 64124
rect 405260 64110 405596 64138
rect 406272 64110 406608 64138
rect 407376 64110 407712 64138
rect 408388 64110 408448 64138
rect 409400 64110 409828 64138
rect 410412 64110 410748 64138
rect 411424 64110 411760 64138
rect 412436 64110 412588 64138
rect 413448 64110 413968 64138
rect 414460 64110 414796 64138
rect 415472 64110 415808 64138
rect 416484 64110 416636 64138
rect 417496 64110 417832 64138
rect 418600 64110 418936 64138
rect 419612 64110 419948 64138
rect 420624 64110 420868 64138
rect 421636 64110 422248 64138
rect 422648 64110 422984 64138
rect 423660 64110 423996 64138
rect 424672 64110 425008 64138
rect 425684 64110 426388 64138
rect 426696 64110 427032 64138
rect 427708 64110 427768 64138
rect 428720 64110 429148 64138
rect 429824 64110 430160 64138
rect 430836 64110 431172 64138
rect 404188 63838 404262 63866
rect 403532 60784 403584 60790
rect 403532 60726 403584 60732
rect 400220 3664 400272 3670
rect 400220 3606 400272 3612
rect 401508 3664 401560 3670
rect 401508 3606 401560 3612
rect 400232 480 400260 3606
rect 404188 3466 404216 63838
rect 405568 61470 405596 64110
rect 405556 61464 405608 61470
rect 405556 61406 405608 61412
rect 406580 60790 406608 64110
rect 407684 60790 407712 64110
rect 408420 61402 408448 64110
rect 408408 61396 408460 61402
rect 408408 61338 408460 61344
rect 404268 60784 404320 60790
rect 404268 60726 404320 60732
rect 406568 60784 406620 60790
rect 406568 60726 406620 60732
rect 407028 60784 407080 60790
rect 407028 60726 407080 60732
rect 407672 60784 407724 60790
rect 407672 60726 407724 60732
rect 408408 60784 408460 60790
rect 408408 60726 408460 60732
rect 404176 3460 404228 3466
rect 404176 3402 404228 3408
rect 404280 3262 404308 60726
rect 404912 3800 404964 3806
rect 404912 3742 404964 3748
rect 403716 3256 403768 3262
rect 403716 3198 403768 3204
rect 404268 3256 404320 3262
rect 404268 3198 404320 3204
rect 402520 3052 402572 3058
rect 402520 2994 402572 3000
rect 401324 2984 401376 2990
rect 401324 2926 401376 2932
rect 401336 480 401364 2926
rect 402532 480 402560 2994
rect 403728 480 403756 3198
rect 404924 480 404952 3742
rect 407040 3330 407068 60726
rect 408420 3806 408448 60726
rect 408500 4004 408552 4010
rect 408500 3946 408552 3952
rect 408408 3800 408460 3806
rect 408408 3742 408460 3748
rect 407304 3596 407356 3602
rect 407304 3538 407356 3544
rect 406108 3324 406160 3330
rect 406108 3266 406160 3272
rect 407028 3324 407080 3330
rect 407028 3266 407080 3272
rect 406120 480 406148 3266
rect 407316 480 407344 3538
rect 408512 480 408540 3946
rect 409800 3602 409828 64110
rect 410720 60790 410748 64110
rect 411732 61538 411760 64110
rect 411720 61532 411772 61538
rect 411720 61474 411772 61480
rect 410708 60784 410760 60790
rect 410708 60726 410760 60732
rect 411168 60784 411220 60790
rect 411168 60726 411220 60732
rect 411180 4010 411208 60726
rect 411168 4004 411220 4010
rect 411168 3946 411220 3952
rect 409788 3596 409840 3602
rect 409788 3538 409840 3544
rect 412088 3528 412140 3534
rect 412088 3470 412140 3476
rect 409696 3392 409748 3398
rect 409696 3334 409748 3340
rect 409708 480 409736 3334
rect 410892 3120 410944 3126
rect 410892 3062 410944 3068
rect 410904 480 410932 3062
rect 412100 480 412128 3470
rect 412560 3398 412588 64110
rect 413940 3738 413968 64110
rect 414768 61810 414796 64110
rect 414756 61804 414808 61810
rect 414756 61746 414808 61752
rect 415780 60790 415808 64110
rect 415768 60784 415820 60790
rect 415768 60726 415820 60732
rect 414480 4140 414532 4146
rect 414480 4082 414532 4088
rect 413284 3732 413336 3738
rect 413284 3674 413336 3680
rect 413928 3732 413980 3738
rect 413928 3674 413980 3680
rect 412548 3392 412600 3398
rect 412548 3334 412600 3340
rect 413296 480 413324 3674
rect 414492 480 414520 4082
rect 415676 3936 415728 3942
rect 415676 3878 415728 3884
rect 415688 480 415716 3878
rect 416608 3534 416636 64110
rect 417804 61674 417832 64110
rect 418252 61736 418304 61742
rect 418252 61678 418304 61684
rect 417792 61668 417844 61674
rect 417792 61610 417844 61616
rect 416688 60784 416740 60790
rect 416688 60726 416740 60732
rect 416596 3528 416648 3534
rect 416596 3470 416648 3476
rect 416700 3058 416728 60726
rect 416872 3868 416924 3874
rect 416872 3810 416924 3816
rect 416688 3052 416740 3058
rect 416688 2994 416740 3000
rect 416884 480 416912 3810
rect 417976 3188 418028 3194
rect 417976 3130 418028 3136
rect 417988 480 418016 3130
rect 418264 610 418292 61678
rect 418908 60790 418936 64110
rect 419920 60790 419948 64110
rect 420840 61742 420868 64110
rect 420828 61736 420880 61742
rect 420828 61678 420880 61684
rect 418896 60784 418948 60790
rect 418896 60726 418948 60732
rect 419448 60784 419500 60790
rect 419448 60726 419500 60732
rect 419908 60784 419960 60790
rect 419908 60726 419960 60732
rect 420828 60784 420880 60790
rect 420828 60726 420880 60732
rect 419460 3942 419488 60726
rect 420840 4146 420868 60726
rect 420828 4140 420880 4146
rect 420828 4082 420880 4088
rect 420368 4072 420420 4078
rect 420368 4014 420420 4020
rect 419448 3936 419500 3942
rect 419448 3878 419500 3884
rect 418252 604 418304 610
rect 418252 546 418304 552
rect 419172 604 419224 610
rect 419172 546 419224 552
rect 419184 480 419212 546
rect 420380 480 420408 4014
rect 421564 3664 421616 3670
rect 421564 3606 421616 3612
rect 421576 480 421604 3606
rect 422220 3126 422248 64110
rect 422392 61600 422444 61606
rect 422392 61542 422444 61548
rect 422300 3392 422352 3398
rect 422300 3334 422352 3340
rect 422312 3194 422340 3334
rect 422300 3188 422352 3194
rect 422300 3130 422352 3136
rect 422208 3120 422260 3126
rect 422208 3062 422260 3068
rect 422404 626 422432 61542
rect 422956 60790 422984 64110
rect 423968 61946 423996 64110
rect 423956 61940 424008 61946
rect 423956 61882 424008 61888
rect 422944 60784 422996 60790
rect 422944 60726 422996 60732
rect 423588 60784 423640 60790
rect 423588 60726 423640 60732
rect 423600 4078 423628 60726
rect 423588 4072 423640 4078
rect 423588 4014 423640 4020
rect 424980 3874 425008 64110
rect 425152 61464 425204 61470
rect 425152 61406 425204 61412
rect 424968 3868 425020 3874
rect 424968 3810 425020 3816
rect 425164 3466 425192 61406
rect 426360 3618 426388 64110
rect 427004 61470 427032 64110
rect 426992 61464 427044 61470
rect 426992 61406 427044 61412
rect 426360 3590 426480 3618
rect 426452 3466 426480 3590
rect 425060 3460 425112 3466
rect 425060 3402 425112 3408
rect 425152 3460 425204 3466
rect 425152 3402 425204 3408
rect 426348 3460 426400 3466
rect 426348 3402 426400 3408
rect 426440 3460 426492 3466
rect 426440 3402 426492 3408
rect 425072 3346 425100 3402
rect 425072 3318 425192 3346
rect 423956 3256 424008 3262
rect 423956 3198 424008 3204
rect 422404 598 422800 626
rect 422772 480 422800 598
rect 423968 480 423996 3198
rect 425164 480 425192 3318
rect 426360 480 426388 3402
rect 427544 3324 427596 3330
rect 427544 3266 427596 3272
rect 427556 480 427584 3266
rect 427740 3262 427768 64110
rect 428740 3800 428792 3806
rect 428740 3742 428792 3748
rect 427728 3256 427780 3262
rect 427728 3198 427780 3204
rect 428752 480 428780 3742
rect 429120 3670 429148 64110
rect 430132 61606 430160 64110
rect 430120 61600 430172 61606
rect 430120 61542 430172 61548
rect 429200 61396 429252 61402
rect 429200 61338 429252 61344
rect 429108 3664 429160 3670
rect 429108 3606 429160 3612
rect 429212 610 429240 61338
rect 431144 60790 431172 64110
rect 431834 63866 431862 64124
rect 432860 64110 433196 64138
rect 433872 64110 434208 64138
rect 434884 64110 435220 64138
rect 435896 64110 436048 64138
rect 436908 64110 437428 64138
rect 437920 64110 438256 64138
rect 438932 64110 439268 64138
rect 440036 64110 440188 64138
rect 441048 64110 441568 64138
rect 442060 64110 442396 64138
rect 443072 64110 443408 64138
rect 444084 64110 444236 64138
rect 445096 64110 445432 64138
rect 446108 64110 446444 64138
rect 447120 64110 447456 64138
rect 448132 64110 448376 64138
rect 449144 64110 449848 64138
rect 450156 64110 450492 64138
rect 451260 64110 451596 64138
rect 452272 64110 452608 64138
rect 453284 64110 453988 64138
rect 454296 64110 454632 64138
rect 455308 64110 455368 64138
rect 456320 64110 456748 64138
rect 457332 64110 457668 64138
rect 458344 64110 458680 64138
rect 459356 64110 459508 64138
rect 460368 64110 460704 64138
rect 461380 64110 461716 64138
rect 462484 64110 462820 64138
rect 463496 64110 463648 64138
rect 464508 64110 465028 64138
rect 465520 64110 465856 64138
rect 466532 64110 466868 64138
rect 467544 64110 467788 64138
rect 468556 64110 469168 64138
rect 469568 64110 469904 64138
rect 470580 64110 470916 64138
rect 471592 64110 471928 64138
rect 472604 64110 473308 64138
rect 473708 64110 474044 64138
rect 474720 64110 475056 64138
rect 475732 64110 476068 64138
rect 476744 64110 477448 64138
rect 477756 64110 478092 64138
rect 478768 64110 478828 64138
rect 479780 64110 480208 64138
rect 480792 64110 481128 64138
rect 481804 64110 482140 64138
rect 482816 64110 482968 64138
rect 483828 64110 484164 64138
rect 484932 64110 485268 64138
rect 485944 64110 486280 64138
rect 486956 64110 487108 64138
rect 487968 64110 488488 64138
rect 488980 64110 489316 64138
rect 489992 64110 490328 64138
rect 491004 64110 491248 64138
rect 492016 64110 492628 64138
rect 493028 64110 493364 64138
rect 494040 64110 494376 64138
rect 495052 64110 495388 64138
rect 496156 64110 496492 64138
rect 497168 64110 497504 64138
rect 498180 64110 498516 64138
rect 499192 64110 499436 64138
rect 500204 64110 500908 64138
rect 501216 64110 501552 64138
rect 502228 64110 502288 64138
rect 503240 64110 503576 64138
rect 504252 64110 504588 64138
rect 505264 64110 505600 64138
rect 506276 64110 506428 64138
rect 507380 64110 507808 64138
rect 508392 64110 508728 64138
rect 509404 64110 509740 64138
rect 510416 64110 510568 64138
rect 511428 64110 511948 64138
rect 512440 64110 512776 64138
rect 513452 64110 513788 64138
rect 514464 64110 514708 64138
rect 515476 64110 515812 64138
rect 516488 64110 516824 64138
rect 517500 64110 517836 64138
rect 518604 64110 518756 64138
rect 519616 64110 519952 64138
rect 520628 64110 520964 64138
rect 521640 64110 521976 64138
rect 522652 64110 522988 64138
rect 523664 64110 524368 64138
rect 524676 64110 525012 64138
rect 525688 64110 525748 64138
rect 526700 64110 527036 64138
rect 527712 64110 528048 64138
rect 528724 64110 529060 64138
rect 529828 64110 529888 64138
rect 530840 64110 531176 64138
rect 531852 64110 532188 64138
rect 532864 64110 533200 64138
rect 533876 64110 534028 64138
rect 534888 64110 535224 64138
rect 535900 64110 536236 64138
rect 536912 64110 537248 64138
rect 537924 64110 538076 64138
rect 431788 63838 431862 63866
rect 431132 60784 431184 60790
rect 431132 60726 431184 60732
rect 431788 3602 431816 63838
rect 433168 61402 433196 64110
rect 433432 61532 433484 61538
rect 433432 61474 433484 61480
rect 433156 61396 433208 61402
rect 433156 61338 433208 61344
rect 431868 60784 431920 60790
rect 431868 60726 431920 60732
rect 431880 3806 431908 60726
rect 432328 4004 432380 4010
rect 432328 3946 432380 3952
rect 431868 3800 431920 3806
rect 431868 3742 431920 3748
rect 431132 3596 431184 3602
rect 431132 3538 431184 3544
rect 431776 3596 431828 3602
rect 431776 3538 431828 3544
rect 429200 604 429252 610
rect 429200 546 429252 552
rect 429936 604 429988 610
rect 429936 546 429988 552
rect 429948 480 429976 546
rect 431144 480 431172 3538
rect 432340 480 432368 3946
rect 433444 3482 433472 61474
rect 434180 60790 434208 64110
rect 435192 60790 435220 64110
rect 436020 61538 436048 64110
rect 436192 61804 436244 61810
rect 436192 61746 436244 61752
rect 436008 61532 436060 61538
rect 436008 61474 436060 61480
rect 434168 60784 434220 60790
rect 434168 60726 434220 60732
rect 434628 60784 434680 60790
rect 434628 60726 434680 60732
rect 435180 60784 435232 60790
rect 435180 60726 435232 60732
rect 436008 60784 436060 60790
rect 436008 60726 436060 60732
rect 434640 3482 434668 60726
rect 435824 3732 435876 3738
rect 435824 3674 435876 3680
rect 433444 3454 433564 3482
rect 434640 3454 434760 3482
rect 433536 480 433564 3454
rect 434732 3398 434760 3454
rect 434720 3392 434772 3398
rect 434720 3334 434772 3340
rect 434628 3324 434680 3330
rect 434628 3266 434680 3272
rect 434640 480 434668 3266
rect 435836 480 435864 3674
rect 436020 3194 436048 60726
rect 436008 3188 436060 3194
rect 436008 3130 436060 3136
rect 436204 610 436232 61746
rect 437400 3330 437428 64110
rect 438228 60790 438256 64110
rect 439240 61878 439268 64110
rect 439228 61872 439280 61878
rect 439228 61814 439280 61820
rect 438216 60784 438268 60790
rect 438216 60726 438268 60732
rect 438768 60784 438820 60790
rect 438768 60726 438820 60732
rect 438780 4010 438808 60726
rect 438768 4004 438820 4010
rect 438768 3946 438820 3952
rect 440160 3534 440188 64110
rect 440332 61668 440384 61674
rect 440332 61610 440384 61616
rect 439412 3528 439464 3534
rect 439412 3470 439464 3476
rect 440148 3528 440200 3534
rect 440148 3470 440200 3476
rect 437388 3324 437440 3330
rect 437388 3266 437440 3272
rect 438216 3052 438268 3058
rect 438216 2994 438268 3000
rect 436192 604 436244 610
rect 436192 546 436244 552
rect 437020 604 437072 610
rect 437020 546 437072 552
rect 437032 480 437060 546
rect 438228 480 438256 2994
rect 439424 480 439452 3470
rect 440344 626 440372 61610
rect 441540 3738 441568 64110
rect 442368 61810 442396 64110
rect 442356 61804 442408 61810
rect 442356 61746 442408 61752
rect 443184 61736 443236 61742
rect 443184 61678 443236 61684
rect 443000 4140 443052 4146
rect 443000 4082 443052 4088
rect 441804 3936 441856 3942
rect 441804 3878 441856 3884
rect 441528 3732 441580 3738
rect 441528 3674 441580 3680
rect 440344 598 440648 626
rect 440620 480 440648 598
rect 441816 480 441844 3878
rect 443012 480 443040 4082
rect 443196 3210 443224 61678
rect 443380 60790 443408 64110
rect 443368 60784 443420 60790
rect 443368 60726 443420 60732
rect 444208 3942 444236 64110
rect 445404 61742 445432 64110
rect 445392 61736 445444 61742
rect 445392 61678 445444 61684
rect 446416 60790 446444 64110
rect 447140 61940 447192 61946
rect 447140 61882 447192 61888
rect 444288 60784 444340 60790
rect 444288 60726 444340 60732
rect 446404 60784 446456 60790
rect 446404 60726 446456 60732
rect 447048 60784 447100 60790
rect 447048 60726 447100 60732
rect 444196 3936 444248 3942
rect 444196 3878 444248 3884
rect 443196 3182 444236 3210
rect 444208 480 444236 3182
rect 444300 2854 444328 60726
rect 447060 4078 447088 60726
rect 446588 4072 446640 4078
rect 446588 4014 446640 4020
rect 447048 4072 447100 4078
rect 447048 4014 447100 4020
rect 445392 3120 445444 3126
rect 445392 3062 445444 3068
rect 444288 2848 444340 2854
rect 444288 2790 444340 2796
rect 445404 480 445432 3062
rect 446600 480 446628 4014
rect 447152 610 447180 61882
rect 447428 60790 447456 64110
rect 447416 60784 447468 60790
rect 447416 60726 447468 60732
rect 448348 4826 448376 64110
rect 448428 60784 448480 60790
rect 448428 60726 448480 60732
rect 448336 4820 448388 4826
rect 448336 4762 448388 4768
rect 448440 2922 448468 60726
rect 449820 4146 449848 64110
rect 450464 60790 450492 64110
rect 451464 61464 451516 61470
rect 451464 61406 451516 61412
rect 450452 60784 450504 60790
rect 450452 60726 450504 60732
rect 451188 60784 451240 60790
rect 451188 60726 451240 60732
rect 449808 4140 449860 4146
rect 449808 4082 449860 4088
rect 448980 3868 449032 3874
rect 448980 3810 449032 3816
rect 448428 2916 448480 2922
rect 448428 2858 448480 2864
rect 447140 604 447192 610
rect 447140 546 447192 552
rect 447784 604 447836 610
rect 447784 546 447836 552
rect 447796 480 447824 546
rect 448992 480 449020 3810
rect 450176 3460 450228 3466
rect 450176 3402 450228 3408
rect 450188 480 450216 3402
rect 451200 2990 451228 60726
rect 451188 2984 451240 2990
rect 451188 2926 451240 2932
rect 451476 626 451504 61406
rect 451568 60790 451596 64110
rect 451556 60784 451608 60790
rect 451556 60726 451608 60732
rect 452476 60784 452528 60790
rect 452476 60726 452528 60732
rect 452488 6882 452516 60726
rect 452304 6854 452516 6882
rect 452304 3058 452332 6854
rect 452580 3262 452608 64110
rect 453960 3670 453988 64110
rect 454604 61674 454632 64110
rect 454592 61668 454644 61674
rect 454592 61610 454644 61616
rect 454224 61600 454276 61606
rect 454224 61542 454276 61548
rect 453672 3664 453724 3670
rect 453672 3606 453724 3612
rect 453948 3664 454000 3670
rect 453948 3606 454000 3612
rect 452476 3256 452528 3262
rect 452476 3198 452528 3204
rect 452568 3256 452620 3262
rect 452568 3198 452620 3204
rect 452292 3052 452344 3058
rect 452292 2994 452344 3000
rect 451384 598 451504 626
rect 451384 592 451412 598
rect 451292 564 451412 592
rect 451292 480 451320 564
rect 452488 480 452516 3198
rect 453684 480 453712 3606
rect 454236 610 454264 61542
rect 455340 3466 455368 64110
rect 456720 3806 456748 64110
rect 457640 61606 457668 64110
rect 457628 61600 457680 61606
rect 457628 61542 457680 61548
rect 458364 61396 458416 61402
rect 458364 61338 458416 61344
rect 456064 3800 456116 3806
rect 456064 3742 456116 3748
rect 456708 3800 456760 3806
rect 456708 3742 456760 3748
rect 455328 3460 455380 3466
rect 455328 3402 455380 3408
rect 454224 604 454276 610
rect 454224 546 454276 552
rect 454868 604 454920 610
rect 454868 546 454920 552
rect 454880 480 454908 546
rect 456076 480 456104 3742
rect 457260 3596 457312 3602
rect 457260 3538 457312 3544
rect 457272 480 457300 3538
rect 458376 592 458404 61338
rect 458652 60790 458680 64110
rect 458640 60784 458692 60790
rect 458640 60726 458692 60732
rect 459376 60784 459428 60790
rect 459376 60726 459428 60732
rect 459388 3126 459416 60726
rect 459480 3874 459508 64110
rect 460676 61470 460704 64110
rect 461032 61532 461084 61538
rect 461032 61474 461084 61480
rect 460664 61464 460716 61470
rect 460664 61406 460716 61412
rect 459468 3868 459520 3874
rect 459468 3810 459520 3816
rect 459652 3392 459704 3398
rect 459652 3334 459704 3340
rect 459376 3120 459428 3126
rect 459376 3062 459428 3068
rect 458376 564 458496 592
rect 458468 480 458496 564
rect 459664 480 459692 3334
rect 460848 3188 460900 3194
rect 460848 3130 460900 3136
rect 460860 480 460888 3130
rect 461044 610 461072 61474
rect 461688 60790 461716 64110
rect 462792 60790 462820 64110
rect 463620 61402 463648 64110
rect 463608 61396 463660 61402
rect 463608 61338 463660 61344
rect 461676 60784 461728 60790
rect 461676 60726 461728 60732
rect 462228 60784 462280 60790
rect 462228 60726 462280 60732
rect 462780 60784 462832 60790
rect 462780 60726 462832 60732
rect 463608 60784 463660 60790
rect 463608 60726 463660 60732
rect 462240 3194 462268 60726
rect 463620 3398 463648 60726
rect 465000 4010 465028 64110
rect 465172 61872 465224 61878
rect 465172 61814 465224 61820
rect 464436 4004 464488 4010
rect 464436 3946 464488 3952
rect 464988 4004 465040 4010
rect 464988 3946 465040 3952
rect 463608 3392 463660 3398
rect 463608 3334 463660 3340
rect 463240 3324 463292 3330
rect 463240 3266 463292 3272
rect 462228 3188 462280 3194
rect 462228 3130 462280 3136
rect 461032 604 461084 610
rect 461032 546 461084 552
rect 462044 604 462096 610
rect 462044 546 462096 552
rect 462056 480 462084 546
rect 463252 480 463280 3266
rect 464448 480 464476 3946
rect 465184 626 465212 61814
rect 465828 60790 465856 64110
rect 466840 61538 466868 64110
rect 466828 61532 466880 61538
rect 466828 61474 466880 61480
rect 465816 60784 465868 60790
rect 465816 60726 465868 60732
rect 466368 60784 466420 60790
rect 466368 60726 466420 60732
rect 466380 3330 466408 60726
rect 467760 3602 467788 64110
rect 467932 61804 467984 61810
rect 467932 61746 467984 61752
rect 467840 3732 467892 3738
rect 467840 3674 467892 3680
rect 467748 3596 467800 3602
rect 467748 3538 467800 3544
rect 466828 3528 466880 3534
rect 466828 3470 466880 3476
rect 466368 3324 466420 3330
rect 466368 3266 466420 3272
rect 465184 598 465672 626
rect 465644 480 465672 598
rect 466840 480 466868 3470
rect 467852 3346 467880 3674
rect 467944 3534 467972 61746
rect 469140 3738 469168 64110
rect 469876 60790 469904 64110
rect 470888 60790 470916 64110
rect 471900 61810 471928 64110
rect 471888 61804 471940 61810
rect 471888 61746 471940 61752
rect 472072 61736 472124 61742
rect 472072 61678 472124 61684
rect 469864 60784 469916 60790
rect 469864 60726 469916 60732
rect 470508 60784 470560 60790
rect 470508 60726 470560 60732
rect 470876 60784 470928 60790
rect 470876 60726 470928 60732
rect 471888 60784 471940 60790
rect 471888 60726 471940 60732
rect 470520 5030 470548 60726
rect 470508 5024 470560 5030
rect 470508 4966 470560 4972
rect 471900 4010 471928 60726
rect 469496 4004 469548 4010
rect 469496 3946 469548 3952
rect 471888 4004 471940 4010
rect 471888 3946 471940 3952
rect 469128 3732 469180 3738
rect 469128 3674 469180 3680
rect 469312 3596 469364 3602
rect 469312 3538 469364 3544
rect 467932 3528 467984 3534
rect 467932 3470 467984 3476
rect 469128 3528 469180 3534
rect 469128 3470 469180 3476
rect 467852 3318 467972 3346
rect 467944 480 467972 3318
rect 469140 480 469168 3470
rect 469324 3398 469352 3538
rect 469312 3392 469364 3398
rect 469312 3334 469364 3340
rect 469404 3392 469456 3398
rect 469404 3334 469456 3340
rect 469416 3194 469444 3334
rect 469508 3194 469536 3946
rect 471520 3936 471572 3942
rect 471520 3878 471572 3884
rect 469404 3188 469456 3194
rect 469404 3130 469456 3136
rect 469496 3188 469548 3194
rect 469496 3130 469548 3136
rect 470324 2848 470376 2854
rect 470324 2790 470376 2796
rect 470336 480 470364 2790
rect 471532 480 471560 3878
rect 472084 610 472112 61678
rect 473280 5302 473308 64110
rect 474016 60790 474044 64110
rect 475028 62014 475056 64110
rect 475016 62008 475068 62014
rect 475016 61950 475068 61956
rect 474004 60784 474056 60790
rect 474004 60726 474056 60732
rect 474648 60784 474700 60790
rect 474648 60726 474700 60732
rect 473268 5296 473320 5302
rect 473268 5238 473320 5244
rect 474660 4078 474688 60726
rect 476040 5166 476068 64110
rect 476028 5160 476080 5166
rect 476028 5102 476080 5108
rect 476304 4820 476356 4826
rect 476304 4762 476356 4768
rect 473912 4072 473964 4078
rect 473912 4014 473964 4020
rect 474648 4072 474700 4078
rect 474648 4014 474700 4020
rect 472072 604 472124 610
rect 472072 546 472124 552
rect 472716 604 472768 610
rect 472716 546 472768 552
rect 472728 480 472756 546
rect 473924 480 473952 4014
rect 475108 2916 475160 2922
rect 475108 2858 475160 2864
rect 475120 480 475148 2858
rect 476316 480 476344 4762
rect 477420 3942 477448 64110
rect 478064 61742 478092 64110
rect 478052 61736 478104 61742
rect 478052 61678 478104 61684
rect 478800 5234 478828 64110
rect 478788 5228 478840 5234
rect 478788 5170 478840 5176
rect 480180 4146 480208 64110
rect 481100 60790 481128 64110
rect 482112 60790 482140 64110
rect 481088 60784 481140 60790
rect 481088 60726 481140 60732
rect 481548 60784 481600 60790
rect 481548 60726 481600 60732
rect 482100 60784 482152 60790
rect 482100 60726 482152 60732
rect 482836 60784 482888 60790
rect 482836 60726 482888 60732
rect 477500 4140 477552 4146
rect 477500 4082 477552 4088
rect 480168 4140 480220 4146
rect 480168 4082 480220 4088
rect 477408 3936 477460 3942
rect 477408 3878 477460 3884
rect 477512 480 477540 4082
rect 481560 3262 481588 60726
rect 482848 5370 482876 60726
rect 482836 5364 482888 5370
rect 482836 5306 482888 5312
rect 482940 3670 482968 64110
rect 484136 61946 484164 64110
rect 484124 61940 484176 61946
rect 484124 61882 484176 61888
rect 483664 61804 483716 61810
rect 483664 61746 483716 61752
rect 483020 61668 483072 61674
rect 483020 61610 483072 61616
rect 482284 3664 482336 3670
rect 482284 3606 482336 3612
rect 482928 3664 482980 3670
rect 482928 3606 482980 3612
rect 481088 3256 481140 3262
rect 481088 3198 481140 3204
rect 481548 3256 481600 3262
rect 481548 3198 481600 3204
rect 479892 3052 479944 3058
rect 479892 2994 479944 3000
rect 478696 2984 478748 2990
rect 478696 2926 478748 2932
rect 478708 480 478736 2926
rect 479904 480 479932 2994
rect 481100 480 481128 3198
rect 482296 480 482324 3606
rect 483032 626 483060 61610
rect 483676 3058 483704 61746
rect 485240 60790 485268 64110
rect 485872 61600 485924 61606
rect 485872 61542 485924 61548
rect 485228 60784 485280 60790
rect 485228 60726 485280 60732
rect 485688 60784 485740 60790
rect 485688 60726 485740 60732
rect 485700 4962 485728 60726
rect 485688 4956 485740 4962
rect 485688 4898 485740 4904
rect 485780 3800 485832 3806
rect 485780 3742 485832 3748
rect 484584 3460 484636 3466
rect 484584 3402 484636 3408
rect 483664 3052 483716 3058
rect 483664 2994 483716 3000
rect 483032 598 483520 626
rect 483492 480 483520 598
rect 484596 480 484624 3402
rect 485792 480 485820 3742
rect 485884 610 485912 61542
rect 486252 60790 486280 64110
rect 487080 61878 487108 64110
rect 487068 61872 487120 61878
rect 487068 61814 487120 61820
rect 486240 60784 486292 60790
rect 486240 60726 486292 60732
rect 487068 60784 487120 60790
rect 487068 60726 487120 60732
rect 487080 3806 487108 60726
rect 488460 4894 488488 64110
rect 489288 60790 489316 64110
rect 490300 61810 490328 64110
rect 490288 61804 490340 61810
rect 490288 61746 490340 61752
rect 491220 61606 491248 64110
rect 491208 61600 491260 61606
rect 491208 61542 491260 61548
rect 489920 61464 489972 61470
rect 489920 61406 489972 61412
rect 489276 60784 489328 60790
rect 489276 60726 489328 60732
rect 489828 60784 489880 60790
rect 489828 60726 489880 60732
rect 488448 4888 488500 4894
rect 488448 4830 488500 4836
rect 489840 3874 489868 60726
rect 489368 3868 489420 3874
rect 489368 3810 489420 3816
rect 489828 3868 489880 3874
rect 489828 3810 489880 3816
rect 487068 3800 487120 3806
rect 487068 3742 487120 3748
rect 488172 3120 488224 3126
rect 488172 3062 488224 3068
rect 485872 604 485924 610
rect 485872 546 485924 552
rect 486976 604 487028 610
rect 486976 546 487028 552
rect 486988 480 487016 546
rect 488184 480 488212 3062
rect 489380 480 489408 3810
rect 489932 610 489960 61406
rect 492600 3466 492628 64110
rect 493336 60790 493364 64110
rect 494244 61396 494296 61402
rect 494244 61338 494296 61344
rect 493324 60784 493376 60790
rect 493324 60726 493376 60732
rect 493968 60784 494020 60790
rect 493968 60726 494020 60732
rect 492956 3596 493008 3602
rect 492956 3538 493008 3544
rect 492588 3460 492640 3466
rect 492588 3402 492640 3408
rect 491760 3392 491812 3398
rect 491760 3334 491812 3340
rect 489920 604 489972 610
rect 489920 546 489972 552
rect 490564 604 490616 610
rect 490564 546 490616 552
rect 490576 480 490604 546
rect 491772 480 491800 3334
rect 492968 480 492996 3538
rect 493980 3126 494008 60726
rect 493968 3120 494020 3126
rect 493968 3062 494020 3068
rect 494256 626 494284 61338
rect 494348 60790 494376 64110
rect 494336 60784 494388 60790
rect 494336 60726 494388 60732
rect 495256 60784 495308 60790
rect 495256 60726 495308 60732
rect 495268 4826 495296 60726
rect 495256 4820 495308 4826
rect 495256 4762 495308 4768
rect 495360 3602 495388 64110
rect 496084 62008 496136 62014
rect 496084 61950 496136 61956
rect 495348 3596 495400 3602
rect 495348 3538 495400 3544
rect 496096 3398 496124 61950
rect 496464 61674 496492 64110
rect 496452 61668 496504 61674
rect 496452 61610 496504 61616
rect 496820 61532 496872 61538
rect 496820 61474 496872 61480
rect 496084 3392 496136 3398
rect 496084 3334 496136 3340
rect 496544 3324 496596 3330
rect 496544 3266 496596 3272
rect 495348 3188 495400 3194
rect 495348 3130 495400 3136
rect 494164 598 494284 626
rect 494164 480 494192 598
rect 495360 480 495388 3130
rect 496556 480 496584 3266
rect 496832 610 496860 61474
rect 497476 61130 497504 64110
rect 497464 61124 497516 61130
rect 497464 61066 497516 61072
rect 498488 60790 498516 64110
rect 498476 60784 498528 60790
rect 498476 60726 498528 60732
rect 499408 3534 499436 64110
rect 499488 60784 499540 60790
rect 499488 60726 499540 60732
rect 498936 3528 498988 3534
rect 498936 3470 498988 3476
rect 499396 3528 499448 3534
rect 499396 3470 499448 3476
rect 496820 604 496872 610
rect 496820 546 496872 552
rect 497740 604 497792 610
rect 497740 546 497792 552
rect 497752 480 497780 546
rect 498948 480 498976 3470
rect 499500 3194 499528 60726
rect 500880 5098 500908 64110
rect 501524 60790 501552 64110
rect 502260 61402 502288 64110
rect 502248 61396 502300 61402
rect 502248 61338 502300 61344
rect 501604 61124 501656 61130
rect 501604 61066 501656 61072
rect 501512 60784 501564 60790
rect 501512 60726 501564 60732
rect 501616 5506 501644 61066
rect 503548 60858 503576 64110
rect 503536 60852 503588 60858
rect 503536 60794 503588 60800
rect 504560 60790 504588 64110
rect 505572 61470 505600 64110
rect 505560 61464 505612 61470
rect 505560 61406 505612 61412
rect 505744 60852 505796 60858
rect 505744 60794 505796 60800
rect 502248 60784 502300 60790
rect 502248 60726 502300 60732
rect 504548 60784 504600 60790
rect 504548 60726 504600 60732
rect 505008 60784 505060 60790
rect 505008 60726 505060 60732
rect 501604 5500 501656 5506
rect 501604 5442 501656 5448
rect 500868 5092 500920 5098
rect 500868 5034 500920 5040
rect 501236 5024 501288 5030
rect 501236 4966 501288 4972
rect 500132 3732 500184 3738
rect 500132 3674 500184 3680
rect 499488 3188 499540 3194
rect 499488 3130 499540 3136
rect 500144 480 500172 3674
rect 501248 480 501276 4966
rect 502260 3330 502288 60726
rect 504824 5296 504876 5302
rect 504824 5238 504876 5244
rect 502432 4004 502484 4010
rect 502432 3946 502484 3952
rect 502248 3324 502300 3330
rect 502248 3266 502300 3272
rect 502444 480 502472 3946
rect 503628 3052 503680 3058
rect 503628 2994 503680 3000
rect 503640 480 503668 2994
rect 504836 480 504864 5238
rect 505020 3738 505048 60726
rect 505756 5302 505784 60794
rect 506400 60790 506428 64110
rect 506388 60784 506440 60790
rect 506388 60726 506440 60732
rect 507124 60784 507176 60790
rect 507124 60726 507176 60732
rect 505744 5296 505796 5302
rect 505744 5238 505796 5244
rect 507136 5030 507164 60726
rect 507124 5024 507176 5030
rect 507124 4966 507176 4972
rect 507780 4078 507808 64110
rect 508504 61736 508556 61742
rect 508504 61678 508556 61684
rect 508412 5160 508464 5166
rect 508412 5102 508464 5108
rect 506020 4072 506072 4078
rect 506020 4014 506072 4020
rect 507768 4072 507820 4078
rect 507768 4014 507820 4020
rect 505008 3732 505060 3738
rect 505008 3674 505060 3680
rect 506032 480 506060 4014
rect 507308 4004 507360 4010
rect 507308 3946 507360 3952
rect 507320 3398 507348 3946
rect 507216 3392 507268 3398
rect 507216 3334 507268 3340
rect 507308 3392 507360 3398
rect 507308 3334 507360 3340
rect 507228 480 507256 3334
rect 508424 480 508452 5102
rect 508516 4146 508544 61678
rect 508700 61538 508728 64110
rect 508688 61532 508740 61538
rect 508688 61474 508740 61480
rect 509712 60790 509740 64110
rect 509700 60784 509752 60790
rect 509700 60726 509752 60732
rect 508504 4140 508556 4146
rect 508504 4082 508556 4088
rect 510540 4010 510568 64110
rect 511264 60784 511316 60790
rect 511264 60726 511316 60732
rect 511276 5166 511304 60726
rect 511264 5160 511316 5166
rect 511264 5102 511316 5108
rect 510804 4140 510856 4146
rect 510804 4082 510856 4088
rect 510528 4004 510580 4010
rect 510528 3946 510580 3952
rect 509608 3392 509660 3398
rect 509608 3334 509660 3340
rect 509620 480 509648 3334
rect 510816 480 510844 4082
rect 511920 3398 511948 64110
rect 512644 61940 512696 61946
rect 512644 61882 512696 61888
rect 512000 5228 512052 5234
rect 512000 5170 512052 5176
rect 511908 3392 511960 3398
rect 511908 3334 511960 3340
rect 512012 480 512040 5170
rect 512656 3058 512684 61882
rect 512748 60858 512776 64110
rect 512736 60852 512788 60858
rect 512736 60794 512788 60800
rect 513760 60790 513788 64110
rect 514680 61742 514708 64110
rect 515784 61946 515812 64110
rect 516796 62014 516824 64110
rect 517808 62082 517836 64110
rect 517796 62076 517848 62082
rect 517796 62018 517848 62024
rect 516784 62008 516836 62014
rect 516784 61950 516836 61956
rect 515772 61940 515824 61946
rect 515772 61882 515824 61888
rect 516876 61872 516928 61878
rect 516876 61814 516928 61820
rect 514668 61736 514720 61742
rect 514668 61678 514720 61684
rect 515404 60852 515456 60858
rect 515404 60794 515456 60800
rect 513748 60784 513800 60790
rect 513748 60726 513800 60732
rect 514668 60784 514720 60790
rect 514668 60726 514720 60732
rect 514680 4146 514708 60726
rect 515416 5234 515444 60794
rect 516888 51202 516916 61814
rect 516876 51196 516928 51202
rect 516876 51138 516928 51144
rect 516968 51060 517020 51066
rect 516968 51002 517020 51008
rect 516980 48362 517008 51002
rect 516888 48334 517008 48362
rect 516888 48278 516916 48334
rect 516692 48272 516744 48278
rect 516692 48214 516744 48220
rect 516876 48272 516928 48278
rect 516876 48214 516928 48220
rect 516704 31754 516732 48214
rect 516692 31748 516744 31754
rect 516692 31690 516744 31696
rect 516876 31748 516928 31754
rect 516876 31690 516928 31696
rect 516888 28966 516916 31690
rect 516600 28960 516652 28966
rect 516600 28902 516652 28908
rect 516876 28960 516928 28966
rect 516876 28902 516928 28908
rect 516612 19378 516640 28902
rect 516600 19372 516652 19378
rect 516600 19314 516652 19320
rect 516784 19372 516836 19378
rect 516784 19314 516836 19320
rect 516796 12458 516824 19314
rect 516796 12430 517008 12458
rect 515588 5364 515640 5370
rect 515588 5306 515640 5312
rect 515404 5228 515456 5234
rect 515404 5170 515456 5176
rect 514668 4140 514720 4146
rect 514668 4082 514720 4088
rect 514852 4004 514904 4010
rect 514852 3946 514904 3952
rect 513196 3936 513248 3942
rect 513196 3878 513248 3884
rect 512644 3052 512696 3058
rect 512644 2994 512696 3000
rect 513208 480 513236 3878
rect 514484 3800 514536 3806
rect 514484 3742 514536 3748
rect 514496 3262 514524 3742
rect 514392 3256 514444 3262
rect 514392 3198 514444 3204
rect 514484 3256 514536 3262
rect 514484 3198 514536 3204
rect 514404 480 514432 3198
rect 514864 2922 514892 3946
rect 514852 2916 514904 2922
rect 514852 2858 514904 2864
rect 515600 480 515628 5306
rect 516980 4078 517008 12430
rect 518728 6254 518756 64110
rect 518808 62076 518860 62082
rect 518808 62018 518860 62024
rect 518716 6248 518768 6254
rect 518716 6190 518768 6196
rect 516876 4072 516928 4078
rect 516876 4014 516928 4020
rect 516968 4072 517020 4078
rect 516968 4014 517020 4020
rect 516784 3664 516836 3670
rect 516784 3606 516836 3612
rect 516796 480 516824 3606
rect 516888 2990 516916 4014
rect 518820 3942 518848 62018
rect 519544 62008 519596 62014
rect 519544 61950 519596 61956
rect 519556 10554 519584 61950
rect 519924 60858 519952 64110
rect 520832 61804 520884 61810
rect 520832 61746 520884 61752
rect 519912 60852 519964 60858
rect 519912 60794 519964 60800
rect 520844 60722 520872 61746
rect 520936 61266 520964 64110
rect 521948 62082 521976 64110
rect 521936 62076 521988 62082
rect 521936 62018 521988 62024
rect 522856 62076 522908 62082
rect 522856 62018 522908 62024
rect 522304 61940 522356 61946
rect 522304 61882 522356 61888
rect 520924 61260 520976 61266
rect 520924 61202 520976 61208
rect 521568 61260 521620 61266
rect 521568 61202 521620 61208
rect 520832 60716 520884 60722
rect 520832 60658 520884 60664
rect 520924 60648 520976 60654
rect 520924 60590 520976 60596
rect 520936 53174 520964 60590
rect 520740 53168 520792 53174
rect 520740 53110 520792 53116
rect 520924 53168 520976 53174
rect 520924 53110 520976 53116
rect 520752 48346 520780 53110
rect 520740 48340 520792 48346
rect 520740 48282 520792 48288
rect 520924 48340 520976 48346
rect 520924 48282 520976 48288
rect 520936 38706 520964 48282
rect 520936 38678 521056 38706
rect 521028 31822 521056 38678
rect 521016 31816 521068 31822
rect 521016 31758 521068 31764
rect 521016 31680 521068 31686
rect 521016 31622 521068 31628
rect 521028 28966 521056 31622
rect 520924 28960 520976 28966
rect 520924 28902 520976 28908
rect 521016 28960 521068 28966
rect 521016 28902 521068 28908
rect 520936 12458 520964 28902
rect 520936 12430 521148 12458
rect 519464 10526 519584 10554
rect 519084 4956 519136 4962
rect 519084 4898 519136 4904
rect 518808 3936 518860 3942
rect 518808 3878 518860 3884
rect 517888 3052 517940 3058
rect 517888 2994 517940 3000
rect 516876 2984 516928 2990
rect 516876 2926 516928 2932
rect 517900 480 517928 2994
rect 519096 480 519124 4898
rect 519464 3670 519492 10526
rect 519452 3664 519504 3670
rect 519452 3606 519504 3612
rect 520372 3664 520424 3670
rect 520372 3606 520424 3612
rect 520384 3262 520412 3606
rect 520280 3256 520332 3262
rect 520280 3198 520332 3204
rect 520372 3256 520424 3262
rect 520372 3198 520424 3204
rect 520292 480 520320 3198
rect 521120 3058 521148 12430
rect 521476 4072 521528 4078
rect 521476 4014 521528 4020
rect 521108 3052 521160 3058
rect 521108 2994 521160 3000
rect 521488 480 521516 4014
rect 521580 3806 521608 61202
rect 522316 5370 522344 61882
rect 522304 5364 522356 5370
rect 522304 5306 522356 5312
rect 522868 4894 522896 62018
rect 522672 4888 522724 4894
rect 522672 4830 522724 4836
rect 522856 4888 522908 4894
rect 522856 4830 522908 4836
rect 521568 3800 521620 3806
rect 521568 3742 521620 3748
rect 522684 480 522712 4830
rect 522960 3670 522988 64110
rect 524340 3874 524368 64110
rect 524984 62014 525012 64110
rect 524972 62008 525024 62014
rect 524972 61950 525024 61956
rect 525720 61878 525748 64110
rect 525708 61872 525760 61878
rect 525708 61814 525760 61820
rect 527008 61810 527036 64110
rect 526996 61804 527048 61810
rect 526996 61746 527048 61752
rect 525800 61600 525852 61606
rect 525800 61542 525852 61548
rect 523868 3868 523920 3874
rect 523868 3810 523920 3816
rect 524328 3868 524380 3874
rect 524328 3810 524380 3816
rect 522948 3664 523000 3670
rect 522948 3606 523000 3612
rect 523880 480 523908 3810
rect 525064 3052 525116 3058
rect 525064 2994 525116 3000
rect 525076 480 525104 2994
rect 525812 610 525840 61542
rect 526444 60852 526496 60858
rect 526444 60794 526496 60800
rect 526456 3058 526484 60794
rect 528020 60790 528048 64110
rect 529032 60926 529060 64110
rect 529204 61668 529256 61674
rect 529204 61610 529256 61616
rect 529020 60920 529072 60926
rect 529020 60862 529072 60868
rect 528008 60784 528060 60790
rect 528008 60726 528060 60732
rect 528468 60784 528520 60790
rect 528468 60726 528520 60732
rect 528480 6186 528508 60726
rect 528468 6180 528520 6186
rect 528468 6122 528520 6128
rect 528468 4072 528520 4078
rect 528468 4014 528520 4020
rect 528376 4004 528428 4010
rect 528376 3946 528428 3952
rect 527456 3460 527508 3466
rect 527456 3402 527508 3408
rect 526444 3052 526496 3058
rect 526444 2994 526496 3000
rect 525800 604 525852 610
rect 525800 546 525852 552
rect 526260 604 526312 610
rect 526260 546 526312 552
rect 526272 480 526300 546
rect 527468 480 527496 3402
rect 528388 2922 528416 3946
rect 528480 2990 528508 4014
rect 528652 3120 528704 3126
rect 528652 3062 528704 3068
rect 528468 2984 528520 2990
rect 528468 2926 528520 2932
rect 528376 2916 528428 2922
rect 528376 2858 528428 2864
rect 528664 480 528692 3062
rect 529216 2922 529244 61610
rect 529860 5114 529888 64110
rect 531148 60858 531176 64110
rect 531964 62008 532016 62014
rect 531964 61950 532016 61956
rect 531136 60852 531188 60858
rect 531136 60794 531188 60800
rect 531976 5438 532004 61950
rect 532160 60790 532188 64110
rect 533172 61674 533200 64110
rect 533160 61668 533212 61674
rect 533160 61610 533212 61616
rect 533344 60852 533396 60858
rect 533344 60794 533396 60800
rect 532148 60784 532200 60790
rect 532148 60726 532200 60732
rect 532608 60784 532660 60790
rect 532608 60726 532660 60732
rect 531964 5432 532016 5438
rect 531964 5374 532016 5380
rect 529676 5086 529888 5114
rect 529676 3466 529704 5086
rect 529848 4820 529900 4826
rect 529848 4762 529900 4768
rect 529664 3460 529716 3466
rect 529664 3402 529716 3408
rect 529204 2916 529256 2922
rect 529204 2858 529256 2864
rect 529860 480 529888 4762
rect 532620 3602 532648 60726
rect 533356 4962 533384 60794
rect 534000 60790 534028 64110
rect 534724 61872 534776 61878
rect 534724 61814 534776 61820
rect 533988 60784 534040 60790
rect 533988 60726 534040 60732
rect 533436 5500 533488 5506
rect 533436 5442 533488 5448
rect 533344 4956 533396 4962
rect 533344 4898 533396 4904
rect 531044 3596 531096 3602
rect 531044 3538 531096 3544
rect 532608 3596 532660 3602
rect 532608 3538 532660 3544
rect 531056 480 531084 3538
rect 532240 2916 532292 2922
rect 532240 2858 532292 2864
rect 532252 480 532280 2858
rect 533448 480 533476 5442
rect 534540 3188 534592 3194
rect 534540 3130 534592 3136
rect 534552 480 534580 3130
rect 534736 3126 534764 61814
rect 535196 61062 535224 64110
rect 535184 61056 535236 61062
rect 535184 60998 535236 61004
rect 536208 60790 536236 64110
rect 537220 61606 537248 64110
rect 538048 61878 538076 64110
rect 538036 61872 538088 61878
rect 538036 61814 538088 61820
rect 537208 61600 537260 61606
rect 537208 61542 537260 61548
rect 537484 60920 537536 60926
rect 537484 60862 537536 60868
rect 536104 60784 536156 60790
rect 536104 60726 536156 60732
rect 536196 60784 536248 60790
rect 536196 60726 536248 60732
rect 536748 60784 536800 60790
rect 536748 60726 536800 60732
rect 536116 4826 536144 60726
rect 536104 4820 536156 4826
rect 536104 4762 536156 4768
rect 536760 3534 536788 60726
rect 536932 5092 536984 5098
rect 536932 5034 536984 5040
rect 535736 3528 535788 3534
rect 535736 3470 535788 3476
rect 536748 3528 536800 3534
rect 536748 3470 536800 3476
rect 534724 3120 534776 3126
rect 534724 3062 534776 3068
rect 535748 480 535776 3470
rect 536944 480 536972 5034
rect 537496 3194 537524 60862
rect 538232 22098 538260 683318
rect 538876 218006 538904 686394
rect 538968 264926 538996 686462
rect 539060 311846 539088 686598
rect 539140 683732 539192 683738
rect 539140 683674 539192 683680
rect 539152 358766 539180 683674
rect 539232 683596 539284 683602
rect 539232 683538 539284 683544
rect 539244 369850 539272 683538
rect 539336 452606 539364 686870
rect 540336 686860 540388 686866
rect 540336 686802 540388 686808
rect 539508 685568 539560 685574
rect 539508 685510 539560 685516
rect 539416 685364 539468 685370
rect 539416 685306 539468 685312
rect 539428 487150 539456 685306
rect 539520 534070 539548 685510
rect 540242 684584 540298 684593
rect 540242 684519 540298 684528
rect 539508 534064 539560 534070
rect 539508 534006 539560 534012
rect 539416 487144 539468 487150
rect 539416 487086 539468 487092
rect 539324 452600 539376 452606
rect 539324 452542 539376 452548
rect 539232 369844 539284 369850
rect 539232 369786 539284 369792
rect 539140 358760 539192 358766
rect 539140 358702 539192 358708
rect 539048 311840 539100 311846
rect 539048 311782 539100 311788
rect 538956 264920 539008 264926
rect 538956 264862 539008 264868
rect 538864 218000 538916 218006
rect 538864 217942 538916 217948
rect 540256 64870 540284 684519
rect 540348 463690 540376 686802
rect 541716 686792 541768 686798
rect 541716 686734 541768 686740
rect 540888 685840 540940 685846
rect 540888 685782 540940 685788
rect 540704 685772 540756 685778
rect 540704 685714 540756 685720
rect 540520 685704 540572 685710
rect 540520 685646 540572 685652
rect 540426 684856 540482 684865
rect 540426 684791 540482 684800
rect 540336 463684 540388 463690
rect 540336 463626 540388 463632
rect 540440 111790 540468 684791
rect 540532 580990 540560 685646
rect 540610 684992 540666 685001
rect 540610 684927 540666 684936
rect 540520 580984 540572 580990
rect 540520 580926 540572 580932
rect 540624 158710 540652 684927
rect 540716 627910 540744 685714
rect 540794 685400 540850 685409
rect 540794 685335 540850 685344
rect 540704 627904 540756 627910
rect 540704 627846 540756 627852
rect 540808 299470 540836 685335
rect 540900 674830 540928 685782
rect 541624 684956 541676 684962
rect 541624 684898 541676 684904
rect 540888 674824 540940 674830
rect 540888 674766 540940 674772
rect 541636 393310 541664 684898
rect 541728 405686 541756 686734
rect 577780 686248 577832 686254
rect 577780 686190 577832 686196
rect 577502 686080 577558 686089
rect 577502 686015 577558 686024
rect 577688 686044 577740 686050
rect 543096 684480 543148 684486
rect 543096 684422 543148 684428
rect 543004 684276 543056 684282
rect 543004 684218 543056 684224
rect 541808 684140 541860 684146
rect 541808 684082 541860 684088
rect 541820 546446 541848 684082
rect 543016 593366 543044 684218
rect 543108 640286 543136 684422
rect 543096 640280 543148 640286
rect 543096 640222 543148 640228
rect 543004 593360 543056 593366
rect 543004 593302 543056 593308
rect 541808 546440 541860 546446
rect 541808 546382 541860 546388
rect 541716 405680 541768 405686
rect 541716 405622 541768 405628
rect 541624 393304 541676 393310
rect 541624 393246 541676 393252
rect 540796 299464 540848 299470
rect 540796 299406 540848 299412
rect 540612 158704 540664 158710
rect 540612 158646 540664 158652
rect 540428 111784 540480 111790
rect 540428 111726 540480 111732
rect 540244 64864 540296 64870
rect 540244 64806 540296 64812
rect 538936 64110 539272 64138
rect 539244 61402 539272 64110
rect 541624 61872 541676 61878
rect 541624 61814 541676 61820
rect 538312 61396 538364 61402
rect 538312 61338 538364 61344
rect 539232 61396 539284 61402
rect 539232 61338 539284 61344
rect 538220 22092 538272 22098
rect 538220 22034 538272 22040
rect 538128 3324 538180 3330
rect 538128 3266 538180 3272
rect 537484 3188 537536 3194
rect 537484 3130 537536 3136
rect 538140 480 538168 3266
rect 538324 610 538352 61338
rect 540244 61056 540296 61062
rect 540244 60998 540296 61004
rect 540256 2990 540284 60998
rect 540520 5296 540572 5302
rect 540520 5238 540572 5244
rect 540244 2984 540296 2990
rect 540244 2926 540296 2932
rect 538312 604 538364 610
rect 538312 546 538364 552
rect 539324 604 539376 610
rect 539324 546 539376 552
rect 539336 480 539364 546
rect 540532 480 540560 5238
rect 541636 2922 541664 61814
rect 547236 61804 547288 61810
rect 547236 61746 547288 61752
rect 545764 61736 545816 61742
rect 545764 61678 545816 61684
rect 544384 61532 544436 61538
rect 544384 61474 544436 61480
rect 542360 61464 542412 61470
rect 542360 61406 542412 61412
rect 541716 3732 541768 3738
rect 541716 3674 541768 3680
rect 541624 2916 541676 2922
rect 541624 2858 541676 2864
rect 541728 480 541756 3674
rect 542372 610 542400 61406
rect 544108 5024 544160 5030
rect 544108 4966 544160 4972
rect 543004 4004 543056 4010
rect 543004 3946 543056 3952
rect 543016 3738 543044 3946
rect 543004 3732 543056 3738
rect 543004 3674 543056 3680
rect 542360 604 542412 610
rect 542360 546 542412 552
rect 542912 604 542964 610
rect 542912 546 542964 552
rect 542924 480 542952 546
rect 544120 480 544148 4966
rect 544396 3330 544424 61474
rect 545304 4072 545356 4078
rect 545304 4014 545356 4020
rect 544384 3324 544436 3330
rect 544384 3266 544436 3272
rect 545316 480 545344 4014
rect 545776 2854 545804 61678
rect 547144 61668 547196 61674
rect 547144 61610 547196 61616
rect 547156 4078 547184 61610
rect 547144 4072 547196 4078
rect 547144 4014 547196 4020
rect 546500 3324 546552 3330
rect 546500 3266 546552 3272
rect 546592 3324 546644 3330
rect 546592 3266 546644 3272
rect 545764 2848 545816 2854
rect 545764 2790 545816 2796
rect 546512 480 546540 3266
rect 546604 2990 546632 3266
rect 546592 2984 546644 2990
rect 546592 2926 546644 2932
rect 547248 2922 547276 61746
rect 567844 61600 567896 61606
rect 567844 61542 567896 61548
rect 548524 61396 548576 61402
rect 548524 61338 548576 61344
rect 547696 5160 547748 5166
rect 547696 5102 547748 5108
rect 547236 2916 547288 2922
rect 547236 2858 547288 2864
rect 547708 480 547736 5102
rect 548536 4010 548564 61338
rect 558368 6248 558420 6254
rect 558368 6190 558420 6196
rect 554780 5364 554832 5370
rect 554780 5306 554832 5312
rect 551192 5228 551244 5234
rect 551192 5170 551244 5176
rect 548524 4004 548576 4010
rect 548524 3946 548576 3952
rect 548892 3732 548944 3738
rect 548892 3674 548944 3680
rect 548904 480 548932 3674
rect 550088 3392 550140 3398
rect 550088 3334 550140 3340
rect 550100 480 550128 3334
rect 551204 480 551232 5170
rect 552388 4140 552440 4146
rect 552388 4082 552440 4088
rect 552400 480 552428 4082
rect 552664 3732 552716 3738
rect 552664 3674 552716 3680
rect 552676 2990 552704 3674
rect 552664 2984 552716 2990
rect 552664 2926 552716 2932
rect 553584 2848 553636 2854
rect 553584 2790 553636 2796
rect 553596 480 553624 2790
rect 554792 480 554820 5306
rect 557172 3936 557224 3942
rect 557172 3878 557224 3884
rect 555976 3256 556028 3262
rect 555976 3198 556028 3204
rect 555988 480 556016 3198
rect 557184 480 557212 3878
rect 558380 480 558408 6190
rect 565544 5432 565596 5438
rect 565544 5374 565596 5380
rect 561956 4888 562008 4894
rect 561956 4830 562008 4836
rect 560760 3800 560812 3806
rect 560760 3742 560812 3748
rect 559564 3052 559616 3058
rect 559564 2994 559616 3000
rect 559576 480 559604 2994
rect 560772 480 560800 3742
rect 561968 480 561996 4830
rect 564348 3868 564400 3874
rect 564348 3810 564400 3816
rect 563152 3664 563204 3670
rect 563152 3606 563204 3612
rect 563164 480 563192 3606
rect 564360 480 564388 3810
rect 565556 480 565584 5374
rect 567856 3670 567884 61542
rect 577516 41410 577544 686015
rect 577688 685986 577740 685992
rect 577596 685908 577648 685914
rect 577596 685850 577648 685856
rect 577608 205630 577636 685850
rect 577700 252550 577728 685986
rect 577792 346390 577820 686190
rect 578148 685500 578200 685506
rect 578148 685442 578200 685448
rect 578056 685296 578108 685302
rect 578056 685238 578108 685244
rect 577964 685160 578016 685166
rect 577964 685102 578016 685108
rect 577872 684684 577924 684690
rect 577872 684626 577924 684632
rect 577884 440230 577912 684626
rect 577976 557394 578004 685102
rect 578068 604450 578096 685238
rect 578160 651370 578188 685442
rect 579988 685228 580040 685234
rect 579988 685170 580040 685176
rect 579804 684888 579856 684894
rect 579804 684830 579856 684836
rect 579712 674824 579764 674830
rect 579712 674766 579764 674772
rect 579724 674665 579752 674766
rect 579710 674656 579766 674665
rect 579710 674591 579766 674600
rect 578148 651364 578200 651370
rect 578148 651306 578200 651312
rect 579620 651364 579672 651370
rect 579620 651306 579672 651312
rect 579632 651137 579660 651306
rect 579618 651128 579674 651137
rect 579618 651063 579674 651072
rect 579712 640280 579764 640286
rect 579712 640222 579764 640228
rect 579724 639441 579752 640222
rect 579710 639432 579766 639441
rect 579710 639367 579766 639376
rect 579712 627904 579764 627910
rect 579712 627846 579764 627852
rect 579724 627745 579752 627846
rect 579710 627736 579766 627745
rect 579710 627671 579766 627680
rect 578056 604444 578108 604450
rect 578056 604386 578108 604392
rect 579620 604444 579672 604450
rect 579620 604386 579672 604392
rect 579632 604217 579660 604386
rect 579618 604208 579674 604217
rect 579618 604143 579674 604152
rect 579712 593360 579764 593366
rect 579712 593302 579764 593308
rect 579724 592521 579752 593302
rect 579710 592512 579766 592521
rect 579710 592447 579766 592456
rect 579712 580984 579764 580990
rect 579712 580926 579764 580932
rect 579724 580825 579752 580926
rect 579710 580816 579766 580825
rect 579710 580751 579766 580760
rect 577964 557388 578016 557394
rect 577964 557330 578016 557336
rect 579620 557388 579672 557394
rect 579620 557330 579672 557336
rect 579632 557297 579660 557330
rect 579618 557288 579674 557297
rect 579618 557223 579674 557232
rect 579712 546440 579764 546446
rect 579712 546382 579764 546388
rect 579724 545601 579752 546382
rect 579710 545592 579766 545601
rect 579710 545527 579766 545536
rect 579712 534064 579764 534070
rect 579712 534006 579764 534012
rect 579724 533905 579752 534006
rect 579710 533896 579766 533905
rect 579710 533831 579766 533840
rect 579816 510377 579844 684830
rect 579896 683664 579948 683670
rect 579896 683606 579948 683612
rect 579802 510368 579858 510377
rect 579802 510303 579858 510312
rect 579908 498681 579936 683606
rect 579894 498672 579950 498681
rect 579894 498607 579950 498616
rect 579896 487144 579948 487150
rect 579896 487086 579948 487092
rect 579908 486849 579936 487086
rect 579894 486840 579950 486849
rect 579894 486775 579950 486784
rect 579896 463684 579948 463690
rect 579896 463626 579948 463632
rect 579908 463457 579936 463626
rect 579894 463448 579950 463457
rect 579894 463383 579950 463392
rect 579896 452600 579948 452606
rect 579896 452542 579948 452548
rect 579908 451761 579936 452542
rect 579894 451752 579950 451761
rect 579894 451687 579950 451696
rect 577872 440224 577924 440230
rect 577872 440166 577924 440172
rect 579896 440224 579948 440230
rect 579896 440166 579948 440172
rect 579908 439929 579936 440166
rect 579894 439920 579950 439929
rect 579894 439855 579950 439864
rect 580000 416537 580028 685170
rect 579986 416528 580042 416537
rect 579986 416463 580042 416472
rect 579988 405680 580040 405686
rect 579988 405622 580040 405628
rect 580000 404841 580028 405622
rect 579986 404832 580042 404841
rect 579986 404767 580042 404776
rect 579988 393304 580040 393310
rect 579988 393246 580040 393252
rect 580000 393009 580028 393246
rect 579986 393000 580042 393009
rect 579986 392935 580042 392944
rect 579988 369844 580040 369850
rect 579988 369786 580040 369792
rect 580000 369617 580028 369786
rect 579986 369608 580042 369617
rect 579986 369543 580042 369552
rect 579988 358760 580040 358766
rect 579988 358702 580040 358708
rect 580000 357921 580028 358702
rect 579986 357912 580042 357921
rect 579986 357847 580042 357856
rect 577780 346384 577832 346390
rect 577780 346326 577832 346332
rect 579896 346384 579948 346390
rect 579896 346326 579948 346332
rect 579908 346089 579936 346326
rect 579894 346080 579950 346089
rect 579894 346015 579950 346024
rect 577688 252544 577740 252550
rect 577688 252486 577740 252492
rect 579988 252544 580040 252550
rect 579988 252486 580040 252492
rect 580000 252249 580028 252486
rect 579986 252240 580042 252249
rect 579986 252175 580042 252184
rect 577596 205624 577648 205630
rect 577596 205566 577648 205572
rect 580092 181937 580120 686967
rect 580172 686938 580224 686944
rect 580184 686361 580212 686938
rect 580630 686760 580686 686769
rect 580630 686695 580686 686704
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 580446 686080 580502 686089
rect 580446 686015 580502 686024
rect 580262 685944 580318 685953
rect 580262 685879 580318 685888
rect 580172 683868 580224 683874
rect 580172 683810 580224 683816
rect 580184 322697 580212 683810
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 580172 311840 580224 311846
rect 580172 311782 580224 311788
rect 580184 310865 580212 311782
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 299169 580212 299406
rect 580170 299160 580226 299169
rect 580170 299095 580226 299104
rect 580172 264920 580224 264926
rect 580172 264862 580224 264868
rect 580184 263945 580212 264862
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 580078 181928 580134 181937
rect 580078 181863 580134 181872
rect 580172 158704 580224 158710
rect 580172 158646 580224 158652
rect 580184 158409 580212 158646
rect 580170 158400 580226 158409
rect 580170 158335 580226 158344
rect 580172 111784 580224 111790
rect 580172 111726 580224 111732
rect 580184 111489 580212 111726
rect 580170 111480 580226 111489
rect 580170 111415 580226 111424
rect 580172 64864 580224 64870
rect 580172 64806 580224 64812
rect 580184 64569 580212 64806
rect 580170 64560 580226 64569
rect 580170 64495 580226 64504
rect 577504 41404 577556 41410
rect 577504 41346 577556 41352
rect 579896 30320 579948 30326
rect 579896 30262 579948 30268
rect 579908 29345 579936 30262
rect 579894 29336 579950 29345
rect 579894 29271 579950 29280
rect 580276 17649 580304 685879
rect 580354 685536 580410 685545
rect 580354 685471 580410 685480
rect 580368 76265 580396 685471
rect 580460 87961 580488 686015
rect 580540 683188 580592 683194
rect 580540 683130 580592 683136
rect 580552 170105 580580 683130
rect 580538 170096 580594 170105
rect 580538 170031 580594 170040
rect 580644 123185 580672 686695
rect 580814 686488 580870 686497
rect 580814 686423 580870 686432
rect 580724 683256 580776 683262
rect 580724 683198 580776 683204
rect 580736 228857 580764 683198
rect 580722 228848 580778 228857
rect 580722 228783 580778 228792
rect 580724 205624 580776 205630
rect 580724 205566 580776 205572
rect 580736 205329 580764 205566
rect 580722 205320 580778 205329
rect 580722 205255 580778 205264
rect 580828 134881 580856 686423
rect 580908 684344 580960 684350
rect 580908 684286 580960 684292
rect 580920 275777 580948 684286
rect 580906 275768 580962 275777
rect 580906 275703 580962 275712
rect 580814 134872 580870 134881
rect 580814 134807 580870 134816
rect 580630 123176 580686 123185
rect 580630 123111 580686 123120
rect 580446 87952 580502 87961
rect 580446 87887 580502 87896
rect 580354 76256 580410 76265
rect 580354 76191 580410 76200
rect 580540 41404 580592 41410
rect 580540 41346 580592 41352
rect 580552 41041 580580 41346
rect 580538 41032 580594 41041
rect 580538 40967 580594 40976
rect 580262 17640 580318 17649
rect 580262 17575 580318 17584
rect 569040 6180 569092 6186
rect 569040 6122 569092 6128
rect 567844 3664 567896 3670
rect 567844 3606 567896 3612
rect 566740 3120 566792 3126
rect 566740 3062 566792 3068
rect 566752 480 566780 3062
rect 567844 2984 567896 2990
rect 567844 2926 567896 2932
rect 567856 480 567884 2926
rect 569052 480 569080 6122
rect 572628 4956 572680 4962
rect 572628 4898 572680 4904
rect 571432 3460 571484 3466
rect 571432 3402 571484 3408
rect 570236 3188 570288 3194
rect 570236 3130 570288 3136
rect 570248 480 570276 3130
rect 571444 480 571472 3402
rect 572640 480 572668 4898
rect 576216 4820 576268 4826
rect 576216 4762 576268 4768
rect 575020 4072 575072 4078
rect 575020 4014 575072 4020
rect 573824 3596 573876 3602
rect 573824 3538 573876 3544
rect 573836 480 573864 3538
rect 575032 480 575060 4014
rect 576228 480 576256 4762
rect 582196 4004 582248 4010
rect 582196 3946 582248 3952
rect 581000 3732 581052 3738
rect 581000 3674 581052 3680
rect 579804 3664 579856 3670
rect 579804 3606 579856 3612
rect 578608 3528 578660 3534
rect 578608 3470 578660 3476
rect 577412 3324 577464 3330
rect 577412 3266 577464 3272
rect 577424 480 577452 3266
rect 578620 480 578648 3470
rect 579816 480 579844 3606
rect 581012 480 581040 3674
rect 582208 480 582236 3946
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 4802 687112 4858 687168
rect 3698 686840 3754 686896
rect 2778 682252 2780 682272
rect 2780 682252 2832 682272
rect 2832 682252 2834 682272
rect 2778 682216 2834 682252
rect 2778 667936 2834 667992
rect 2778 653520 2834 653576
rect 2778 624860 2780 624880
rect 2780 624860 2832 624880
rect 2832 624860 2834 624880
rect 2778 624824 2834 624860
rect 2778 610444 2780 610464
rect 2780 610444 2832 610464
rect 2832 610444 2834 610464
rect 2778 610408 2834 610444
rect 2778 595992 2834 596048
rect 2778 567332 2780 567352
rect 2780 567332 2832 567352
rect 2832 567332 2834 567352
rect 2778 567296 2834 567332
rect 2778 553016 2834 553072
rect 2778 538600 2834 538656
rect 2778 509940 2780 509960
rect 2780 509940 2832 509960
rect 2832 509940 2834 509960
rect 2778 509904 2834 509940
rect 2870 495488 2926 495544
rect 2870 481072 2926 481128
rect 2870 452412 2872 452432
rect 2872 452412 2924 452432
rect 2924 452412 2926 452432
rect 2870 452376 2926 452412
rect 2778 437960 2834 438016
rect 2870 423680 2926 423736
rect 2870 395020 2872 395040
rect 2872 395020 2924 395040
rect 2924 395020 2926 395040
rect 2870 394984 2926 395020
rect 2962 380568 3018 380624
rect 2962 366152 3018 366208
rect 2962 337456 3018 337512
rect 2962 323076 2964 323096
rect 2964 323076 3016 323096
rect 3016 323076 3018 323096
rect 2962 323040 3018 323076
rect 3514 686160 3570 686216
rect 3054 308760 3110 308816
rect 3054 294344 3110 294400
rect 3146 280064 3202 280120
rect 3238 265648 3294 265704
rect 3146 251268 3148 251288
rect 3148 251268 3200 251288
rect 3200 251268 3202 251288
rect 3146 251232 3202 251268
rect 3422 683712 3478 683768
rect 3330 236952 3386 237008
rect 3330 222536 3386 222592
rect 2778 208156 2780 208176
rect 2780 208156 2832 208176
rect 2832 208156 2834 208176
rect 2778 208120 2834 208156
rect 2778 179460 2780 179480
rect 2780 179460 2832 179480
rect 2832 179460 2834 179480
rect 2778 179424 2834 179460
rect 3146 165008 3202 165064
rect 3330 136312 3386 136368
rect 3330 122032 3386 122088
rect 3330 78920 3386 78976
rect 3606 683440 3662 683496
rect 3882 686568 3938 686624
rect 3790 683304 3846 683360
rect 3698 93200 3754 93256
rect 3974 683576 4030 683632
rect 4066 193840 4122 193896
rect 84198 686976 84254 687032
rect 6182 685072 6238 685128
rect 6826 683712 6882 683768
rect 6826 683168 6882 683224
rect 57978 686296 58034 686352
rect 45558 686024 45614 686080
rect 41418 685888 41474 685944
rect 39394 685208 39450 685264
rect 24122 684664 24178 684720
rect 22742 683848 22798 683904
rect 16578 683712 16634 683768
rect 16578 683168 16634 683224
rect 3974 150728 4030 150784
rect 35806 683712 35862 683768
rect 35806 683168 35862 683224
rect 39302 683712 39358 683768
rect 3882 107616 3938 107672
rect 3790 64504 3846 64560
rect 3606 50088 3662 50144
rect 3514 35808 3570 35864
rect 3514 21392 3570 21448
rect 3422 7112 3478 7168
rect 55126 684528 55182 684584
rect 75918 686704 75974 686760
rect 71778 686432 71834 686488
rect 68282 684800 68338 684856
rect 81346 684936 81402 684992
rect 120906 685344 120962 685400
rect 233238 685480 233294 685536
rect 277306 684256 277362 684312
rect 276938 683984 276994 684040
rect 280618 683984 280674 684040
rect 298190 684256 298246 684312
rect 298098 684120 298154 684176
rect 302146 684256 302202 684312
rect 302238 684120 302294 684176
rect 312450 684120 312506 684176
rect 311162 683984 311218 684040
rect 313002 683984 313058 684040
rect 318798 684120 318854 684176
rect 328366 684120 328422 684176
rect 328458 683984 328514 684040
rect 333242 684120 333298 684176
rect 331218 683712 331274 683768
rect 331402 683712 331458 683768
rect 331218 683576 331274 683632
rect 331402 683576 331458 683632
rect 331218 683440 331274 683496
rect 331402 683440 331458 683496
rect 333426 683984 333482 684040
rect 580170 697992 580226 698048
rect 356610 684936 356666 684992
rect 357346 684936 357402 684992
rect 356978 684800 357034 684856
rect 357346 684800 357402 684856
rect 357162 684664 357218 684720
rect 357346 684664 357402 684720
rect 357346 684392 357402 684448
rect 357346 684120 357402 684176
rect 360106 684256 360162 684312
rect 360106 683984 360162 684040
rect 367006 684256 367062 684312
rect 367006 683984 367062 684040
rect 379334 684256 379390 684312
rect 480258 687112 480314 687168
rect 386326 684256 386382 684312
rect 398746 684256 398802 684312
rect 405646 684256 405702 684312
rect 418066 684256 418122 684312
rect 424966 684256 425022 684312
rect 437386 684256 437442 684312
rect 444286 684256 444342 684312
rect 462318 685072 462374 685128
rect 456706 684256 456762 684312
rect 463606 684256 463662 684312
rect 476026 684256 476082 684312
rect 580078 686976 580134 687032
rect 506570 686840 506626 686896
rect 482926 684256 482982 684312
rect 488630 685208 488686 685264
rect 501786 684664 501842 684720
rect 495346 684256 495402 684312
rect 493046 683848 493102 683904
rect 510618 686568 510674 686624
rect 509238 683848 509294 683904
rect 528098 686160 528154 686216
rect 514942 683712 514998 683768
rect 497462 683576 497518 683632
rect 497922 683576 497978 683632
rect 509238 683576 509294 683632
rect 532698 683576 532754 683632
rect 519358 683440 519414 683496
rect 276938 683304 276994 683360
rect 277306 683304 277362 683360
rect 280618 683304 280674 683360
rect 311162 683304 311218 683360
rect 312450 683304 312506 683360
rect 313002 683304 313058 683360
rect 318798 683304 318854 683360
rect 333242 683304 333298 683360
rect 333426 683304 333482 683360
rect 521658 683324 521714 683360
rect 521658 683304 521660 683324
rect 521660 683304 521712 683324
rect 521712 683304 521714 683324
rect 74446 27648 74502 27704
rect 74722 27648 74778 27704
rect 540242 684528 540298 684584
rect 540426 684800 540482 684856
rect 540610 684936 540666 684992
rect 540794 685344 540850 685400
rect 577502 686024 577558 686080
rect 579710 674600 579766 674656
rect 579618 651072 579674 651128
rect 579710 639376 579766 639432
rect 579710 627680 579766 627736
rect 579618 604152 579674 604208
rect 579710 592456 579766 592512
rect 579710 580760 579766 580816
rect 579618 557232 579674 557288
rect 579710 545536 579766 545592
rect 579710 533840 579766 533896
rect 579802 510312 579858 510368
rect 579894 498616 579950 498672
rect 579894 486784 579950 486840
rect 579894 463392 579950 463448
rect 579894 451696 579950 451752
rect 579894 439864 579950 439920
rect 579986 416472 580042 416528
rect 579986 404776 580042 404832
rect 579986 392944 580042 393000
rect 579986 369552 580042 369608
rect 579986 357856 580042 357912
rect 579894 346024 579950 346080
rect 579986 252184 580042 252240
rect 580630 686704 580686 686760
rect 580170 686296 580226 686352
rect 580446 686024 580502 686080
rect 580262 685888 580318 685944
rect 580170 322632 580226 322688
rect 580170 310800 580226 310856
rect 580170 299104 580226 299160
rect 580170 263880 580226 263936
rect 580170 216960 580226 217016
rect 580078 181872 580134 181928
rect 580170 158344 580226 158400
rect 580170 111424 580226 111480
rect 580170 64504 580226 64560
rect 579894 29280 579950 29336
rect 580354 685480 580410 685536
rect 580538 170040 580594 170096
rect 580814 686432 580870 686488
rect 580722 228792 580778 228848
rect 580722 205264 580778 205320
rect 580906 275712 580962 275768
rect 580814 134816 580870 134872
rect 580630 123120 580686 123176
rect 580446 87896 580502 87952
rect 580354 76200 580410 76256
rect 580538 40976 580594 41032
rect 580262 17584 580318 17640
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 4797 687170 4863 687173
rect 480253 687170 480319 687173
rect 4797 687168 480319 687170
rect 4797 687112 4802 687168
rect 4858 687112 480258 687168
rect 480314 687112 480319 687168
rect 4797 687110 480319 687112
rect 4797 687107 4863 687110
rect 480253 687107 480319 687110
rect 84193 687034 84259 687037
rect 580073 687034 580139 687037
rect 84193 687032 580139 687034
rect 84193 686976 84198 687032
rect 84254 686976 580078 687032
rect 580134 686976 580139 687032
rect 84193 686974 580139 686976
rect 84193 686971 84259 686974
rect 580073 686971 580139 686974
rect 3693 686898 3759 686901
rect 506565 686898 506631 686901
rect 3693 686896 506631 686898
rect 3693 686840 3698 686896
rect 3754 686840 506570 686896
rect 506626 686840 506631 686896
rect 3693 686838 506631 686840
rect 3693 686835 3759 686838
rect 506565 686835 506631 686838
rect 75913 686762 75979 686765
rect 580625 686762 580691 686765
rect 75913 686760 580691 686762
rect 75913 686704 75918 686760
rect 75974 686704 580630 686760
rect 580686 686704 580691 686760
rect 75913 686702 580691 686704
rect 75913 686699 75979 686702
rect 580625 686699 580691 686702
rect 3877 686626 3943 686629
rect 510613 686626 510679 686629
rect 3877 686624 510679 686626
rect 3877 686568 3882 686624
rect 3938 686568 510618 686624
rect 510674 686568 510679 686624
rect 3877 686566 510679 686568
rect 3877 686563 3943 686566
rect 510613 686563 510679 686566
rect 71773 686490 71839 686493
rect 580809 686490 580875 686493
rect 71773 686488 580875 686490
rect 71773 686432 71778 686488
rect 71834 686432 580814 686488
rect 580870 686432 580875 686488
rect 71773 686430 580875 686432
rect 71773 686427 71839 686430
rect 580809 686427 580875 686430
rect 57973 686354 58039 686357
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 57973 686352 578618 686354
rect 57973 686296 57978 686352
rect 58034 686296 578618 686352
rect 57973 686294 578618 686296
rect 57973 686291 58039 686294
rect 3509 686218 3575 686221
rect 528093 686218 528159 686221
rect 3509 686216 528159 686218
rect 3509 686160 3514 686216
rect 3570 686160 528098 686216
rect 528154 686160 528159 686216
rect 3509 686158 528159 686160
rect 3509 686155 3575 686158
rect 528093 686155 528159 686158
rect 45553 686082 45619 686085
rect 577497 686082 577563 686085
rect 45553 686080 577563 686082
rect 45553 686024 45558 686080
rect 45614 686024 577502 686080
rect 577558 686024 577563 686080
rect 45553 686022 577563 686024
rect 578558 686082 578618 686294
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 580441 686082 580507 686085
rect 578558 686080 580507 686082
rect 578558 686024 580446 686080
rect 580502 686024 580507 686080
rect 578558 686022 580507 686024
rect 45553 686019 45619 686022
rect 577497 686019 577563 686022
rect 580441 686019 580507 686022
rect 41413 685946 41479 685949
rect 580257 685946 580323 685949
rect 41413 685944 580323 685946
rect 41413 685888 41418 685944
rect 41474 685888 580262 685944
rect 580318 685888 580323 685944
rect 41413 685886 580323 685888
rect 41413 685883 41479 685886
rect 580257 685883 580323 685886
rect 233233 685538 233299 685541
rect 580349 685538 580415 685541
rect 233233 685536 580415 685538
rect 233233 685480 233238 685536
rect 233294 685480 580354 685536
rect 580410 685480 580415 685536
rect 233233 685478 580415 685480
rect 233233 685475 233299 685478
rect 580349 685475 580415 685478
rect 120901 685402 120967 685405
rect 540789 685402 540855 685405
rect 120901 685400 540855 685402
rect 120901 685344 120906 685400
rect 120962 685344 540794 685400
rect 540850 685344 540855 685400
rect 120901 685342 540855 685344
rect 120901 685339 120967 685342
rect 540789 685339 540855 685342
rect 39389 685266 39455 685269
rect 488625 685266 488691 685269
rect 39389 685264 488691 685266
rect 39389 685208 39394 685264
rect 39450 685208 488630 685264
rect 488686 685208 488691 685264
rect 39389 685206 488691 685208
rect 39389 685203 39455 685206
rect 488625 685203 488691 685206
rect 6177 685130 6243 685133
rect 462313 685130 462379 685133
rect 6177 685128 462379 685130
rect 6177 685072 6182 685128
rect 6238 685072 462318 685128
rect 462374 685072 462379 685128
rect 6177 685070 462379 685072
rect 6177 685067 6243 685070
rect 462313 685067 462379 685070
rect 81341 684994 81407 684997
rect 356605 684994 356671 684997
rect 81341 684992 356671 684994
rect 81341 684936 81346 684992
rect 81402 684936 356610 684992
rect 356666 684936 356671 684992
rect 81341 684934 356671 684936
rect 81341 684931 81407 684934
rect 356605 684931 356671 684934
rect 357341 684994 357407 684997
rect 540605 684994 540671 684997
rect 357341 684992 540671 684994
rect 357341 684936 357346 684992
rect 357402 684936 540610 684992
rect 540666 684936 540671 684992
rect 357341 684934 540671 684936
rect 357341 684931 357407 684934
rect 540605 684931 540671 684934
rect 68277 684858 68343 684861
rect 356973 684858 357039 684861
rect 68277 684856 357039 684858
rect 68277 684800 68282 684856
rect 68338 684800 356978 684856
rect 357034 684800 357039 684856
rect 68277 684798 357039 684800
rect 68277 684795 68343 684798
rect 356973 684795 357039 684798
rect 357341 684858 357407 684861
rect 540421 684858 540487 684861
rect 357341 684856 540487 684858
rect 357341 684800 357346 684856
rect 357402 684800 540426 684856
rect 540482 684800 540487 684856
rect 357341 684798 540487 684800
rect 357341 684795 357407 684798
rect 540421 684795 540487 684798
rect 24117 684722 24183 684725
rect 357157 684722 357223 684725
rect 24117 684720 357223 684722
rect 24117 684664 24122 684720
rect 24178 684664 357162 684720
rect 357218 684664 357223 684720
rect 24117 684662 357223 684664
rect 24117 684659 24183 684662
rect 357157 684659 357223 684662
rect 357341 684722 357407 684725
rect 501781 684722 501847 684725
rect 357341 684720 501847 684722
rect 357341 684664 357346 684720
rect 357402 684664 501786 684720
rect 501842 684664 501847 684720
rect 357341 684662 501847 684664
rect 357341 684659 357407 684662
rect 501781 684659 501847 684662
rect 55121 684586 55187 684589
rect 540237 684586 540303 684589
rect 55121 684584 540303 684586
rect 55121 684528 55126 684584
rect 55182 684528 540242 684584
rect 540298 684528 540303 684584
rect 55121 684526 540303 684528
rect 55121 684523 55187 684526
rect 540237 684523 540303 684526
rect 357341 684450 357407 684453
rect 357341 684448 357450 684450
rect 357341 684392 357346 684448
rect 357402 684392 357450 684448
rect 357341 684387 357450 684392
rect 277301 684314 277367 684317
rect 298185 684314 298251 684317
rect 302141 684314 302207 684317
rect 277301 684312 292498 684314
rect 277301 684256 277306 684312
rect 277362 684256 292498 684312
rect 277301 684254 292498 684256
rect 277301 684251 277367 684254
rect 276933 684042 276999 684045
rect 280613 684042 280679 684045
rect 276933 684040 280679 684042
rect 276933 683984 276938 684040
rect 276994 683984 280618 684040
rect 280674 683984 280679 684040
rect 276933 683982 280679 683984
rect 292438 684042 292498 684254
rect 298185 684312 302207 684314
rect 298185 684256 298190 684312
rect 298246 684256 302146 684312
rect 302202 684256 302207 684312
rect 298185 684254 302207 684256
rect 357390 684314 357450 684387
rect 360101 684314 360167 684317
rect 357390 684312 360167 684314
rect 357390 684256 360106 684312
rect 360162 684256 360167 684312
rect 357390 684254 360167 684256
rect 298185 684251 298251 684254
rect 302141 684251 302207 684254
rect 360101 684251 360167 684254
rect 367001 684314 367067 684317
rect 379329 684314 379395 684317
rect 367001 684312 369778 684314
rect 367001 684256 367006 684312
rect 367062 684256 369778 684312
rect 367001 684254 369778 684256
rect 367001 684251 367067 684254
rect 298093 684178 298159 684181
rect 292622 684176 298159 684178
rect 292622 684120 298098 684176
rect 298154 684120 298159 684176
rect 292622 684118 298159 684120
rect 292622 684042 292682 684118
rect 298093 684115 298159 684118
rect 302233 684178 302299 684181
rect 312445 684178 312511 684181
rect 302233 684176 312511 684178
rect 302233 684120 302238 684176
rect 302294 684120 312450 684176
rect 312506 684120 312511 684176
rect 302233 684118 312511 684120
rect 302233 684115 302299 684118
rect 312445 684115 312511 684118
rect 318793 684178 318859 684181
rect 328361 684178 328427 684181
rect 318793 684176 328427 684178
rect 318793 684120 318798 684176
rect 318854 684120 328366 684176
rect 328422 684120 328427 684176
rect 318793 684118 328427 684120
rect 318793 684115 318859 684118
rect 328361 684115 328427 684118
rect 333237 684178 333303 684181
rect 357341 684178 357407 684181
rect 333237 684176 357407 684178
rect 333237 684120 333242 684176
rect 333298 684120 357346 684176
rect 357402 684120 357407 684176
rect 333237 684118 357407 684120
rect 333237 684115 333303 684118
rect 357341 684115 357407 684118
rect 292438 683982 292682 684042
rect 311157 684042 311223 684045
rect 312997 684042 313063 684045
rect 311157 684040 313063 684042
rect 311157 683984 311162 684040
rect 311218 683984 313002 684040
rect 313058 683984 313063 684040
rect 311157 683982 313063 683984
rect 276933 683979 276999 683982
rect 280613 683979 280679 683982
rect 311157 683979 311223 683982
rect 312997 683979 313063 683982
rect 328453 684042 328519 684045
rect 333421 684042 333487 684045
rect 328453 684040 333487 684042
rect 328453 683984 328458 684040
rect 328514 683984 333426 684040
rect 333482 683984 333487 684040
rect 328453 683982 333487 683984
rect 328453 683979 328519 683982
rect 333421 683979 333487 683982
rect 360101 684042 360167 684045
rect 367001 684042 367067 684045
rect 360101 684040 367067 684042
rect 360101 683984 360106 684040
rect 360162 683984 367006 684040
rect 367062 683984 367067 684040
rect 360101 683982 367067 683984
rect 369718 684042 369778 684254
rect 376710 684312 379395 684314
rect 376710 684256 379334 684312
rect 379390 684256 379395 684312
rect 376710 684254 379395 684256
rect 376710 684178 376770 684254
rect 379329 684251 379395 684254
rect 386321 684314 386387 684317
rect 398741 684314 398807 684317
rect 386321 684312 389098 684314
rect 386321 684256 386326 684312
rect 386382 684256 389098 684312
rect 386321 684254 389098 684256
rect 386321 684251 386387 684254
rect 369902 684118 376770 684178
rect 369902 684042 369962 684118
rect 369718 683982 369962 684042
rect 389038 684042 389098 684254
rect 396030 684312 398807 684314
rect 396030 684256 398746 684312
rect 398802 684256 398807 684312
rect 396030 684254 398807 684256
rect 396030 684178 396090 684254
rect 398741 684251 398807 684254
rect 405641 684314 405707 684317
rect 418061 684314 418127 684317
rect 405641 684312 408418 684314
rect 405641 684256 405646 684312
rect 405702 684256 408418 684312
rect 405641 684254 408418 684256
rect 405641 684251 405707 684254
rect 389222 684118 396090 684178
rect 389222 684042 389282 684118
rect 389038 683982 389282 684042
rect 408358 684042 408418 684254
rect 415350 684312 418127 684314
rect 415350 684256 418066 684312
rect 418122 684256 418127 684312
rect 415350 684254 418127 684256
rect 415350 684178 415410 684254
rect 418061 684251 418127 684254
rect 424961 684314 425027 684317
rect 437381 684314 437447 684317
rect 424961 684312 427738 684314
rect 424961 684256 424966 684312
rect 425022 684256 427738 684312
rect 424961 684254 427738 684256
rect 424961 684251 425027 684254
rect 408542 684118 415410 684178
rect 408542 684042 408602 684118
rect 408358 683982 408602 684042
rect 427678 684042 427738 684254
rect 434670 684312 437447 684314
rect 434670 684256 437386 684312
rect 437442 684256 437447 684312
rect 434670 684254 437447 684256
rect 434670 684178 434730 684254
rect 437381 684251 437447 684254
rect 444281 684314 444347 684317
rect 456701 684314 456767 684317
rect 444281 684312 447058 684314
rect 444281 684256 444286 684312
rect 444342 684256 447058 684312
rect 444281 684254 447058 684256
rect 444281 684251 444347 684254
rect 427862 684118 434730 684178
rect 427862 684042 427922 684118
rect 427678 683982 427922 684042
rect 446998 684042 447058 684254
rect 453990 684312 456767 684314
rect 453990 684256 456706 684312
rect 456762 684256 456767 684312
rect 453990 684254 456767 684256
rect 453990 684178 454050 684254
rect 456701 684251 456767 684254
rect 463601 684314 463667 684317
rect 476021 684314 476087 684317
rect 463601 684312 466378 684314
rect 463601 684256 463606 684312
rect 463662 684256 466378 684312
rect 463601 684254 466378 684256
rect 463601 684251 463667 684254
rect 447182 684118 454050 684178
rect 447182 684042 447242 684118
rect 446998 683982 447242 684042
rect 466318 684042 466378 684254
rect 473310 684312 476087 684314
rect 473310 684256 476026 684312
rect 476082 684256 476087 684312
rect 473310 684254 476087 684256
rect 473310 684178 473370 684254
rect 476021 684251 476087 684254
rect 482921 684314 482987 684317
rect 495341 684314 495407 684317
rect 482921 684312 485698 684314
rect 482921 684256 482926 684312
rect 482982 684256 485698 684312
rect 482921 684254 485698 684256
rect 482921 684251 482987 684254
rect 466502 684118 473370 684178
rect 466502 684042 466562 684118
rect 466318 683982 466562 684042
rect 485638 684042 485698 684254
rect 492630 684312 495407 684314
rect 492630 684256 495346 684312
rect 495402 684256 495407 684312
rect 492630 684254 495407 684256
rect 492630 684178 492690 684254
rect 495341 684251 495407 684254
rect 485822 684118 492690 684178
rect 514710 684118 524338 684178
rect 485822 684042 485882 684118
rect 485638 683982 485882 684042
rect 360101 683979 360167 683982
rect 367001 683979 367067 683982
rect 22737 683906 22803 683909
rect 493041 683906 493107 683909
rect 22737 683904 493107 683906
rect 22737 683848 22742 683904
rect 22798 683848 493046 683904
rect 493102 683848 493107 683904
rect 22737 683846 493107 683848
rect 22737 683843 22803 683846
rect 493041 683843 493107 683846
rect 509233 683906 509299 683909
rect 514710 683906 514770 684118
rect 509233 683904 514770 683906
rect 509233 683848 509238 683904
rect 509294 683848 514770 683904
rect 509233 683846 514770 683848
rect 509233 683843 509299 683846
rect 3417 683770 3483 683773
rect 6821 683770 6887 683773
rect 3417 683768 6887 683770
rect 3417 683712 3422 683768
rect 3478 683712 6826 683768
rect 6882 683712 6887 683768
rect 3417 683710 6887 683712
rect 3417 683707 3483 683710
rect 6821 683707 6887 683710
rect 16573 683770 16639 683773
rect 35801 683770 35867 683773
rect 16573 683768 35867 683770
rect 16573 683712 16578 683768
rect 16634 683712 35806 683768
rect 35862 683712 35867 683768
rect 16573 683710 35867 683712
rect 16573 683707 16639 683710
rect 35801 683707 35867 683710
rect 39297 683770 39363 683773
rect 331213 683770 331279 683773
rect 39297 683768 331279 683770
rect 39297 683712 39302 683768
rect 39358 683712 331218 683768
rect 331274 683712 331279 683768
rect 39297 683710 331279 683712
rect 39297 683707 39363 683710
rect 331213 683707 331279 683710
rect 331397 683770 331463 683773
rect 514937 683770 515003 683773
rect 331397 683768 515003 683770
rect 331397 683712 331402 683768
rect 331458 683712 514942 683768
rect 514998 683712 515003 683768
rect 331397 683710 515003 683712
rect 331397 683707 331463 683710
rect 514937 683707 515003 683710
rect 3969 683634 4035 683637
rect 331213 683634 331279 683637
rect 3969 683632 331279 683634
rect 3969 683576 3974 683632
rect 4030 683576 331218 683632
rect 331274 683576 331279 683632
rect 3969 683574 331279 683576
rect 3969 683571 4035 683574
rect 331213 683571 331279 683574
rect 331397 683634 331463 683637
rect 497457 683634 497523 683637
rect 331397 683632 497523 683634
rect 331397 683576 331402 683632
rect 331458 683576 497462 683632
rect 497518 683576 497523 683632
rect 331397 683574 497523 683576
rect 331397 683571 331463 683574
rect 497457 683571 497523 683574
rect 497917 683634 497983 683637
rect 509233 683634 509299 683637
rect 497917 683632 509299 683634
rect 497917 683576 497922 683632
rect 497978 683576 509238 683632
rect 509294 683576 509299 683632
rect 497917 683574 509299 683576
rect 524278 683634 524338 684118
rect 532693 683634 532759 683637
rect 524278 683632 532759 683634
rect 524278 683576 532698 683632
rect 532754 683576 532759 683632
rect 524278 683574 532759 683576
rect 497917 683571 497983 683574
rect 509233 683571 509299 683574
rect 532693 683571 532759 683574
rect 3601 683498 3667 683501
rect 331213 683498 331279 683501
rect 3601 683496 331279 683498
rect 3601 683440 3606 683496
rect 3662 683440 331218 683496
rect 331274 683440 331279 683496
rect 3601 683438 331279 683440
rect 3601 683435 3667 683438
rect 331213 683435 331279 683438
rect 331397 683498 331463 683501
rect 519353 683498 519419 683501
rect 331397 683496 519419 683498
rect 331397 683440 331402 683496
rect 331458 683440 519358 683496
rect 519414 683440 519419 683496
rect 331397 683438 519419 683440
rect 331397 683435 331463 683438
rect 519353 683435 519419 683438
rect 3785 683362 3851 683365
rect 276933 683362 276999 683365
rect 3785 683360 276999 683362
rect 3785 683304 3790 683360
rect 3846 683304 276938 683360
rect 276994 683304 276999 683360
rect 3785 683302 276999 683304
rect 3785 683299 3851 683302
rect 276933 683299 276999 683302
rect 277301 683362 277367 683365
rect 280613 683362 280679 683365
rect 311157 683362 311223 683365
rect 277301 683360 277410 683362
rect 277301 683304 277306 683360
rect 277362 683304 277410 683360
rect 277301 683299 277410 683304
rect 280613 683360 280722 683362
rect 280613 683304 280618 683360
rect 280674 683304 280722 683360
rect 280613 683299 280722 683304
rect 6821 683226 6887 683229
rect 16573 683226 16639 683229
rect 6821 683224 16639 683226
rect 6821 683168 6826 683224
rect 6882 683168 16578 683224
rect 16634 683168 16639 683224
rect 6821 683166 16639 683168
rect 6821 683163 6887 683166
rect 16573 683163 16639 683166
rect 35801 683226 35867 683229
rect 35801 683224 276122 683226
rect 35801 683168 35806 683224
rect 35862 683168 276122 683224
rect 35801 683166 276122 683168
rect 35801 683163 35867 683166
rect 276062 683090 276122 683166
rect 277350 683090 277410 683299
rect 276062 683030 277410 683090
rect 280662 683090 280722 683299
rect 289678 683360 311223 683362
rect 289678 683304 311162 683360
rect 311218 683304 311223 683360
rect 289678 683302 311223 683304
rect 289678 683090 289738 683302
rect 311157 683299 311223 683302
rect 312445 683360 312511 683365
rect 312445 683304 312450 683360
rect 312506 683304 312511 683360
rect 312445 683299 312511 683304
rect 312997 683362 313063 683365
rect 318793 683362 318859 683365
rect 333237 683362 333303 683365
rect 312997 683360 318859 683362
rect 312997 683304 313002 683360
rect 313058 683304 318798 683360
rect 318854 683304 318859 683360
rect 312997 683302 318859 683304
rect 312997 683299 313063 683302
rect 318793 683299 318859 683302
rect 333102 683360 333303 683362
rect 333102 683304 333242 683360
rect 333298 683304 333303 683360
rect 333102 683302 333303 683304
rect 312448 683226 312508 683299
rect 333102 683226 333162 683302
rect 333237 683299 333303 683302
rect 333421 683362 333487 683365
rect 521653 683362 521719 683365
rect 333421 683360 521719 683362
rect 333421 683304 333426 683360
rect 333482 683304 521658 683360
rect 521714 683304 521719 683360
rect 333421 683302 521719 683304
rect 333421 683299 333487 683302
rect 521653 683299 521719 683302
rect 312448 683166 333162 683226
rect 280662 683030 289738 683090
rect -960 682274 480 682364
rect 2773 682274 2839 682277
rect -960 682272 2839 682274
rect -960 682216 2778 682272
rect 2834 682216 2839 682272
rect -960 682214 2839 682216
rect -960 682124 480 682214
rect 2773 682211 2839 682214
rect 579705 674658 579771 674661
rect 583520 674658 584960 674748
rect 579705 674656 584960 674658
rect 579705 674600 579710 674656
rect 579766 674600 584960 674656
rect 579705 674598 584960 674600
rect 579705 674595 579771 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 2773 667994 2839 667997
rect -960 667992 2839 667994
rect -960 667936 2778 667992
rect 2834 667936 2839 667992
rect -960 667934 2839 667936
rect -960 667844 480 667934
rect 2773 667931 2839 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 2773 653578 2839 653581
rect -960 653576 2839 653578
rect -960 653520 2778 653576
rect 2834 653520 2839 653576
rect -960 653518 2839 653520
rect -960 653428 480 653518
rect 2773 653515 2839 653518
rect 579613 651130 579679 651133
rect 583520 651130 584960 651220
rect 579613 651128 584960 651130
rect 579613 651072 579618 651128
rect 579674 651072 584960 651128
rect 579613 651070 584960 651072
rect 579613 651067 579679 651070
rect 583520 650980 584960 651070
rect 579705 639434 579771 639437
rect 583520 639434 584960 639524
rect 579705 639432 584960 639434
rect 579705 639376 579710 639432
rect 579766 639376 584960 639432
rect 579705 639374 584960 639376
rect 579705 639371 579771 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 579705 627738 579771 627741
rect 583520 627738 584960 627828
rect 579705 627736 584960 627738
rect 579705 627680 579710 627736
rect 579766 627680 584960 627736
rect 579705 627678 584960 627680
rect 579705 627675 579771 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 2773 624882 2839 624885
rect -960 624880 2839 624882
rect -960 624824 2778 624880
rect 2834 624824 2839 624880
rect -960 624822 2839 624824
rect -960 624732 480 624822
rect 2773 624819 2839 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 2773 610466 2839 610469
rect -960 610464 2839 610466
rect -960 610408 2778 610464
rect 2834 610408 2839 610464
rect -960 610406 2839 610408
rect -960 610316 480 610406
rect 2773 610403 2839 610406
rect 579613 604210 579679 604213
rect 583520 604210 584960 604300
rect 579613 604208 584960 604210
rect 579613 604152 579618 604208
rect 579674 604152 584960 604208
rect 579613 604150 584960 604152
rect 579613 604147 579679 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 2773 596050 2839 596053
rect -960 596048 2839 596050
rect -960 595992 2778 596048
rect 2834 595992 2839 596048
rect -960 595990 2839 595992
rect -960 595900 480 595990
rect 2773 595987 2839 595990
rect 579705 592514 579771 592517
rect 583520 592514 584960 592604
rect 579705 592512 584960 592514
rect 579705 592456 579710 592512
rect 579766 592456 584960 592512
rect 579705 592454 584960 592456
rect 579705 592451 579771 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 579705 580818 579771 580821
rect 583520 580818 584960 580908
rect 579705 580816 584960 580818
rect 579705 580760 579710 580816
rect 579766 580760 584960 580816
rect 579705 580758 584960 580760
rect 579705 580755 579771 580758
rect 583520 580668 584960 580758
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 2773 567354 2839 567357
rect -960 567352 2839 567354
rect -960 567296 2778 567352
rect 2834 567296 2839 567352
rect -960 567294 2839 567296
rect -960 567204 480 567294
rect 2773 567291 2839 567294
rect 579613 557290 579679 557293
rect 583520 557290 584960 557380
rect 579613 557288 584960 557290
rect 579613 557232 579618 557288
rect 579674 557232 584960 557288
rect 579613 557230 584960 557232
rect 579613 557227 579679 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 2773 553074 2839 553077
rect -960 553072 2839 553074
rect -960 553016 2778 553072
rect 2834 553016 2839 553072
rect -960 553014 2839 553016
rect -960 552924 480 553014
rect 2773 553011 2839 553014
rect 579705 545594 579771 545597
rect 583520 545594 584960 545684
rect 579705 545592 584960 545594
rect 579705 545536 579710 545592
rect 579766 545536 584960 545592
rect 579705 545534 584960 545536
rect 579705 545531 579771 545534
rect 583520 545444 584960 545534
rect -960 538658 480 538748
rect 2773 538658 2839 538661
rect -960 538656 2839 538658
rect -960 538600 2778 538656
rect 2834 538600 2839 538656
rect -960 538598 2839 538600
rect -960 538508 480 538598
rect 2773 538595 2839 538598
rect 579705 533898 579771 533901
rect 583520 533898 584960 533988
rect 579705 533896 584960 533898
rect 579705 533840 579710 533896
rect 579766 533840 584960 533896
rect 579705 533838 584960 533840
rect 579705 533835 579771 533838
rect 583520 533748 584960 533838
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 579797 510370 579863 510373
rect 583520 510370 584960 510460
rect 579797 510368 584960 510370
rect 579797 510312 579802 510368
rect 579858 510312 584960 510368
rect 579797 510310 584960 510312
rect 579797 510307 579863 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 2773 509962 2839 509965
rect -960 509960 2839 509962
rect -960 509904 2778 509960
rect 2834 509904 2839 509960
rect -960 509902 2839 509904
rect -960 509812 480 509902
rect 2773 509899 2839 509902
rect 579889 498674 579955 498677
rect 583520 498674 584960 498764
rect 579889 498672 584960 498674
rect 579889 498616 579894 498672
rect 579950 498616 584960 498672
rect 579889 498614 584960 498616
rect 579889 498611 579955 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 2865 495546 2931 495549
rect -960 495544 2931 495546
rect -960 495488 2870 495544
rect 2926 495488 2931 495544
rect -960 495486 2931 495488
rect -960 495396 480 495486
rect 2865 495483 2931 495486
rect 579889 486842 579955 486845
rect 583520 486842 584960 486932
rect 579889 486840 584960 486842
rect 579889 486784 579894 486840
rect 579950 486784 584960 486840
rect 579889 486782 584960 486784
rect 579889 486779 579955 486782
rect 583520 486692 584960 486782
rect -960 481130 480 481220
rect 2865 481130 2931 481133
rect -960 481128 2931 481130
rect -960 481072 2870 481128
rect 2926 481072 2931 481128
rect -960 481070 2931 481072
rect -960 480980 480 481070
rect 2865 481067 2931 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 579889 463450 579955 463453
rect 583520 463450 584960 463540
rect 579889 463448 584960 463450
rect 579889 463392 579894 463448
rect 579950 463392 584960 463448
rect 579889 463390 584960 463392
rect 579889 463387 579955 463390
rect 583520 463300 584960 463390
rect -960 452434 480 452524
rect 2865 452434 2931 452437
rect -960 452432 2931 452434
rect -960 452376 2870 452432
rect 2926 452376 2931 452432
rect -960 452374 2931 452376
rect -960 452284 480 452374
rect 2865 452371 2931 452374
rect 579889 451754 579955 451757
rect 583520 451754 584960 451844
rect 579889 451752 584960 451754
rect 579889 451696 579894 451752
rect 579950 451696 584960 451752
rect 579889 451694 584960 451696
rect 579889 451691 579955 451694
rect 583520 451604 584960 451694
rect 579889 439922 579955 439925
rect 583520 439922 584960 440012
rect 579889 439920 584960 439922
rect 579889 439864 579894 439920
rect 579950 439864 584960 439920
rect 579889 439862 584960 439864
rect 579889 439859 579955 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 2773 438018 2839 438021
rect -960 438016 2839 438018
rect -960 437960 2778 438016
rect 2834 437960 2839 438016
rect -960 437958 2839 437960
rect -960 437868 480 437958
rect 2773 437955 2839 437958
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 2865 423738 2931 423741
rect -960 423736 2931 423738
rect -960 423680 2870 423736
rect 2926 423680 2931 423736
rect -960 423678 2931 423680
rect -960 423588 480 423678
rect 2865 423675 2931 423678
rect 579981 416530 580047 416533
rect 583520 416530 584960 416620
rect 579981 416528 584960 416530
rect 579981 416472 579986 416528
rect 580042 416472 584960 416528
rect 579981 416470 584960 416472
rect 579981 416467 580047 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 579981 404834 580047 404837
rect 583520 404834 584960 404924
rect 579981 404832 584960 404834
rect 579981 404776 579986 404832
rect 580042 404776 584960 404832
rect 579981 404774 584960 404776
rect 579981 404771 580047 404774
rect 583520 404684 584960 404774
rect -960 395042 480 395132
rect 2865 395042 2931 395045
rect -960 395040 2931 395042
rect -960 394984 2870 395040
rect 2926 394984 2931 395040
rect -960 394982 2931 394984
rect -960 394892 480 394982
rect 2865 394979 2931 394982
rect 579981 393002 580047 393005
rect 583520 393002 584960 393092
rect 579981 393000 584960 393002
rect 579981 392944 579986 393000
rect 580042 392944 584960 393000
rect 579981 392942 584960 392944
rect 579981 392939 580047 392942
rect 583520 392852 584960 392942
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 2957 380626 3023 380629
rect -960 380624 3023 380626
rect -960 380568 2962 380624
rect 3018 380568 3023 380624
rect -960 380566 3023 380568
rect -960 380476 480 380566
rect 2957 380563 3023 380566
rect 579981 369610 580047 369613
rect 583520 369610 584960 369700
rect 579981 369608 584960 369610
rect 579981 369552 579986 369608
rect 580042 369552 584960 369608
rect 579981 369550 584960 369552
rect 579981 369547 580047 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 2957 366210 3023 366213
rect -960 366208 3023 366210
rect -960 366152 2962 366208
rect 3018 366152 3023 366208
rect -960 366150 3023 366152
rect -960 366060 480 366150
rect 2957 366147 3023 366150
rect 579981 357914 580047 357917
rect 583520 357914 584960 358004
rect 579981 357912 584960 357914
rect 579981 357856 579986 357912
rect 580042 357856 584960 357912
rect 579981 357854 584960 357856
rect 579981 357851 580047 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 579889 346082 579955 346085
rect 583520 346082 584960 346172
rect 579889 346080 584960 346082
rect 579889 346024 579894 346080
rect 579950 346024 584960 346080
rect 579889 346022 584960 346024
rect 579889 346019 579955 346022
rect 583520 345932 584960 346022
rect -960 337514 480 337604
rect 2957 337514 3023 337517
rect -960 337512 3023 337514
rect -960 337456 2962 337512
rect 3018 337456 3023 337512
rect -960 337454 3023 337456
rect -960 337364 480 337454
rect 2957 337451 3023 337454
rect 583520 334236 584960 334476
rect -960 323098 480 323188
rect 2957 323098 3023 323101
rect -960 323096 3023 323098
rect -960 323040 2962 323096
rect 3018 323040 3023 323096
rect -960 323038 3023 323040
rect -960 322948 480 323038
rect 2957 323035 3023 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3049 308818 3115 308821
rect -960 308816 3115 308818
rect -960 308760 3054 308816
rect 3110 308760 3115 308816
rect -960 308758 3115 308760
rect -960 308668 480 308758
rect 3049 308755 3115 308758
rect 580165 299162 580231 299165
rect 583520 299162 584960 299252
rect 580165 299160 584960 299162
rect 580165 299104 580170 299160
rect 580226 299104 584960 299160
rect 580165 299102 584960 299104
rect 580165 299099 580231 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 3049 294402 3115 294405
rect -960 294400 3115 294402
rect -960 294344 3054 294400
rect 3110 294344 3115 294400
rect -960 294342 3115 294344
rect -960 294252 480 294342
rect 3049 294339 3115 294342
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 3141 280122 3207 280125
rect -960 280120 3207 280122
rect -960 280064 3146 280120
rect 3202 280064 3207 280120
rect -960 280062 3207 280064
rect -960 279972 480 280062
rect 3141 280059 3207 280062
rect 580901 275770 580967 275773
rect 583520 275770 584960 275860
rect 580901 275768 584960 275770
rect 580901 275712 580906 275768
rect 580962 275712 584960 275768
rect 580901 275710 584960 275712
rect 580901 275707 580967 275710
rect 583520 275620 584960 275710
rect -960 265706 480 265796
rect 3233 265706 3299 265709
rect -960 265704 3299 265706
rect -960 265648 3238 265704
rect 3294 265648 3299 265704
rect -960 265646 3299 265648
rect -960 265556 480 265646
rect 3233 265643 3299 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 579981 252242 580047 252245
rect 583520 252242 584960 252332
rect 579981 252240 584960 252242
rect 579981 252184 579986 252240
rect 580042 252184 584960 252240
rect 579981 252182 584960 252184
rect 579981 252179 580047 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3141 251290 3207 251293
rect -960 251288 3207 251290
rect -960 251232 3146 251288
rect 3202 251232 3207 251288
rect -960 251230 3207 251232
rect -960 251140 480 251230
rect 3141 251227 3207 251230
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 3325 237010 3391 237013
rect -960 237008 3391 237010
rect -960 236952 3330 237008
rect 3386 236952 3391 237008
rect -960 236950 3391 236952
rect -960 236860 480 236950
rect 3325 236947 3391 236950
rect 580717 228850 580783 228853
rect 583520 228850 584960 228940
rect 580717 228848 584960 228850
rect 580717 228792 580722 228848
rect 580778 228792 584960 228848
rect 580717 228790 584960 228792
rect 580717 228787 580783 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 3325 222594 3391 222597
rect -960 222592 3391 222594
rect -960 222536 3330 222592
rect 3386 222536 3391 222592
rect -960 222534 3391 222536
rect -960 222444 480 222534
rect 3325 222531 3391 222534
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect -960 208178 480 208268
rect 2773 208178 2839 208181
rect -960 208176 2839 208178
rect -960 208120 2778 208176
rect 2834 208120 2839 208176
rect -960 208118 2839 208120
rect -960 208028 480 208118
rect 2773 208115 2839 208118
rect 580717 205322 580783 205325
rect 583520 205322 584960 205412
rect 580717 205320 584960 205322
rect 580717 205264 580722 205320
rect 580778 205264 584960 205320
rect 580717 205262 584960 205264
rect 580717 205259 580783 205262
rect 583520 205172 584960 205262
rect -960 193898 480 193988
rect 4061 193898 4127 193901
rect -960 193896 4127 193898
rect -960 193840 4066 193896
rect 4122 193840 4127 193896
rect -960 193838 4127 193840
rect -960 193748 480 193838
rect 4061 193835 4127 193838
rect 583520 193476 584960 193716
rect 580073 181930 580139 181933
rect 583520 181930 584960 182020
rect 580073 181928 584960 181930
rect 580073 181872 580078 181928
rect 580134 181872 584960 181928
rect 580073 181870 584960 181872
rect 580073 181867 580139 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 2773 179482 2839 179485
rect -960 179480 2839 179482
rect -960 179424 2778 179480
rect 2834 179424 2839 179480
rect -960 179422 2839 179424
rect -960 179332 480 179422
rect 2773 179419 2839 179422
rect 580533 170098 580599 170101
rect 583520 170098 584960 170188
rect 580533 170096 584960 170098
rect 580533 170040 580538 170096
rect 580594 170040 584960 170096
rect 580533 170038 584960 170040
rect 580533 170035 580599 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 3141 165066 3207 165069
rect -960 165064 3207 165066
rect -960 165008 3146 165064
rect 3202 165008 3207 165064
rect -960 165006 3207 165008
rect -960 164916 480 165006
rect 3141 165003 3207 165006
rect 580165 158402 580231 158405
rect 583520 158402 584960 158492
rect 580165 158400 584960 158402
rect 580165 158344 580170 158400
rect 580226 158344 584960 158400
rect 580165 158342 584960 158344
rect 580165 158339 580231 158342
rect 583520 158252 584960 158342
rect -960 150786 480 150876
rect 3969 150786 4035 150789
rect -960 150784 4035 150786
rect -960 150728 3974 150784
rect 4030 150728 4035 150784
rect -960 150726 4035 150728
rect -960 150636 480 150726
rect 3969 150723 4035 150726
rect 583520 146556 584960 146796
rect -960 136370 480 136460
rect 3325 136370 3391 136373
rect -960 136368 3391 136370
rect -960 136312 3330 136368
rect 3386 136312 3391 136368
rect -960 136310 3391 136312
rect -960 136220 480 136310
rect 3325 136307 3391 136310
rect 580809 134874 580875 134877
rect 583520 134874 584960 134964
rect 580809 134872 584960 134874
rect 580809 134816 580814 134872
rect 580870 134816 584960 134872
rect 580809 134814 584960 134816
rect 580809 134811 580875 134814
rect 583520 134724 584960 134814
rect 580625 123178 580691 123181
rect 583520 123178 584960 123268
rect 580625 123176 584960 123178
rect 580625 123120 580630 123176
rect 580686 123120 584960 123176
rect 580625 123118 584960 123120
rect 580625 123115 580691 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3325 122090 3391 122093
rect -960 122088 3391 122090
rect -960 122032 3330 122088
rect 3386 122032 3391 122088
rect -960 122030 3391 122032
rect -960 121940 480 122030
rect 3325 122027 3391 122030
rect 580165 111482 580231 111485
rect 583520 111482 584960 111572
rect 580165 111480 584960 111482
rect 580165 111424 580170 111480
rect 580226 111424 584960 111480
rect 580165 111422 584960 111424
rect 580165 111419 580231 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3877 107674 3943 107677
rect -960 107672 3943 107674
rect -960 107616 3882 107672
rect 3938 107616 3943 107672
rect -960 107614 3943 107616
rect -960 107524 480 107614
rect 3877 107611 3943 107614
rect 583520 99636 584960 99876
rect -960 93258 480 93348
rect 3693 93258 3759 93261
rect -960 93256 3759 93258
rect -960 93200 3698 93256
rect 3754 93200 3759 93256
rect -960 93198 3759 93200
rect -960 93108 480 93198
rect 3693 93195 3759 93198
rect 580441 87954 580507 87957
rect 583520 87954 584960 88044
rect 580441 87952 584960 87954
rect 580441 87896 580446 87952
rect 580502 87896 584960 87952
rect 580441 87894 584960 87896
rect 580441 87891 580507 87894
rect 583520 87804 584960 87894
rect -960 78978 480 79068
rect 3325 78978 3391 78981
rect -960 78976 3391 78978
rect -960 78920 3330 78976
rect 3386 78920 3391 78976
rect -960 78918 3391 78920
rect -960 78828 480 78918
rect 3325 78915 3391 78918
rect 580349 76258 580415 76261
rect 583520 76258 584960 76348
rect 580349 76256 584960 76258
rect 580349 76200 580354 76256
rect 580410 76200 584960 76256
rect 580349 76198 584960 76200
rect 580349 76195 580415 76198
rect 583520 76108 584960 76198
rect -960 64562 480 64652
rect 3785 64562 3851 64565
rect -960 64560 3851 64562
rect -960 64504 3790 64560
rect 3846 64504 3851 64560
rect -960 64502 3851 64504
rect -960 64412 480 64502
rect 3785 64499 3851 64502
rect 580165 64562 580231 64565
rect 583520 64562 584960 64652
rect 580165 64560 584960 64562
rect 580165 64504 580170 64560
rect 580226 64504 584960 64560
rect 580165 64502 584960 64504
rect 580165 64499 580231 64502
rect 583520 64412 584960 64502
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3601 50146 3667 50149
rect -960 50144 3667 50146
rect -960 50088 3606 50144
rect 3662 50088 3667 50144
rect -960 50086 3667 50088
rect -960 49996 480 50086
rect 3601 50083 3667 50086
rect 580533 41034 580599 41037
rect 583520 41034 584960 41124
rect 580533 41032 584960 41034
rect 580533 40976 580538 41032
rect 580594 40976 584960 41032
rect 580533 40974 584960 40976
rect 580533 40971 580599 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 3509 35866 3575 35869
rect -960 35864 3575 35866
rect -960 35808 3514 35864
rect 3570 35808 3575 35864
rect -960 35806 3575 35808
rect -960 35716 480 35806
rect 3509 35803 3575 35806
rect 579889 29338 579955 29341
rect 583520 29338 584960 29428
rect 579889 29336 584960 29338
rect 579889 29280 579894 29336
rect 579950 29280 584960 29336
rect 579889 29278 584960 29280
rect 579889 29275 579955 29278
rect 583520 29188 584960 29278
rect 74441 27706 74507 27709
rect 74717 27706 74783 27709
rect 74441 27704 74783 27706
rect 74441 27648 74446 27704
rect 74502 27648 74722 27704
rect 74778 27648 74783 27704
rect 74441 27646 74783 27648
rect 74441 27643 74507 27646
rect 74717 27643 74783 27646
rect -960 21450 480 21540
rect 3509 21450 3575 21453
rect -960 21448 3575 21450
rect -960 21392 3514 21448
rect 3570 21392 3575 21448
rect -960 21390 3575 21392
rect -960 21300 480 21390
rect 3509 21387 3575 21390
rect 580257 17642 580323 17645
rect 583520 17642 584960 17732
rect 580257 17640 584960 17642
rect 580257 17584 580262 17640
rect 580318 17584 584960 17640
rect 580257 17582 584960 17584
rect 580257 17579 580323 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 684000 41004 689498
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 684000 44604 693098
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 684000 48204 696698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 684000 55404 705222
rect 58404 684000 59004 707102
rect 62004 684000 62604 708982
rect 65604 684000 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 684000 73404 685898
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 684000 77004 689498
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 684000 80604 693098
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 684000 84204 696698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 684000 91404 705222
rect 94404 684000 95004 707102
rect 98004 684000 98604 708982
rect 101604 684000 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 684000 109404 685898
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 684000 113004 689498
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 684000 116604 693098
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 684000 120204 696698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 684000 127404 705222
rect 130404 684000 131004 707102
rect 134004 684000 134604 708982
rect 137604 684000 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 684000 145404 685898
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 684000 149004 689498
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 684000 152604 693098
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 684000 156204 696698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 684000 163404 705222
rect 166404 684000 167004 707102
rect 170004 684000 170604 708982
rect 173604 684000 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 684000 181404 685898
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 684000 185004 689498
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 684000 188604 693098
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 684000 192204 696698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 684000 199404 705222
rect 202404 684000 203004 707102
rect 206004 684000 206604 708982
rect 209604 684000 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 684000 217404 685898
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 684000 221004 689498
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 684000 224604 693098
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 684000 228204 696698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 684000 235404 705222
rect 238404 684000 239004 707102
rect 242004 684000 242604 708982
rect 245604 684000 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 684000 253404 685898
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 684000 257004 689498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 684000 260604 693098
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 684000 264204 696698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 684000 271404 705222
rect 274404 684000 275004 707102
rect 278004 684000 278604 708982
rect 281604 684000 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 684000 289404 685898
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 684000 293004 689498
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 684000 296604 693098
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 684000 300204 696698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 684000 307404 705222
rect 310404 684000 311004 707102
rect 314004 684000 314604 708982
rect 317604 684000 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 684000 325404 685898
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 684000 329004 689498
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 684000 332604 693098
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 684000 336204 696698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 684000 343404 705222
rect 346404 684000 347004 707102
rect 350004 684000 350604 708982
rect 353604 684000 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 684000 361404 685898
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 684000 365004 689498
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 684000 368604 693098
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 684000 372204 696698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 684000 379404 705222
rect 382404 684000 383004 707102
rect 386004 684000 386604 708982
rect 389604 684000 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 684000 397404 685898
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 684000 401004 689498
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 684000 404604 693098
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 684000 408204 696698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 684000 415404 705222
rect 418404 684000 419004 707102
rect 422004 684000 422604 708982
rect 425604 684000 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 684000 433404 685898
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 684000 437004 689498
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 684000 440604 693098
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 684000 444204 696698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 684000 451404 705222
rect 454404 684000 455004 707102
rect 458004 684000 458604 708982
rect 461604 684000 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 684000 469404 685898
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 684000 473004 689498
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 684000 476604 693098
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 684000 480204 696698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 684000 487404 705222
rect 490404 684000 491004 707102
rect 494004 684000 494604 708982
rect 497604 684000 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 684000 505404 685898
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 684000 509004 689498
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 684000 512604 693098
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 684000 516204 696698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 684000 523404 705222
rect 526404 684000 527004 707102
rect 530004 684000 530604 708982
rect 533604 684000 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 59096 668454 59416 668476
rect 59096 668218 59138 668454
rect 59374 668218 59416 668454
rect 59096 668134 59416 668218
rect 59096 667898 59138 668134
rect 59374 667898 59416 668134
rect 59096 667876 59416 667898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 43736 650454 44056 650476
rect 43736 650218 43778 650454
rect 44014 650218 44056 650454
rect 43736 650134 44056 650218
rect 43736 649898 43778 650134
rect 44014 649898 44056 650134
rect 43736 649876 44056 649898
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 59096 632454 59416 632476
rect 59096 632218 59138 632454
rect 59374 632218 59416 632454
rect 59096 632134 59416 632218
rect 59096 631898 59138 632134
rect 59374 631898 59416 632134
rect 59096 631876 59416 631898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 43736 614454 44056 614476
rect 43736 614218 43778 614454
rect 44014 614218 44056 614454
rect 43736 614134 44056 614218
rect 43736 613898 43778 614134
rect 44014 613898 44056 614134
rect 43736 613876 44056 613898
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 59096 596454 59416 596476
rect 59096 596218 59138 596454
rect 59374 596218 59416 596454
rect 59096 596134 59416 596218
rect 59096 595898 59138 596134
rect 59374 595898 59416 596134
rect 59096 595876 59416 595898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 43736 578454 44056 578476
rect 43736 578218 43778 578454
rect 44014 578218 44056 578454
rect 43736 578134 44056 578218
rect 43736 577898 43778 578134
rect 44014 577898 44056 578134
rect 43736 577876 44056 577898
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 59096 560454 59416 560476
rect 59096 560218 59138 560454
rect 59374 560218 59416 560454
rect 59096 560134 59416 560218
rect 59096 559898 59138 560134
rect 59374 559898 59416 560134
rect 59096 559876 59416 559898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 43736 542454 44056 542476
rect 43736 542218 43778 542454
rect 44014 542218 44056 542454
rect 43736 542134 44056 542218
rect 43736 541898 43778 542134
rect 44014 541898 44056 542134
rect 43736 541876 44056 541898
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 59096 524454 59416 524476
rect 59096 524218 59138 524454
rect 59374 524218 59416 524454
rect 59096 524134 59416 524218
rect 59096 523898 59138 524134
rect 59374 523898 59416 524134
rect 59096 523876 59416 523898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 43736 506454 44056 506476
rect 43736 506218 43778 506454
rect 44014 506218 44056 506454
rect 43736 506134 44056 506218
rect 43736 505898 43778 506134
rect 44014 505898 44056 506134
rect 43736 505876 44056 505898
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 59096 488454 59416 488476
rect 59096 488218 59138 488454
rect 59374 488218 59416 488454
rect 59096 488134 59416 488218
rect 59096 487898 59138 488134
rect 59374 487898 59416 488134
rect 59096 487876 59416 487898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 43736 470454 44056 470476
rect 43736 470218 43778 470454
rect 44014 470218 44056 470454
rect 43736 470134 44056 470218
rect 43736 469898 43778 470134
rect 44014 469898 44056 470134
rect 43736 469876 44056 469898
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 59096 452454 59416 452476
rect 59096 452218 59138 452454
rect 59374 452218 59416 452454
rect 59096 452134 59416 452218
rect 59096 451898 59138 452134
rect 59374 451898 59416 452134
rect 59096 451876 59416 451898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 43736 434454 44056 434476
rect 43736 434218 43778 434454
rect 44014 434218 44056 434454
rect 43736 434134 44056 434218
rect 43736 433898 43778 434134
rect 44014 433898 44056 434134
rect 43736 433876 44056 433898
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 59096 416454 59416 416476
rect 59096 416218 59138 416454
rect 59374 416218 59416 416454
rect 59096 416134 59416 416218
rect 59096 415898 59138 416134
rect 59374 415898 59416 416134
rect 59096 415876 59416 415898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 43736 398454 44056 398476
rect 43736 398218 43778 398454
rect 44014 398218 44056 398454
rect 43736 398134 44056 398218
rect 43736 397898 43778 398134
rect 44014 397898 44056 398134
rect 43736 397876 44056 397898
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 59096 380454 59416 380476
rect 59096 380218 59138 380454
rect 59374 380218 59416 380454
rect 59096 380134 59416 380218
rect 59096 379898 59138 380134
rect 59374 379898 59416 380134
rect 59096 379876 59416 379898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 43736 362454 44056 362476
rect 43736 362218 43778 362454
rect 44014 362218 44056 362454
rect 43736 362134 44056 362218
rect 43736 361898 43778 362134
rect 44014 361898 44056 362134
rect 43736 361876 44056 361898
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 59096 344454 59416 344476
rect 59096 344218 59138 344454
rect 59374 344218 59416 344454
rect 59096 344134 59416 344218
rect 59096 343898 59138 344134
rect 59374 343898 59416 344134
rect 59096 343876 59416 343898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 43736 326454 44056 326476
rect 43736 326218 43778 326454
rect 44014 326218 44056 326454
rect 43736 326134 44056 326218
rect 43736 325898 43778 326134
rect 44014 325898 44056 326134
rect 43736 325876 44056 325898
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 59096 308454 59416 308476
rect 59096 308218 59138 308454
rect 59374 308218 59416 308454
rect 59096 308134 59416 308218
rect 59096 307898 59138 308134
rect 59374 307898 59416 308134
rect 59096 307876 59416 307898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 43736 290454 44056 290476
rect 43736 290218 43778 290454
rect 44014 290218 44056 290454
rect 43736 290134 44056 290218
rect 43736 289898 43778 290134
rect 44014 289898 44056 290134
rect 43736 289876 44056 289898
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 59096 272454 59416 272476
rect 59096 272218 59138 272454
rect 59374 272218 59416 272454
rect 59096 272134 59416 272218
rect 59096 271898 59138 272134
rect 59374 271898 59416 272134
rect 59096 271876 59416 271898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 43736 254454 44056 254476
rect 43736 254218 43778 254454
rect 44014 254218 44056 254454
rect 43736 254134 44056 254218
rect 43736 253898 43778 254134
rect 44014 253898 44056 254134
rect 43736 253876 44056 253898
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 59096 236454 59416 236476
rect 59096 236218 59138 236454
rect 59374 236218 59416 236454
rect 59096 236134 59416 236218
rect 59096 235898 59138 236134
rect 59374 235898 59416 236134
rect 59096 235876 59416 235898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 43736 218454 44056 218476
rect 43736 218218 43778 218454
rect 44014 218218 44056 218454
rect 43736 218134 44056 218218
rect 43736 217898 43778 218134
rect 44014 217898 44056 218134
rect 43736 217876 44056 217898
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 59096 200454 59416 200476
rect 59096 200218 59138 200454
rect 59374 200218 59416 200454
rect 59096 200134 59416 200218
rect 59096 199898 59138 200134
rect 59374 199898 59416 200134
rect 59096 199876 59416 199898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 43736 182454 44056 182476
rect 43736 182218 43778 182454
rect 44014 182218 44056 182454
rect 43736 182134 44056 182218
rect 43736 181898 43778 182134
rect 44014 181898 44056 182134
rect 43736 181876 44056 181898
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 59096 164454 59416 164476
rect 59096 164218 59138 164454
rect 59374 164218 59416 164454
rect 59096 164134 59416 164218
rect 59096 163898 59138 164134
rect 59374 163898 59416 164134
rect 59096 163876 59416 163898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 43736 146454 44056 146476
rect 43736 146218 43778 146454
rect 44014 146218 44056 146454
rect 43736 146134 44056 146218
rect 43736 145898 43778 146134
rect 44014 145898 44056 146134
rect 43736 145876 44056 145898
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 59096 128454 59416 128476
rect 59096 128218 59138 128454
rect 59374 128218 59416 128454
rect 59096 128134 59416 128218
rect 59096 127898 59138 128134
rect 59374 127898 59416 128134
rect 59096 127876 59416 127898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 43736 110454 44056 110476
rect 43736 110218 43778 110454
rect 44014 110218 44056 110454
rect 43736 110134 44056 110218
rect 43736 109898 43778 110134
rect 44014 109898 44056 110134
rect 43736 109876 44056 109898
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 59096 92454 59416 92476
rect 59096 92218 59138 92454
rect 59374 92218 59416 92454
rect 59096 92134 59416 92218
rect 59096 91898 59138 92134
rect 59374 91898 59416 92134
rect 59096 91876 59416 91898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 43736 74454 44056 74476
rect 43736 74218 43778 74454
rect 44014 74218 44056 74454
rect 43736 74134 44056 74218
rect 43736 73898 43778 74134
rect 44014 73898 44056 74134
rect 43736 73876 44056 73898
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 42054 41004 64000
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 45654 44604 64000
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 49254 48204 64000
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 56454 55404 64000
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 60054 59004 64000
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 63654 62604 64000
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 31254 66204 64000
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 38454 73404 64000
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 42054 77004 64000
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 45654 80604 64000
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 49254 84204 64000
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 56454 91404 64000
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 60054 95004 64000
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 63654 98604 64000
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 31254 102204 64000
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 38454 109404 64000
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 42054 113004 64000
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 45654 116604 64000
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 49254 120204 64000
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 56454 127404 64000
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 60054 131004 64000
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 63654 134604 64000
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 31254 138204 64000
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 38454 145404 64000
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 42054 149004 64000
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 45654 152604 64000
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 49254 156204 64000
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 56454 163404 64000
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 60054 167004 64000
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 63654 170604 64000
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 31254 174204 64000
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 38454 181404 64000
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 42054 185004 64000
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 45654 188604 64000
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 49254 192204 64000
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 56454 199404 64000
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 60054 203004 64000
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 63654 206604 64000
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 31254 210204 64000
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 38454 217404 64000
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 42054 221004 64000
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 45654 224604 64000
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 49254 228204 64000
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 56454 235404 64000
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 60054 239004 64000
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 63654 242604 64000
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 31254 246204 64000
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 38454 253404 64000
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 42054 257004 64000
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 45654 260604 64000
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 49254 264204 64000
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 56454 271404 64000
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 60054 275004 64000
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 63654 278604 64000
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 31254 282204 64000
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 38454 289404 64000
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 42054 293004 64000
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 45654 296604 64000
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 49254 300204 64000
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 56454 307404 64000
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 60054 311004 64000
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 63654 314604 64000
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 31254 318204 64000
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 38454 325404 64000
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 42054 329004 64000
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 45654 332604 64000
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 49254 336204 64000
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 56454 343404 64000
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 60054 347004 64000
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 63654 350604 64000
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 31254 354204 64000
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 38454 361404 64000
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 42054 365004 64000
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 45654 368604 64000
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 49254 372204 64000
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 56454 379404 64000
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 60054 383004 64000
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 63654 386604 64000
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 31254 390204 64000
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 38454 397404 64000
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 42054 401004 64000
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 45654 404604 64000
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 49254 408204 64000
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 56454 415404 64000
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 60054 419004 64000
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 63654 422604 64000
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 31254 426204 64000
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 38454 433404 64000
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 42054 437004 64000
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 45654 440604 64000
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 49254 444204 64000
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 56454 451404 64000
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 60054 455004 64000
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 63654 458604 64000
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 31254 462204 64000
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 38454 469404 64000
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 42054 473004 64000
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 45654 476604 64000
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 49254 480204 64000
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 56454 487404 64000
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 60054 491004 64000
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 63654 494604 64000
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 31254 498204 64000
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 38454 505404 64000
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 42054 509004 64000
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 45654 512604 64000
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 49254 516204 64000
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 56454 523404 64000
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 60054 527004 64000
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 63654 530604 64000
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 31254 534204 64000
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 59138 668218 59374 668454
rect 59138 667898 59374 668134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 43778 650218 44014 650454
rect 43778 649898 44014 650134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 59138 632218 59374 632454
rect 59138 631898 59374 632134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 43778 614218 44014 614454
rect 43778 613898 44014 614134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 59138 596218 59374 596454
rect 59138 595898 59374 596134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 43778 578218 44014 578454
rect 43778 577898 44014 578134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 59138 560218 59374 560454
rect 59138 559898 59374 560134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 43778 542218 44014 542454
rect 43778 541898 44014 542134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 59138 524218 59374 524454
rect 59138 523898 59374 524134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 43778 506218 44014 506454
rect 43778 505898 44014 506134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 59138 488218 59374 488454
rect 59138 487898 59374 488134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 43778 470218 44014 470454
rect 43778 469898 44014 470134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 59138 452218 59374 452454
rect 59138 451898 59374 452134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 43778 434218 44014 434454
rect 43778 433898 44014 434134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 59138 416218 59374 416454
rect 59138 415898 59374 416134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 43778 398218 44014 398454
rect 43778 397898 44014 398134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 59138 380218 59374 380454
rect 59138 379898 59374 380134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 43778 362218 44014 362454
rect 43778 361898 44014 362134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 59138 344218 59374 344454
rect 59138 343898 59374 344134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 43778 326218 44014 326454
rect 43778 325898 44014 326134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 59138 308218 59374 308454
rect 59138 307898 59374 308134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 43778 290218 44014 290454
rect 43778 289898 44014 290134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 59138 272218 59374 272454
rect 59138 271898 59374 272134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 43778 254218 44014 254454
rect 43778 253898 44014 254134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 59138 236218 59374 236454
rect 59138 235898 59374 236134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 43778 218218 44014 218454
rect 43778 217898 44014 218134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 59138 200218 59374 200454
rect 59138 199898 59374 200134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 43778 182218 44014 182454
rect 43778 181898 44014 182134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 59138 164218 59374 164454
rect 59138 163898 59374 164134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 43778 146218 44014 146454
rect 43778 145898 44014 146134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 59138 128218 59374 128454
rect 59138 127898 59374 128134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 43778 110218 44014 110454
rect 43778 109898 44014 110134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 59138 92218 59374 92454
rect 59138 91898 59374 92134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 43778 74218 44014 74454
rect 43778 73898 44014 74134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 59096 668476 59416 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 59138 668454
rect 59374 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 59138 668134
rect 59374 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 59096 667874 59416 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 43736 650476 44056 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 43778 650454
rect 44014 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 43778 650134
rect 44014 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 43736 649874 44056 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 59096 632476 59416 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 59138 632454
rect 59374 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 59138 632134
rect 59374 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 59096 631874 59416 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 43736 614476 44056 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 43778 614454
rect 44014 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 43778 614134
rect 44014 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 43736 613874 44056 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 59096 596476 59416 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 59138 596454
rect 59374 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 59138 596134
rect 59374 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 59096 595874 59416 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 43736 578476 44056 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 43778 578454
rect 44014 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 43778 578134
rect 44014 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 43736 577874 44056 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 59096 560476 59416 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 59138 560454
rect 59374 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 59138 560134
rect 59374 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 59096 559874 59416 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 43736 542476 44056 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 43778 542454
rect 44014 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 43778 542134
rect 44014 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 43736 541874 44056 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 59096 524476 59416 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 59138 524454
rect 59374 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 59138 524134
rect 59374 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 59096 523874 59416 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 43736 506476 44056 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 43778 506454
rect 44014 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 43778 506134
rect 44014 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 43736 505874 44056 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 59096 488476 59416 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 59138 488454
rect 59374 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 59138 488134
rect 59374 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 59096 487874 59416 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 43736 470476 44056 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 43778 470454
rect 44014 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 43778 470134
rect 44014 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 43736 469874 44056 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 59096 452476 59416 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 59138 452454
rect 59374 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 59138 452134
rect 59374 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 59096 451874 59416 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 43736 434476 44056 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 43778 434454
rect 44014 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 43778 434134
rect 44014 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 43736 433874 44056 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 59096 416476 59416 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 59138 416454
rect 59374 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 59138 416134
rect 59374 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 59096 415874 59416 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 43736 398476 44056 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 43778 398454
rect 44014 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 43778 398134
rect 44014 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 43736 397874 44056 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 59096 380476 59416 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 59138 380454
rect 59374 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 59138 380134
rect 59374 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 59096 379874 59416 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 43736 362476 44056 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 43778 362454
rect 44014 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 43778 362134
rect 44014 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 43736 361874 44056 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 59096 344476 59416 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 59138 344454
rect 59374 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 59138 344134
rect 59374 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 59096 343874 59416 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 43736 326476 44056 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 43778 326454
rect 44014 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 43778 326134
rect 44014 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 43736 325874 44056 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 59096 308476 59416 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 59138 308454
rect 59374 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 59138 308134
rect 59374 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 59096 307874 59416 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 43736 290476 44056 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 43778 290454
rect 44014 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 43778 290134
rect 44014 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 43736 289874 44056 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 59096 272476 59416 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 59138 272454
rect 59374 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 59138 272134
rect 59374 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 59096 271874 59416 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 43736 254476 44056 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 43778 254454
rect 44014 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 43778 254134
rect 44014 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 43736 253874 44056 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 59096 236476 59416 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 59138 236454
rect 59374 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 59138 236134
rect 59374 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 59096 235874 59416 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 43736 218476 44056 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 43778 218454
rect 44014 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 43778 218134
rect 44014 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 43736 217874 44056 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 59096 200476 59416 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 59138 200454
rect 59374 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 59138 200134
rect 59374 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 59096 199874 59416 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 43736 182476 44056 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 43778 182454
rect 44014 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 43778 182134
rect 44014 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 43736 181874 44056 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 59096 164476 59416 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 59138 164454
rect 59374 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 59138 164134
rect 59374 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 59096 163874 59416 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 43736 146476 44056 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 43778 146454
rect 44014 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 43778 146134
rect 44014 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 43736 145874 44056 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 59096 128476 59416 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 59138 128454
rect 59374 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 59138 128134
rect 59374 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 59096 127874 59416 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 43736 110476 44056 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 43778 110454
rect 44014 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 43778 110134
rect 44014 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 43736 109874 44056 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 59096 92476 59416 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 59138 92454
rect 59374 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 59138 92134
rect 59374 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 59096 91874 59416 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 43736 74476 44056 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 43778 74454
rect 44014 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 43778 74134
rect 44014 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 43736 73874 44056 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use user_proj_example  mprj
timestamp 1608291739
transform 1 0 39999 0 1 64000
box 1 0 498978 620000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
