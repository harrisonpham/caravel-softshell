VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2694.290 89.660 2694.610 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2694.290 89.520 2899.310 89.660 ;
        RECT 2694.290 89.460 2694.610 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2694.320 89.460 2694.580 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 307.840 3298.410 308.120 3300.000 ;
        RECT 309.670 3298.410 309.950 3298.525 ;
        RECT 307.840 3298.270 309.950 3298.410 ;
        RECT 307.840 3296.000 308.120 3298.270 ;
        RECT 309.670 3298.155 309.950 3298.270 ;
        RECT 2694.310 3298.155 2694.590 3298.525 ;
        RECT 2694.380 89.750 2694.520 3298.155 ;
        RECT 2694.320 89.430 2694.580 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 309.670 3298.200 309.950 3298.480 ;
        RECT 2694.310 3298.200 2694.590 3298.480 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 309.645 3298.490 309.975 3298.505 ;
        RECT 2694.285 3298.490 2694.615 3298.505 ;
        RECT 309.645 3298.190 2694.615 3298.490 ;
        RECT 309.645 3298.175 309.975 3298.190 ;
        RECT 2694.285 3298.175 2694.615 3298.190 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 938.930 3304.020 939.250 3304.080 ;
        RECT 2693.370 3304.020 2693.690 3304.080 ;
        RECT 938.930 3303.880 2693.690 3304.020 ;
        RECT 938.930 3303.820 939.250 3303.880 ;
        RECT 2693.370 3303.820 2693.690 3303.880 ;
        RECT 2693.370 2435.660 2693.690 2435.720 ;
        RECT 2900.830 2435.660 2901.150 2435.720 ;
        RECT 2693.370 2435.520 2901.150 2435.660 ;
        RECT 2693.370 2435.460 2693.690 2435.520 ;
        RECT 2900.830 2435.460 2901.150 2435.520 ;
      LAYER via ;
        RECT 938.960 3303.820 939.220 3304.080 ;
        RECT 2693.400 3303.820 2693.660 3304.080 ;
        RECT 2693.400 2435.460 2693.660 2435.720 ;
        RECT 2900.860 2435.460 2901.120 2435.720 ;
      LAYER met2 ;
        RECT 938.960 3303.790 939.220 3304.110 ;
        RECT 2693.400 3303.790 2693.660 3304.110 ;
        RECT 939.020 3300.000 939.160 3303.790 ;
        RECT 938.960 3296.000 939.240 3300.000 ;
        RECT 2693.460 2435.750 2693.600 3303.790 ;
        RECT 2693.400 2435.430 2693.660 2435.750 ;
        RECT 2900.860 2435.430 2901.120 2435.750 ;
        RECT 2900.920 2434.245 2901.060 2435.430 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1002.410 3304.360 1002.730 3304.420 ;
        RECT 2692.910 3304.360 2693.230 3304.420 ;
        RECT 1002.410 3304.220 2693.230 3304.360 ;
        RECT 1002.410 3304.160 1002.730 3304.220 ;
        RECT 2692.910 3304.160 2693.230 3304.220 ;
        RECT 2692.910 2670.260 2693.230 2670.320 ;
        RECT 2900.830 2670.260 2901.150 2670.320 ;
        RECT 2692.910 2670.120 2901.150 2670.260 ;
        RECT 2692.910 2670.060 2693.230 2670.120 ;
        RECT 2900.830 2670.060 2901.150 2670.120 ;
      LAYER via ;
        RECT 1002.440 3304.160 1002.700 3304.420 ;
        RECT 2692.940 3304.160 2693.200 3304.420 ;
        RECT 2692.940 2670.060 2693.200 2670.320 ;
        RECT 2900.860 2670.060 2901.120 2670.320 ;
      LAYER met2 ;
        RECT 1002.440 3304.130 1002.700 3304.450 ;
        RECT 2692.940 3304.130 2693.200 3304.450 ;
        RECT 1002.500 3300.000 1002.640 3304.130 ;
        RECT 1002.440 3296.000 1002.720 3300.000 ;
        RECT 2693.000 2670.350 2693.140 3304.130 ;
        RECT 2692.940 2670.030 2693.200 2670.350 ;
        RECT 2900.860 2670.030 2901.120 2670.350 ;
        RECT 2900.920 2669.525 2901.060 2670.030 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
      LAYER met3 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1065.430 3304.700 1065.750 3304.760 ;
        RECT 2692.450 3304.700 2692.770 3304.760 ;
        RECT 1065.430 3304.560 2692.770 3304.700 ;
        RECT 1065.430 3304.500 1065.750 3304.560 ;
        RECT 2692.450 3304.500 2692.770 3304.560 ;
        RECT 2692.450 2904.860 2692.770 2904.920 ;
        RECT 2900.370 2904.860 2900.690 2904.920 ;
        RECT 2692.450 2904.720 2900.690 2904.860 ;
        RECT 2692.450 2904.660 2692.770 2904.720 ;
        RECT 2900.370 2904.660 2900.690 2904.720 ;
      LAYER via ;
        RECT 1065.460 3304.500 1065.720 3304.760 ;
        RECT 2692.480 3304.500 2692.740 3304.760 ;
        RECT 2692.480 2904.660 2692.740 2904.920 ;
        RECT 2900.400 2904.660 2900.660 2904.920 ;
      LAYER met2 ;
        RECT 1065.460 3304.470 1065.720 3304.790 ;
        RECT 2692.480 3304.470 2692.740 3304.790 ;
        RECT 1065.520 3300.000 1065.660 3304.470 ;
        RECT 1065.460 3296.000 1065.740 3300.000 ;
        RECT 2692.540 2904.950 2692.680 3304.470 ;
        RECT 2692.480 2904.630 2692.740 2904.950 ;
        RECT 2900.400 2904.630 2900.660 2904.950 ;
        RECT 2900.460 2904.125 2900.600 2904.630 ;
        RECT 2900.390 2903.755 2900.670 2904.125 ;
      LAYER via2 ;
        RECT 2900.390 2903.800 2900.670 2904.080 ;
      LAYER met3 ;
        RECT 2900.365 2904.090 2900.695 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.365 2903.790 2924.800 2904.090 ;
        RECT 2900.365 2903.775 2900.695 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1128.450 3305.040 1128.770 3305.100 ;
        RECT 2691.990 3305.040 2692.310 3305.100 ;
        RECT 1128.450 3304.900 2692.310 3305.040 ;
        RECT 1128.450 3304.840 1128.770 3304.900 ;
        RECT 2691.990 3304.840 2692.310 3304.900 ;
        RECT 2697.970 3139.460 2698.290 3139.520 ;
        RECT 2900.370 3139.460 2900.690 3139.520 ;
        RECT 2697.970 3139.320 2900.690 3139.460 ;
        RECT 2697.970 3139.260 2698.290 3139.320 ;
        RECT 2900.370 3139.260 2900.690 3139.320 ;
      LAYER via ;
        RECT 1128.480 3304.840 1128.740 3305.100 ;
        RECT 2692.020 3304.840 2692.280 3305.100 ;
        RECT 2698.000 3139.260 2698.260 3139.520 ;
        RECT 2900.400 3139.260 2900.660 3139.520 ;
      LAYER met2 ;
        RECT 1128.480 3304.810 1128.740 3305.130 ;
        RECT 2692.020 3304.810 2692.280 3305.130 ;
        RECT 1128.540 3300.000 1128.680 3304.810 ;
        RECT 1128.480 3296.000 1128.760 3300.000 ;
        RECT 2692.080 3139.405 2692.220 3304.810 ;
        RECT 2698.000 3139.405 2698.260 3139.550 ;
        RECT 2692.010 3139.035 2692.290 3139.405 ;
        RECT 2697.990 3139.035 2698.270 3139.405 ;
        RECT 2900.400 3139.230 2900.660 3139.550 ;
        RECT 2900.460 3138.725 2900.600 3139.230 ;
        RECT 2900.390 3138.355 2900.670 3138.725 ;
      LAYER via2 ;
        RECT 2692.010 3139.080 2692.290 3139.360 ;
        RECT 2697.990 3139.080 2698.270 3139.360 ;
        RECT 2900.390 3138.400 2900.670 3138.680 ;
      LAYER met3 ;
        RECT 2691.985 3139.370 2692.315 3139.385 ;
        RECT 2697.965 3139.370 2698.295 3139.385 ;
        RECT 2691.985 3139.070 2698.295 3139.370 ;
        RECT 2691.985 3139.055 2692.315 3139.070 ;
        RECT 2697.965 3139.055 2698.295 3139.070 ;
        RECT 2900.365 3138.690 2900.695 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.365 3138.390 2924.800 3138.690 ;
        RECT 2900.365 3138.375 2900.695 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1193.310 3367.600 1193.630 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 1193.310 3367.460 2901.150 3367.600 ;
        RECT 1193.310 3367.400 1193.630 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
      LAYER via ;
        RECT 1193.340 3367.400 1193.600 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 1193.340 3367.370 1193.600 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 1191.960 3299.770 1192.240 3300.000 ;
        RECT 1193.400 3299.770 1193.540 3367.370 ;
        RECT 1191.960 3299.630 1193.540 3299.770 ;
        RECT 1191.960 3296.000 1192.240 3299.630 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1254.950 3315.240 1255.270 3315.300 ;
        RECT 2795.030 3315.240 2795.350 3315.300 ;
        RECT 1254.950 3315.100 2795.350 3315.240 ;
        RECT 1254.950 3315.040 1255.270 3315.100 ;
        RECT 2795.030 3315.040 2795.350 3315.100 ;
      LAYER via ;
        RECT 1254.980 3315.040 1255.240 3315.300 ;
        RECT 2795.060 3315.040 2795.320 3315.300 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3443.930 2798.480 3517.600 ;
        RECT 2796.500 3443.790 2798.480 3443.930 ;
        RECT 2796.500 3443.250 2796.640 3443.790 ;
        RECT 2796.040 3443.110 2796.640 3443.250 ;
        RECT 2796.040 3346.690 2796.180 3443.110 ;
        RECT 2795.120 3346.550 2796.180 3346.690 ;
        RECT 2795.120 3315.330 2795.260 3346.550 ;
        RECT 1254.980 3315.010 1255.240 3315.330 ;
        RECT 2795.060 3315.010 2795.320 3315.330 ;
        RECT 1255.040 3300.000 1255.180 3315.010 ;
        RECT 1254.980 3296.000 1255.260 3300.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2470.345 3332.765 2470.515 3380.875 ;
      LAYER mcon ;
        RECT 2470.345 3380.705 2470.515 3380.875 ;
      LAYER met1 ;
        RECT 2470.270 3380.860 2470.590 3380.920 ;
        RECT 2470.075 3380.720 2470.590 3380.860 ;
        RECT 2470.270 3380.660 2470.590 3380.720 ;
        RECT 2470.285 3332.920 2470.575 3332.965 ;
        RECT 2470.730 3332.920 2471.050 3332.980 ;
        RECT 2470.285 3332.780 2471.050 3332.920 ;
        RECT 2470.285 3332.735 2470.575 3332.780 ;
        RECT 2470.730 3332.720 2471.050 3332.780 ;
        RECT 1317.970 3315.580 1318.290 3315.640 ;
        RECT 2470.730 3315.580 2471.050 3315.640 ;
        RECT 1317.970 3315.440 2471.050 3315.580 ;
        RECT 1317.970 3315.380 1318.290 3315.440 ;
        RECT 2470.730 3315.380 2471.050 3315.440 ;
      LAYER via ;
        RECT 2470.300 3380.660 2470.560 3380.920 ;
        RECT 2470.760 3332.720 2471.020 3332.980 ;
        RECT 1318.000 3315.380 1318.260 3315.640 ;
        RECT 2470.760 3315.380 2471.020 3315.640 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3430.445 2474.640 3517.230 ;
        RECT 2474.430 3430.075 2474.710 3430.445 ;
        RECT 2471.210 3429.395 2471.490 3429.765 ;
        RECT 2471.280 3394.970 2471.420 3429.395 ;
        RECT 2470.360 3394.830 2471.420 3394.970 ;
        RECT 2470.360 3380.950 2470.500 3394.830 ;
        RECT 2470.300 3380.630 2470.560 3380.950 ;
        RECT 2470.760 3332.690 2471.020 3333.010 ;
        RECT 2470.820 3315.670 2470.960 3332.690 ;
        RECT 1318.000 3315.350 1318.260 3315.670 ;
        RECT 2470.760 3315.350 2471.020 3315.670 ;
        RECT 1318.060 3300.000 1318.200 3315.350 ;
        RECT 1318.000 3296.000 1318.280 3300.000 ;
      LAYER via2 ;
        RECT 2474.430 3430.120 2474.710 3430.400 ;
        RECT 2471.210 3429.440 2471.490 3429.720 ;
      LAYER met3 ;
        RECT 2474.405 3430.410 2474.735 3430.425 ;
        RECT 2470.510 3430.110 2474.735 3430.410 ;
        RECT 2470.510 3429.730 2470.810 3430.110 ;
        RECT 2474.405 3430.095 2474.735 3430.110 ;
        RECT 2471.185 3429.730 2471.515 3429.745 ;
        RECT 2470.510 3429.430 2471.515 3429.730 ;
        RECT 2471.185 3429.415 2471.515 3429.430 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1380.990 3315.920 1381.310 3315.980 ;
        RECT 2146.430 3315.920 2146.750 3315.980 ;
        RECT 1380.990 3315.780 2146.750 3315.920 ;
        RECT 1380.990 3315.720 1381.310 3315.780 ;
        RECT 2146.430 3315.720 2146.750 3315.780 ;
      LAYER via ;
        RECT 1381.020 3315.720 1381.280 3315.980 ;
        RECT 2146.460 3315.720 2146.720 3315.980 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3444.610 2149.420 3517.600 ;
        RECT 2147.900 3444.470 2149.420 3444.610 ;
        RECT 2147.900 3443.250 2148.040 3444.470 ;
        RECT 2147.440 3443.110 2148.040 3443.250 ;
        RECT 2147.440 3346.690 2147.580 3443.110 ;
        RECT 2146.520 3346.550 2147.580 3346.690 ;
        RECT 2146.520 3316.010 2146.660 3346.550 ;
        RECT 1381.020 3315.690 1381.280 3316.010 ;
        RECT 2146.460 3315.690 2146.720 3316.010 ;
        RECT 1381.080 3300.000 1381.220 3315.690 ;
        RECT 1381.020 3296.000 1381.300 3300.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1821.670 3464.160 1821.990 3464.220 ;
        RECT 1825.350 3464.160 1825.670 3464.220 ;
        RECT 1821.670 3464.020 1825.670 3464.160 ;
        RECT 1821.670 3463.960 1821.990 3464.020 ;
        RECT 1825.350 3463.960 1825.670 3464.020 ;
        RECT 1821.670 3415.540 1821.990 3415.600 ;
        RECT 1823.050 3415.540 1823.370 3415.600 ;
        RECT 1821.670 3415.400 1823.370 3415.540 ;
        RECT 1821.670 3415.340 1821.990 3415.400 ;
        RECT 1823.050 3415.340 1823.370 3415.400 ;
        RECT 1821.670 3367.940 1821.990 3368.000 ;
        RECT 1823.050 3367.940 1823.370 3368.000 ;
        RECT 1821.670 3367.800 1823.370 3367.940 ;
        RECT 1821.670 3367.740 1821.990 3367.800 ;
        RECT 1823.050 3367.740 1823.370 3367.800 ;
        RECT 1821.670 3343.120 1821.990 3343.180 ;
        RECT 1822.590 3343.120 1822.910 3343.180 ;
        RECT 1821.670 3342.980 1822.910 3343.120 ;
        RECT 1821.670 3342.920 1821.990 3342.980 ;
        RECT 1822.590 3342.920 1822.910 3342.980 ;
        RECT 1444.470 3316.600 1444.790 3316.660 ;
        RECT 1822.590 3316.600 1822.910 3316.660 ;
        RECT 1444.470 3316.460 1822.910 3316.600 ;
        RECT 1444.470 3316.400 1444.790 3316.460 ;
        RECT 1822.590 3316.400 1822.910 3316.460 ;
      LAYER via ;
        RECT 1821.700 3463.960 1821.960 3464.220 ;
        RECT 1825.380 3463.960 1825.640 3464.220 ;
        RECT 1821.700 3415.340 1821.960 3415.600 ;
        RECT 1823.080 3415.340 1823.340 3415.600 ;
        RECT 1821.700 3367.740 1821.960 3368.000 ;
        RECT 1823.080 3367.740 1823.340 3368.000 ;
        RECT 1821.700 3342.920 1821.960 3343.180 ;
        RECT 1822.620 3342.920 1822.880 3343.180 ;
        RECT 1444.500 3316.400 1444.760 3316.660 ;
        RECT 1822.620 3316.400 1822.880 3316.660 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3517.370 1825.120 3517.600 ;
        RECT 1824.980 3517.230 1825.580 3517.370 ;
        RECT 1825.440 3464.250 1825.580 3517.230 ;
        RECT 1821.700 3463.930 1821.960 3464.250 ;
        RECT 1825.380 3463.930 1825.640 3464.250 ;
        RECT 1821.760 3415.630 1821.900 3463.930 ;
        RECT 1821.700 3415.310 1821.960 3415.630 ;
        RECT 1823.080 3415.310 1823.340 3415.630 ;
        RECT 1823.140 3368.030 1823.280 3415.310 ;
        RECT 1821.700 3367.710 1821.960 3368.030 ;
        RECT 1823.080 3367.710 1823.340 3368.030 ;
        RECT 1821.760 3343.210 1821.900 3367.710 ;
        RECT 1821.700 3342.890 1821.960 3343.210 ;
        RECT 1822.620 3342.890 1822.880 3343.210 ;
        RECT 1822.680 3316.690 1822.820 3342.890 ;
        RECT 1444.500 3316.370 1444.760 3316.690 ;
        RECT 1822.620 3316.370 1822.880 3316.690 ;
        RECT 1444.560 3300.000 1444.700 3316.370 ;
        RECT 1444.500 3296.000 1444.780 3300.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3499.180 1500.910 3499.240 ;
        RECT 1503.810 3499.180 1504.130 3499.240 ;
        RECT 1500.590 3499.040 1504.130 3499.180 ;
        RECT 1500.590 3498.980 1500.910 3499.040 ;
        RECT 1503.810 3498.980 1504.130 3499.040 ;
        RECT 1503.810 3314.220 1504.130 3314.280 ;
        RECT 1507.490 3314.220 1507.810 3314.280 ;
        RECT 1503.810 3314.080 1507.810 3314.220 ;
        RECT 1503.810 3314.020 1504.130 3314.080 ;
        RECT 1507.490 3314.020 1507.810 3314.080 ;
      LAYER via ;
        RECT 1500.620 3498.980 1500.880 3499.240 ;
        RECT 1503.840 3498.980 1504.100 3499.240 ;
        RECT 1503.840 3314.020 1504.100 3314.280 ;
        RECT 1507.520 3314.020 1507.780 3314.280 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3499.270 1500.820 3517.600 ;
        RECT 1500.620 3498.950 1500.880 3499.270 ;
        RECT 1503.840 3498.950 1504.100 3499.270 ;
        RECT 1503.900 3314.310 1504.040 3498.950 ;
        RECT 1503.840 3313.990 1504.100 3314.310 ;
        RECT 1507.520 3313.990 1507.780 3314.310 ;
        RECT 1507.580 3300.000 1507.720 3313.990 ;
        RECT 1507.520 3296.000 1507.800 3300.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2695.210 324.260 2695.530 324.320 ;
        RECT 2898.070 324.260 2898.390 324.320 ;
        RECT 2695.210 324.120 2898.390 324.260 ;
        RECT 2695.210 324.060 2695.530 324.120 ;
        RECT 2898.070 324.060 2898.390 324.120 ;
      LAYER via ;
        RECT 2695.240 324.060 2695.500 324.320 ;
        RECT 2898.100 324.060 2898.360 324.320 ;
      LAYER met2 ;
        RECT 370.860 3299.770 371.140 3300.000 ;
        RECT 371.770 3299.770 372.050 3299.885 ;
        RECT 370.860 3299.630 372.050 3299.770 ;
        RECT 370.860 3296.000 371.140 3299.630 ;
        RECT 371.770 3299.515 372.050 3299.630 ;
        RECT 2695.230 3299.515 2695.510 3299.885 ;
        RECT 2695.300 324.350 2695.440 3299.515 ;
        RECT 2695.240 324.030 2695.500 324.350 ;
        RECT 2898.100 324.030 2898.360 324.350 ;
        RECT 2898.160 322.845 2898.300 324.030 ;
        RECT 2898.090 322.475 2898.370 322.845 ;
      LAYER via2 ;
        RECT 371.770 3299.560 372.050 3299.840 ;
        RECT 2695.230 3299.560 2695.510 3299.840 ;
        RECT 2898.090 322.520 2898.370 322.800 ;
      LAYER met3 ;
        RECT 371.745 3299.850 372.075 3299.865 ;
        RECT 2695.205 3299.850 2695.535 3299.865 ;
        RECT 371.745 3299.550 2695.535 3299.850 ;
        RECT 371.745 3299.535 372.075 3299.550 ;
        RECT 2695.205 3299.535 2695.535 3299.550 ;
        RECT 2898.065 322.810 2898.395 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.065 322.510 2924.800 322.810 ;
        RECT 2898.065 322.495 2898.395 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1179.510 3316.260 1179.830 3316.320 ;
        RECT 1570.510 3316.260 1570.830 3316.320 ;
        RECT 1179.510 3316.120 1570.830 3316.260 ;
        RECT 1179.510 3316.060 1179.830 3316.120 ;
        RECT 1570.510 3316.060 1570.830 3316.120 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1179.540 3316.060 1179.800 3316.320 ;
        RECT 1570.540 3316.060 1570.800 3316.320 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 3316.350 1179.740 3498.270 ;
        RECT 1179.540 3316.030 1179.800 3316.350 ;
        RECT 1570.540 3316.030 1570.800 3316.350 ;
        RECT 1570.600 3300.000 1570.740 3316.030 ;
        RECT 1570.540 3296.000 1570.820 3300.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3501.220 851.850 3501.280 ;
        RECT 1628.470 3501.220 1628.790 3501.280 ;
        RECT 851.530 3501.080 1628.790 3501.220 ;
        RECT 851.530 3501.020 851.850 3501.080 ;
        RECT 1628.470 3501.020 1628.790 3501.080 ;
      LAYER via ;
        RECT 851.560 3501.020 851.820 3501.280 ;
        RECT 1628.500 3501.020 1628.760 3501.280 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3501.310 851.760 3517.600 ;
        RECT 851.560 3500.990 851.820 3501.310 ;
        RECT 1628.500 3500.990 1628.760 3501.310 ;
        RECT 1628.560 3300.450 1628.700 3500.990 ;
        RECT 1628.560 3300.310 1631.460 3300.450 ;
        RECT 1631.320 3299.090 1631.460 3300.310 ;
        RECT 1634.020 3299.090 1634.300 3300.000 ;
        RECT 1631.320 3298.950 1634.300 3299.090 ;
        RECT 1634.020 3296.000 1634.300 3298.950 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3503.600 527.550 3503.660 ;
        RECT 1690.570 3503.600 1690.890 3503.660 ;
        RECT 527.230 3503.460 1690.890 3503.600 ;
        RECT 527.230 3503.400 527.550 3503.460 ;
        RECT 1690.570 3503.400 1690.890 3503.460 ;
      LAYER via ;
        RECT 527.260 3503.400 527.520 3503.660 ;
        RECT 1690.600 3503.400 1690.860 3503.660 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3503.690 527.460 3517.600 ;
        RECT 527.260 3503.370 527.520 3503.690 ;
        RECT 1690.600 3503.370 1690.860 3503.690 ;
        RECT 1690.660 3300.450 1690.800 3503.370 ;
        RECT 1690.660 3300.310 1694.940 3300.450 ;
        RECT 1694.800 3299.090 1694.940 3300.310 ;
        RECT 1697.040 3299.090 1697.320 3300.000 ;
        RECT 1694.800 3298.950 1697.320 3299.090 ;
        RECT 1697.040 3296.000 1697.320 3298.950 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 1759.570 3501.900 1759.890 3501.960 ;
        RECT 202.470 3501.760 1759.890 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 1759.570 3501.700 1759.890 3501.760 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 1759.600 3501.700 1759.860 3501.960 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 1759.600 3501.670 1759.860 3501.990 ;
        RECT 1759.660 3299.770 1759.800 3501.670 ;
        RECT 1760.060 3299.770 1760.340 3300.000 ;
        RECT 1759.660 3299.630 1760.340 3299.770 ;
        RECT 1760.060 3296.000 1760.340 3299.630 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 1822.130 3408.740 1822.450 3408.800 ;
        RECT 17.550 3408.600 1822.450 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 1822.130 3408.540 1822.450 3408.600 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 1822.160 3408.540 1822.420 3408.800 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 1822.160 3408.510 1822.420 3408.830 ;
        RECT 1822.220 3299.770 1822.360 3408.510 ;
        RECT 1823.080 3299.770 1823.360 3300.000 ;
        RECT 1822.220 3299.630 1823.360 3299.770 ;
        RECT 1823.080 3296.000 1823.360 3299.630 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 41.010 3303.680 41.330 3303.740 ;
        RECT 1886.530 3303.680 1886.850 3303.740 ;
        RECT 41.010 3303.540 1886.850 3303.680 ;
        RECT 41.010 3303.480 41.330 3303.540 ;
        RECT 1886.530 3303.480 1886.850 3303.540 ;
        RECT 15.710 3124.500 16.030 3124.560 ;
        RECT 41.010 3124.500 41.330 3124.560 ;
        RECT 15.710 3124.360 41.330 3124.500 ;
        RECT 15.710 3124.300 16.030 3124.360 ;
        RECT 41.010 3124.300 41.330 3124.360 ;
      LAYER via ;
        RECT 41.040 3303.480 41.300 3303.740 ;
        RECT 1886.560 3303.480 1886.820 3303.740 ;
        RECT 15.740 3124.300 16.000 3124.560 ;
        RECT 41.040 3124.300 41.300 3124.560 ;
      LAYER met2 ;
        RECT 41.040 3303.450 41.300 3303.770 ;
        RECT 1886.560 3303.450 1886.820 3303.770 ;
        RECT 41.100 3124.590 41.240 3303.450 ;
        RECT 1886.620 3300.000 1886.760 3303.450 ;
        RECT 1886.560 3296.000 1886.840 3300.000 ;
        RECT 15.740 3124.445 16.000 3124.590 ;
        RECT 15.730 3124.075 16.010 3124.445 ;
        RECT 41.040 3124.270 41.300 3124.590 ;
      LAYER via2 ;
        RECT 15.730 3124.120 16.010 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 15.705 3124.410 16.035 3124.425 ;
        RECT -4.800 3124.110 16.035 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 15.705 3124.095 16.035 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 40.550 3303.340 40.870 3303.400 ;
        RECT 1949.550 3303.340 1949.870 3303.400 ;
        RECT 40.550 3303.200 1949.870 3303.340 ;
        RECT 40.550 3303.140 40.870 3303.200 ;
        RECT 1949.550 3303.140 1949.870 3303.200 ;
        RECT 15.710 2837.880 16.030 2837.940 ;
        RECT 40.550 2837.880 40.870 2837.940 ;
        RECT 15.710 2837.740 40.870 2837.880 ;
        RECT 15.710 2837.680 16.030 2837.740 ;
        RECT 40.550 2837.680 40.870 2837.740 ;
      LAYER via ;
        RECT 40.580 3303.140 40.840 3303.400 ;
        RECT 1949.580 3303.140 1949.840 3303.400 ;
        RECT 15.740 2837.680 16.000 2837.940 ;
        RECT 40.580 2837.680 40.840 2837.940 ;
      LAYER met2 ;
        RECT 40.580 3303.110 40.840 3303.430 ;
        RECT 1949.580 3303.110 1949.840 3303.430 ;
        RECT 40.640 2837.970 40.780 3303.110 ;
        RECT 1949.640 3300.000 1949.780 3303.110 ;
        RECT 1949.580 3296.000 1949.860 3300.000 ;
        RECT 15.740 2837.650 16.000 2837.970 ;
        RECT 40.580 2837.650 40.840 2837.970 ;
        RECT 15.800 2836.805 15.940 2837.650 ;
        RECT 15.730 2836.435 16.010 2836.805 ;
      LAYER via2 ;
        RECT 15.730 2836.480 16.010 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 15.705 2836.770 16.035 2836.785 ;
        RECT -4.800 2836.470 16.035 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 15.705 2836.455 16.035 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 40.090 3302.660 40.410 3302.720 ;
        RECT 2012.570 3302.660 2012.890 3302.720 ;
        RECT 40.090 3302.520 2012.890 3302.660 ;
        RECT 40.090 3302.460 40.410 3302.520 ;
        RECT 2012.570 3302.460 2012.890 3302.520 ;
        RECT 16.170 2550.240 16.490 2550.300 ;
        RECT 40.090 2550.240 40.410 2550.300 ;
        RECT 16.170 2550.100 40.410 2550.240 ;
        RECT 16.170 2550.040 16.490 2550.100 ;
        RECT 40.090 2550.040 40.410 2550.100 ;
      LAYER via ;
        RECT 40.120 3302.460 40.380 3302.720 ;
        RECT 2012.600 3302.460 2012.860 3302.720 ;
        RECT 16.200 2550.040 16.460 2550.300 ;
        RECT 40.120 2550.040 40.380 2550.300 ;
      LAYER met2 ;
        RECT 40.120 3302.430 40.380 3302.750 ;
        RECT 2012.600 3302.430 2012.860 3302.750 ;
        RECT 40.180 2550.330 40.320 3302.430 ;
        RECT 2012.660 3300.000 2012.800 3302.430 ;
        RECT 2012.600 3296.000 2012.880 3300.000 ;
        RECT 16.200 2550.010 16.460 2550.330 ;
        RECT 40.120 2550.010 40.380 2550.330 ;
        RECT 16.260 2549.845 16.400 2550.010 ;
        RECT 16.190 2549.475 16.470 2549.845 ;
      LAYER via2 ;
        RECT 16.190 2549.520 16.470 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 16.165 2549.810 16.495 2549.825 ;
        RECT -4.800 2549.510 16.495 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 16.165 2549.495 16.495 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 39.630 3302.320 39.950 3302.380 ;
        RECT 2076.050 3302.320 2076.370 3302.380 ;
        RECT 39.630 3302.180 2076.370 3302.320 ;
        RECT 39.630 3302.120 39.950 3302.180 ;
        RECT 2076.050 3302.120 2076.370 3302.180 ;
        RECT 16.170 2262.260 16.490 2262.320 ;
        RECT 39.630 2262.260 39.950 2262.320 ;
        RECT 16.170 2262.120 39.950 2262.260 ;
        RECT 16.170 2262.060 16.490 2262.120 ;
        RECT 39.630 2262.060 39.950 2262.120 ;
      LAYER via ;
        RECT 39.660 3302.120 39.920 3302.380 ;
        RECT 2076.080 3302.120 2076.340 3302.380 ;
        RECT 16.200 2262.060 16.460 2262.320 ;
        RECT 39.660 2262.060 39.920 2262.320 ;
      LAYER met2 ;
        RECT 39.660 3302.090 39.920 3302.410 ;
        RECT 2076.080 3302.090 2076.340 3302.410 ;
        RECT 39.720 2262.350 39.860 3302.090 ;
        RECT 2076.140 3300.000 2076.280 3302.090 ;
        RECT 2076.080 3296.000 2076.360 3300.000 ;
        RECT 16.200 2262.205 16.460 2262.350 ;
        RECT 16.190 2261.835 16.470 2262.205 ;
        RECT 39.660 2262.030 39.920 2262.350 ;
      LAYER via2 ;
        RECT 16.190 2261.880 16.470 2262.160 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 16.165 2262.170 16.495 2262.185 ;
        RECT -4.800 2261.870 16.495 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 16.165 2261.855 16.495 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 39.170 3300.620 39.490 3300.680 ;
        RECT 2139.070 3300.620 2139.390 3300.680 ;
        RECT 39.170 3300.480 2139.390 3300.620 ;
        RECT 39.170 3300.420 39.490 3300.480 ;
        RECT 2139.070 3300.420 2139.390 3300.480 ;
        RECT 16.630 1976.320 16.950 1976.380 ;
        RECT 39.170 1976.320 39.490 1976.380 ;
        RECT 16.630 1976.180 39.490 1976.320 ;
        RECT 16.630 1976.120 16.950 1976.180 ;
        RECT 39.170 1976.120 39.490 1976.180 ;
      LAYER via ;
        RECT 39.200 3300.420 39.460 3300.680 ;
        RECT 2139.100 3300.420 2139.360 3300.680 ;
        RECT 16.660 1976.120 16.920 1976.380 ;
        RECT 39.200 1976.120 39.460 1976.380 ;
      LAYER met2 ;
        RECT 39.200 3300.390 39.460 3300.710 ;
        RECT 2139.100 3300.390 2139.360 3300.710 ;
        RECT 39.260 1976.410 39.400 3300.390 ;
        RECT 2139.160 3300.000 2139.300 3300.390 ;
        RECT 2139.100 3296.000 2139.380 3300.000 ;
        RECT 16.660 1976.090 16.920 1976.410 ;
        RECT 39.200 1976.090 39.460 1976.410 ;
        RECT 16.720 1975.245 16.860 1976.090 ;
        RECT 16.650 1974.875 16.930 1975.245 ;
      LAYER via2 ;
        RECT 16.650 1974.920 16.930 1975.200 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 16.625 1975.210 16.955 1975.225 ;
        RECT -4.800 1974.910 16.955 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 16.625 1974.895 16.955 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2696.130 558.860 2696.450 558.920 ;
        RECT 2900.830 558.860 2901.150 558.920 ;
        RECT 2696.130 558.720 2901.150 558.860 ;
        RECT 2696.130 558.660 2696.450 558.720 ;
        RECT 2900.830 558.660 2901.150 558.720 ;
      LAYER via ;
        RECT 2696.160 558.660 2696.420 558.920 ;
        RECT 2900.860 558.660 2901.120 558.920 ;
      LAYER met2 ;
        RECT 433.870 3300.195 434.150 3300.565 ;
        RECT 2696.150 3300.195 2696.430 3300.565 ;
        RECT 433.940 3300.000 434.080 3300.195 ;
        RECT 433.880 3296.000 434.160 3300.000 ;
        RECT 2696.220 558.950 2696.360 3300.195 ;
        RECT 2696.160 558.630 2696.420 558.950 ;
        RECT 2900.860 558.630 2901.120 558.950 ;
        RECT 2900.920 557.445 2901.060 558.630 ;
        RECT 2900.850 557.075 2901.130 557.445 ;
      LAYER via2 ;
        RECT 433.870 3300.240 434.150 3300.520 ;
        RECT 2696.150 3300.240 2696.430 3300.520 ;
        RECT 2900.850 557.120 2901.130 557.400 ;
      LAYER met3 ;
        RECT 433.845 3300.530 434.175 3300.545 ;
        RECT 2696.125 3300.530 2696.455 3300.545 ;
        RECT 433.845 3300.230 2696.455 3300.530 ;
        RECT 433.845 3300.215 434.175 3300.230 ;
        RECT 2696.125 3300.215 2696.455 3300.230 ;
        RECT 2900.825 557.410 2901.155 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2900.825 557.110 2924.800 557.410 ;
        RECT 2900.825 557.095 2901.155 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.710 3300.280 39.030 3300.340 ;
        RECT 2201.170 3300.280 2201.490 3300.340 ;
        RECT 38.710 3300.140 2201.490 3300.280 ;
        RECT 38.710 3300.080 39.030 3300.140 ;
        RECT 2201.170 3300.080 2201.490 3300.140 ;
        RECT 16.630 1687.660 16.950 1687.720 ;
        RECT 38.710 1687.660 39.030 1687.720 ;
        RECT 16.630 1687.520 39.030 1687.660 ;
        RECT 16.630 1687.460 16.950 1687.520 ;
        RECT 38.710 1687.460 39.030 1687.520 ;
      LAYER via ;
        RECT 38.740 3300.080 39.000 3300.340 ;
        RECT 2201.200 3300.080 2201.460 3300.340 ;
        RECT 16.660 1687.460 16.920 1687.720 ;
        RECT 38.740 1687.460 39.000 1687.720 ;
      LAYER met2 ;
        RECT 38.740 3300.050 39.000 3300.370 ;
        RECT 2201.200 3300.050 2201.460 3300.370 ;
        RECT 38.800 1687.750 38.940 3300.050 ;
        RECT 2201.260 3299.770 2201.400 3300.050 ;
        RECT 2202.120 3299.770 2202.400 3300.000 ;
        RECT 2201.260 3299.630 2202.400 3299.770 ;
        RECT 2202.120 3296.000 2202.400 3299.630 ;
        RECT 16.660 1687.605 16.920 1687.750 ;
        RECT 16.650 1687.235 16.930 1687.605 ;
        RECT 38.740 1687.430 39.000 1687.750 ;
      LAYER via2 ;
        RECT 16.650 1687.280 16.930 1687.560 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 16.625 1687.570 16.955 1687.585 ;
        RECT -4.800 1687.270 16.955 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 16.625 1687.255 16.955 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 3299.600 38.570 3299.660 ;
        RECT 2263.270 3299.600 2263.590 3299.660 ;
        RECT 38.250 3299.460 2263.590 3299.600 ;
        RECT 38.250 3299.400 38.570 3299.460 ;
        RECT 2263.270 3299.400 2263.590 3299.460 ;
        RECT 15.710 1474.140 16.030 1474.200 ;
        RECT 38.250 1474.140 38.570 1474.200 ;
        RECT 15.710 1474.000 38.570 1474.140 ;
        RECT 15.710 1473.940 16.030 1474.000 ;
        RECT 38.250 1473.940 38.570 1474.000 ;
      LAYER via ;
        RECT 38.280 3299.400 38.540 3299.660 ;
        RECT 2263.300 3299.400 2263.560 3299.660 ;
        RECT 15.740 1473.940 16.000 1474.200 ;
        RECT 38.280 1473.940 38.540 1474.200 ;
      LAYER met2 ;
        RECT 2265.140 3299.770 2265.420 3300.000 ;
        RECT 2263.360 3299.690 2265.420 3299.770 ;
        RECT 38.280 3299.370 38.540 3299.690 ;
        RECT 2263.300 3299.630 2265.420 3299.690 ;
        RECT 2263.300 3299.370 2263.560 3299.630 ;
        RECT 38.340 1474.230 38.480 3299.370 ;
        RECT 2265.140 3296.000 2265.420 3299.630 ;
        RECT 15.740 1473.910 16.000 1474.230 ;
        RECT 38.280 1473.910 38.540 1474.230 ;
        RECT 15.800 1472.045 15.940 1473.910 ;
        RECT 15.730 1471.675 16.010 1472.045 ;
      LAYER via2 ;
        RECT 15.730 1471.720 16.010 1472.000 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 15.705 1472.010 16.035 1472.025 ;
        RECT -4.800 1471.710 16.035 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 15.705 1471.695 16.035 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 37.790 3299.260 38.110 3299.320 ;
        RECT 2326.750 3299.260 2327.070 3299.320 ;
        RECT 37.790 3299.120 2327.070 3299.260 ;
        RECT 37.790 3299.060 38.110 3299.120 ;
        RECT 2326.750 3299.060 2327.070 3299.120 ;
        RECT 16.630 1261.300 16.950 1261.360 ;
        RECT 37.790 1261.300 38.110 1261.360 ;
        RECT 16.630 1261.160 38.110 1261.300 ;
        RECT 16.630 1261.100 16.950 1261.160 ;
        RECT 37.790 1261.100 38.110 1261.160 ;
      LAYER via ;
        RECT 37.820 3299.060 38.080 3299.320 ;
        RECT 2326.780 3299.060 2327.040 3299.320 ;
        RECT 16.660 1261.100 16.920 1261.360 ;
        RECT 37.820 1261.100 38.080 1261.360 ;
      LAYER met2 ;
        RECT 37.820 3299.030 38.080 3299.350 ;
        RECT 2326.780 3299.090 2327.040 3299.350 ;
        RECT 2328.620 3299.090 2328.900 3300.000 ;
        RECT 2326.780 3299.030 2328.900 3299.090 ;
        RECT 37.880 1261.390 38.020 3299.030 ;
        RECT 2326.840 3298.950 2328.900 3299.030 ;
        RECT 2328.620 3296.000 2328.900 3298.950 ;
        RECT 16.660 1261.070 16.920 1261.390 ;
        RECT 37.820 1261.070 38.080 1261.390 ;
        RECT 16.720 1256.485 16.860 1261.070 ;
        RECT 16.650 1256.115 16.930 1256.485 ;
      LAYER via2 ;
        RECT 16.650 1256.160 16.930 1256.440 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 16.625 1256.450 16.955 1256.465 ;
        RECT -4.800 1256.150 16.955 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 16.625 1256.135 16.955 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 46.070 3298.920 46.390 3298.980 ;
        RECT 2390.230 3298.920 2390.550 3298.980 ;
        RECT 46.070 3298.780 2390.550 3298.920 ;
        RECT 46.070 3298.720 46.390 3298.780 ;
        RECT 2390.230 3298.720 2390.550 3298.780 ;
        RECT 16.630 1040.980 16.950 1041.040 ;
        RECT 46.070 1040.980 46.390 1041.040 ;
        RECT 16.630 1040.840 46.390 1040.980 ;
        RECT 16.630 1040.780 16.950 1040.840 ;
        RECT 46.070 1040.780 46.390 1040.840 ;
      LAYER via ;
        RECT 46.100 3298.720 46.360 3298.980 ;
        RECT 2390.260 3298.720 2390.520 3298.980 ;
        RECT 16.660 1040.780 16.920 1041.040 ;
        RECT 46.100 1040.780 46.360 1041.040 ;
      LAYER met2 ;
        RECT 2391.640 3299.090 2391.920 3300.000 ;
        RECT 2390.320 3299.010 2391.920 3299.090 ;
        RECT 46.100 3298.690 46.360 3299.010 ;
        RECT 2390.260 3298.950 2391.920 3299.010 ;
        RECT 2390.260 3298.690 2390.520 3298.950 ;
        RECT 46.160 1041.070 46.300 3298.690 ;
        RECT 2391.640 3296.000 2391.920 3298.950 ;
        RECT 16.660 1040.925 16.920 1041.070 ;
        RECT 16.650 1040.555 16.930 1040.925 ;
        RECT 46.100 1040.750 46.360 1041.070 ;
      LAYER via2 ;
        RECT 16.650 1040.600 16.930 1040.880 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 16.625 1040.890 16.955 1040.905 ;
        RECT -4.800 1040.590 16.955 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 16.625 1040.575 16.955 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 30.890 3298.580 31.210 3298.640 ;
        RECT 2452.790 3298.580 2453.110 3298.640 ;
        RECT 30.890 3298.440 2453.110 3298.580 ;
        RECT 30.890 3298.380 31.210 3298.440 ;
        RECT 2452.790 3298.380 2453.110 3298.440 ;
        RECT 15.250 827.460 15.570 827.520 ;
        RECT 30.890 827.460 31.210 827.520 ;
        RECT 15.250 827.320 31.210 827.460 ;
        RECT 15.250 827.260 15.570 827.320 ;
        RECT 30.890 827.260 31.210 827.320 ;
      LAYER via ;
        RECT 30.920 3298.380 31.180 3298.640 ;
        RECT 2452.820 3298.380 2453.080 3298.640 ;
        RECT 15.280 827.260 15.540 827.520 ;
        RECT 30.920 827.260 31.180 827.520 ;
      LAYER met2 ;
        RECT 30.920 3298.350 31.180 3298.670 ;
        RECT 2452.820 3298.410 2453.080 3298.670 ;
        RECT 2454.660 3298.410 2454.940 3300.000 ;
        RECT 2452.820 3298.350 2454.940 3298.410 ;
        RECT 30.980 827.550 31.120 3298.350 ;
        RECT 2452.880 3298.270 2454.940 3298.350 ;
        RECT 2454.660 3296.000 2454.940 3298.270 ;
        RECT 15.280 827.230 15.540 827.550 ;
        RECT 30.920 827.230 31.180 827.550 ;
        RECT 15.340 825.365 15.480 827.230 ;
        RECT 15.270 824.995 15.550 825.365 ;
      LAYER via2 ;
        RECT 15.270 825.040 15.550 825.320 ;
      LAYER met3 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 15.245 825.330 15.575 825.345 ;
        RECT -4.800 825.030 15.575 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 15.245 825.015 15.575 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 613.940 16.950 614.000 ;
        RECT 127.490 613.940 127.810 614.000 ;
        RECT 16.630 613.800 127.810 613.940 ;
        RECT 16.630 613.740 16.950 613.800 ;
        RECT 127.490 613.740 127.810 613.800 ;
      LAYER via ;
        RECT 16.660 613.740 16.920 614.000 ;
        RECT 127.520 613.740 127.780 614.000 ;
      LAYER met2 ;
        RECT 127.510 3298.835 127.790 3299.205 ;
        RECT 2516.290 3299.090 2516.570 3299.205 ;
        RECT 2518.140 3299.090 2518.420 3300.000 ;
        RECT 2516.290 3298.950 2518.420 3299.090 ;
        RECT 2516.290 3298.835 2516.570 3298.950 ;
        RECT 127.580 614.030 127.720 3298.835 ;
        RECT 2518.140 3296.000 2518.420 3298.950 ;
        RECT 16.660 613.710 16.920 614.030 ;
        RECT 127.520 613.710 127.780 614.030 ;
        RECT 16.720 610.485 16.860 613.710 ;
        RECT 16.650 610.115 16.930 610.485 ;
      LAYER via2 ;
        RECT 127.510 3298.880 127.790 3299.160 ;
        RECT 2516.290 3298.880 2516.570 3299.160 ;
        RECT 16.650 610.160 16.930 610.440 ;
      LAYER met3 ;
        RECT 127.485 3299.170 127.815 3299.185 ;
        RECT 2516.265 3299.170 2516.595 3299.185 ;
        RECT 127.485 3298.870 2516.595 3299.170 ;
        RECT 127.485 3298.855 127.815 3298.870 ;
        RECT 2516.265 3298.855 2516.595 3298.870 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 16.625 610.450 16.955 610.465 ;
        RECT -4.800 610.150 16.955 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 16.625 610.135 16.955 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 395.660 16.030 395.720 ;
        RECT 44.690 395.660 45.010 395.720 ;
        RECT 15.710 395.520 45.010 395.660 ;
        RECT 15.710 395.460 16.030 395.520 ;
        RECT 44.690 395.460 45.010 395.520 ;
      LAYER via ;
        RECT 15.740 395.460 16.000 395.720 ;
        RECT 44.720 395.460 44.980 395.720 ;
      LAYER met2 ;
        RECT 2580.690 3297.050 2580.970 3297.165 ;
        RECT 2581.160 3297.050 2581.440 3300.000 ;
        RECT 2580.690 3296.910 2581.440 3297.050 ;
        RECT 2580.690 3296.795 2580.970 3296.910 ;
        RECT 2581.160 3296.000 2581.440 3296.910 ;
        RECT 44.710 3291.355 44.990 3291.725 ;
        RECT 44.780 395.750 44.920 3291.355 ;
        RECT 15.740 395.430 16.000 395.750 ;
        RECT 44.720 395.430 44.980 395.750 ;
        RECT 15.800 394.925 15.940 395.430 ;
        RECT 15.730 394.555 16.010 394.925 ;
      LAYER via2 ;
        RECT 2580.690 3296.840 2580.970 3297.120 ;
        RECT 44.710 3291.400 44.990 3291.680 ;
        RECT 15.730 394.600 16.010 394.880 ;
      LAYER met3 ;
        RECT 2563.390 3297.130 2563.770 3297.140 ;
        RECT 2580.665 3297.130 2580.995 3297.145 ;
        RECT 2563.390 3296.830 2580.995 3297.130 ;
        RECT 2563.390 3296.820 2563.770 3296.830 ;
        RECT 2580.665 3296.815 2580.995 3296.830 ;
        RECT 44.685 3291.690 45.015 3291.705 ;
        RECT 2563.390 3291.690 2563.770 3291.700 ;
        RECT 44.685 3291.390 2563.770 3291.690 ;
        RECT 44.685 3291.375 45.015 3291.390 ;
        RECT 2563.390 3291.380 2563.770 3291.390 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 15.705 394.890 16.035 394.905 ;
        RECT -4.800 394.590 16.035 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 15.705 394.575 16.035 394.590 ;
      LAYER via3 ;
        RECT 2563.420 3296.820 2563.740 3297.140 ;
        RECT 2563.420 3291.380 2563.740 3291.700 ;
      LAYER met4 ;
        RECT 2563.415 3296.815 2563.745 3297.145 ;
        RECT 2563.430 3291.705 2563.730 3296.815 ;
        RECT 2563.415 3291.375 2563.745 3291.705 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2242.570 3306.400 2242.890 3306.460 ;
        RECT 2644.150 3306.400 2644.470 3306.460 ;
        RECT 2242.570 3306.260 2644.470 3306.400 ;
        RECT 2242.570 3306.200 2242.890 3306.260 ;
        RECT 2644.150 3306.200 2644.470 3306.260 ;
      LAYER via ;
        RECT 2242.600 3306.200 2242.860 3306.460 ;
        RECT 2644.180 3306.200 2644.440 3306.460 ;
      LAYER met2 ;
        RECT 2242.600 3306.170 2242.860 3306.490 ;
        RECT 2644.180 3306.170 2644.440 3306.490 ;
        RECT 2242.660 3297.165 2242.800 3306.170 ;
        RECT 2644.240 3300.000 2644.380 3306.170 ;
        RECT 2242.590 3296.795 2242.870 3297.165 ;
        RECT 2644.180 3296.000 2644.460 3300.000 ;
        RECT 17.570 3294.755 17.850 3295.125 ;
        RECT 17.640 179.365 17.780 3294.755 ;
        RECT 17.570 178.995 17.850 179.365 ;
      LAYER via2 ;
        RECT 2242.590 3296.840 2242.870 3297.120 ;
        RECT 17.570 3294.800 17.850 3295.080 ;
        RECT 17.570 179.040 17.850 179.320 ;
      LAYER met3 ;
        RECT 2232.190 3297.130 2232.570 3297.140 ;
        RECT 2242.565 3297.130 2242.895 3297.145 ;
        RECT 2232.190 3296.830 2242.895 3297.130 ;
        RECT 2232.190 3296.820 2232.570 3296.830 ;
        RECT 2242.565 3296.815 2242.895 3296.830 ;
        RECT 17.545 3295.090 17.875 3295.105 ;
        RECT 2232.190 3295.090 2232.570 3295.100 ;
        RECT 17.545 3294.790 2232.570 3295.090 ;
        RECT 17.545 3294.775 17.875 3294.790 ;
        RECT 2232.190 3294.780 2232.570 3294.790 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.545 179.330 17.875 179.345 ;
        RECT -4.800 179.030 17.875 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.545 179.015 17.875 179.030 ;
      LAYER via3 ;
        RECT 2232.220 3296.820 2232.540 3297.140 ;
        RECT 2232.220 3294.780 2232.540 3295.100 ;
      LAYER met4 ;
        RECT 2232.215 3296.815 2232.545 3297.145 ;
        RECT 2232.230 3295.105 2232.530 3296.815 ;
        RECT 2232.215 3294.775 2232.545 3295.105 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 498.250 3299.940 498.570 3300.000 ;
        RECT 2695.670 3299.940 2695.990 3300.000 ;
        RECT 498.250 3299.800 2695.990 3299.940 ;
        RECT 498.250 3299.740 498.570 3299.800 ;
        RECT 2695.670 3299.740 2695.990 3299.800 ;
        RECT 2695.670 793.460 2695.990 793.520 ;
        RECT 2900.830 793.460 2901.150 793.520 ;
        RECT 2695.670 793.320 2901.150 793.460 ;
        RECT 2695.670 793.260 2695.990 793.320 ;
        RECT 2900.830 793.260 2901.150 793.320 ;
      LAYER via ;
        RECT 498.280 3299.740 498.540 3300.000 ;
        RECT 2695.700 3299.740 2695.960 3300.000 ;
        RECT 2695.700 793.260 2695.960 793.520 ;
        RECT 2900.860 793.260 2901.120 793.520 ;
      LAYER met2 ;
        RECT 496.900 3299.770 497.180 3300.000 ;
        RECT 498.280 3299.770 498.540 3300.030 ;
        RECT 496.900 3299.710 498.540 3299.770 ;
        RECT 2695.700 3299.710 2695.960 3300.030 ;
        RECT 496.900 3299.630 498.480 3299.710 ;
        RECT 496.900 3296.000 497.180 3299.630 ;
        RECT 2695.760 793.550 2695.900 3299.710 ;
        RECT 2695.700 793.230 2695.960 793.550 ;
        RECT 2900.860 793.230 2901.120 793.550 ;
        RECT 2900.920 792.045 2901.060 793.230 ;
        RECT 2900.850 791.675 2901.130 792.045 ;
      LAYER via2 ;
        RECT 2900.850 791.720 2901.130 792.000 ;
      LAYER met3 ;
        RECT 2900.825 792.010 2901.155 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2900.825 791.710 2924.800 792.010 ;
        RECT 2900.825 791.695 2901.155 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1845.665 3295.705 1845.835 3298.255 ;
      LAYER mcon ;
        RECT 1845.665 3298.085 1845.835 3298.255 ;
      LAYER met1 ;
        RECT 560.350 3310.480 560.670 3310.540 ;
        RECT 1845.590 3310.480 1845.910 3310.540 ;
        RECT 560.350 3310.340 1845.910 3310.480 ;
        RECT 560.350 3310.280 560.670 3310.340 ;
        RECT 1845.590 3310.280 1845.910 3310.340 ;
        RECT 1845.590 3298.240 1845.910 3298.300 ;
        RECT 1845.395 3298.100 1845.910 3298.240 ;
        RECT 1845.590 3298.040 1845.910 3298.100 ;
        RECT 1845.605 3295.860 1845.895 3295.905 ;
        RECT 2904.050 3295.860 2904.370 3295.920 ;
        RECT 1845.605 3295.720 2904.370 3295.860 ;
        RECT 1845.605 3295.675 1845.895 3295.720 ;
        RECT 2904.050 3295.660 2904.370 3295.720 ;
      LAYER via ;
        RECT 560.380 3310.280 560.640 3310.540 ;
        RECT 1845.620 3310.280 1845.880 3310.540 ;
        RECT 1845.620 3298.040 1845.880 3298.300 ;
        RECT 2904.080 3295.660 2904.340 3295.920 ;
      LAYER met2 ;
        RECT 560.380 3310.250 560.640 3310.570 ;
        RECT 1845.620 3310.250 1845.880 3310.570 ;
        RECT 560.440 3300.000 560.580 3310.250 ;
        RECT 560.380 3296.000 560.660 3300.000 ;
        RECT 1845.680 3298.330 1845.820 3310.250 ;
        RECT 1845.620 3298.010 1845.880 3298.330 ;
        RECT 2904.080 3295.630 2904.340 3295.950 ;
        RECT 2904.140 1026.645 2904.280 3295.630 ;
        RECT 2904.070 1026.275 2904.350 1026.645 ;
      LAYER via2 ;
        RECT 2904.070 1026.320 2904.350 1026.600 ;
      LAYER met3 ;
        RECT 2904.045 1026.610 2904.375 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2904.045 1026.310 2924.800 1026.610 ;
        RECT 2904.045 1026.295 2904.375 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 625.285 3293.665 625.455 3296.555 ;
      LAYER mcon ;
        RECT 625.285 3296.385 625.455 3296.555 ;
      LAYER met1 ;
        RECT 625.210 3296.540 625.530 3296.600 ;
        RECT 625.015 3296.400 625.530 3296.540 ;
        RECT 625.210 3296.340 625.530 3296.400 ;
        RECT 625.225 3293.820 625.515 3293.865 ;
        RECT 2696.590 3293.820 2696.910 3293.880 ;
        RECT 625.225 3293.680 2696.910 3293.820 ;
        RECT 625.225 3293.635 625.515 3293.680 ;
        RECT 2696.590 3293.620 2696.910 3293.680 ;
        RECT 2696.590 1262.660 2696.910 1262.720 ;
        RECT 2900.830 1262.660 2901.150 1262.720 ;
        RECT 2696.590 1262.520 2901.150 1262.660 ;
        RECT 2696.590 1262.460 2696.910 1262.520 ;
        RECT 2900.830 1262.460 2901.150 1262.520 ;
      LAYER via ;
        RECT 625.240 3296.340 625.500 3296.600 ;
        RECT 2696.620 3293.620 2696.880 3293.880 ;
        RECT 2696.620 1262.460 2696.880 1262.720 ;
        RECT 2900.860 1262.460 2901.120 1262.720 ;
      LAYER met2 ;
        RECT 623.400 3296.370 623.680 3300.000 ;
        RECT 625.240 3296.370 625.500 3296.630 ;
        RECT 623.400 3296.310 625.500 3296.370 ;
        RECT 623.400 3296.230 625.440 3296.310 ;
        RECT 623.400 3296.000 623.680 3296.230 ;
        RECT 2696.620 3293.590 2696.880 3293.910 ;
        RECT 2696.680 1262.750 2696.820 3293.590 ;
        RECT 2696.620 1262.430 2696.880 1262.750 ;
        RECT 2900.860 1262.430 2901.120 1262.750 ;
        RECT 2900.920 1261.245 2901.060 1262.430 ;
        RECT 2900.850 1260.875 2901.130 1261.245 ;
      LAYER via2 ;
        RECT 2900.850 1260.920 2901.130 1261.200 ;
      LAYER met3 ;
        RECT 2900.825 1261.210 2901.155 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2900.825 1260.910 2924.800 1261.210 ;
        RECT 2900.825 1260.895 2901.155 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 687.845 3294.685 688.015 3296.555 ;
      LAYER mcon ;
        RECT 687.845 3296.385 688.015 3296.555 ;
      LAYER met1 ;
        RECT 687.770 3296.540 688.090 3296.600 ;
        RECT 687.575 3296.400 688.090 3296.540 ;
        RECT 687.770 3296.340 688.090 3296.400 ;
        RECT 687.785 3294.840 688.075 3294.885 ;
        RECT 2697.050 3294.840 2697.370 3294.900 ;
        RECT 687.785 3294.700 2697.370 3294.840 ;
        RECT 687.785 3294.655 688.075 3294.700 ;
        RECT 2697.050 3294.640 2697.370 3294.700 ;
        RECT 2697.050 1497.260 2697.370 1497.320 ;
        RECT 2900.830 1497.260 2901.150 1497.320 ;
        RECT 2697.050 1497.120 2901.150 1497.260 ;
        RECT 2697.050 1497.060 2697.370 1497.120 ;
        RECT 2900.830 1497.060 2901.150 1497.120 ;
      LAYER via ;
        RECT 687.800 3296.340 688.060 3296.600 ;
        RECT 2697.080 3294.640 2697.340 3294.900 ;
        RECT 2697.080 1497.060 2697.340 1497.320 ;
        RECT 2900.860 1497.060 2901.120 1497.320 ;
      LAYER met2 ;
        RECT 686.420 3296.370 686.700 3300.000 ;
        RECT 687.800 3296.370 688.060 3296.630 ;
        RECT 686.420 3296.310 688.060 3296.370 ;
        RECT 686.420 3296.230 688.000 3296.310 ;
        RECT 686.420 3296.000 686.700 3296.230 ;
        RECT 2697.080 3294.610 2697.340 3294.930 ;
        RECT 2697.140 1497.350 2697.280 3294.610 ;
        RECT 2697.080 1497.030 2697.340 1497.350 ;
        RECT 2900.860 1497.030 2901.120 1497.350 ;
        RECT 2900.920 1495.845 2901.060 1497.030 ;
        RECT 2900.850 1495.475 2901.130 1495.845 ;
      LAYER via2 ;
        RECT 2900.850 1495.520 2901.130 1495.800 ;
      LAYER met3 ;
        RECT 2900.825 1495.810 2901.155 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2900.825 1495.510 2924.800 1495.810 ;
        RECT 2900.825 1495.495 2901.155 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 749.870 3303.000 750.190 3303.060 ;
        RECT 2697.510 3303.000 2697.830 3303.060 ;
        RECT 749.870 3302.860 2697.830 3303.000 ;
        RECT 749.870 3302.800 750.190 3302.860 ;
        RECT 2697.510 3302.800 2697.830 3302.860 ;
        RECT 2697.510 1731.860 2697.830 1731.920 ;
        RECT 2900.830 1731.860 2901.150 1731.920 ;
        RECT 2697.510 1731.720 2901.150 1731.860 ;
        RECT 2697.510 1731.660 2697.830 1731.720 ;
        RECT 2900.830 1731.660 2901.150 1731.720 ;
      LAYER via ;
        RECT 749.900 3302.800 750.160 3303.060 ;
        RECT 2697.540 3302.800 2697.800 3303.060 ;
        RECT 2697.540 1731.660 2697.800 1731.920 ;
        RECT 2900.860 1731.660 2901.120 1731.920 ;
      LAYER met2 ;
        RECT 749.900 3302.770 750.160 3303.090 ;
        RECT 2697.540 3302.770 2697.800 3303.090 ;
        RECT 749.960 3300.000 750.100 3302.770 ;
        RECT 749.900 3296.000 750.180 3300.000 ;
        RECT 2697.600 1731.950 2697.740 3302.770 ;
        RECT 2697.540 1731.630 2697.800 1731.950 ;
        RECT 2900.860 1731.630 2901.120 1731.950 ;
        RECT 2900.920 1730.445 2901.060 1731.630 ;
        RECT 2900.850 1730.075 2901.130 1730.445 ;
      LAYER via2 ;
        RECT 2900.850 1730.120 2901.130 1730.400 ;
      LAYER met3 ;
        RECT 2900.825 1730.410 2901.155 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2900.825 1730.110 2924.800 1730.410 ;
        RECT 2900.825 1730.095 2901.155 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 812.890 3308.780 813.210 3308.840 ;
        RECT 2693.830 3308.780 2694.150 3308.840 ;
        RECT 812.890 3308.640 2694.150 3308.780 ;
        RECT 812.890 3308.580 813.210 3308.640 ;
        RECT 2693.830 3308.580 2694.150 3308.640 ;
        RECT 2693.830 1966.460 2694.150 1966.520 ;
        RECT 2900.830 1966.460 2901.150 1966.520 ;
        RECT 2693.830 1966.320 2901.150 1966.460 ;
        RECT 2693.830 1966.260 2694.150 1966.320 ;
        RECT 2900.830 1966.260 2901.150 1966.320 ;
      LAYER via ;
        RECT 812.920 3308.580 813.180 3308.840 ;
        RECT 2693.860 3308.580 2694.120 3308.840 ;
        RECT 2693.860 1966.260 2694.120 1966.520 ;
        RECT 2900.860 1966.260 2901.120 1966.520 ;
      LAYER met2 ;
        RECT 812.920 3308.550 813.180 3308.870 ;
        RECT 2693.860 3308.550 2694.120 3308.870 ;
        RECT 812.980 3300.000 813.120 3308.550 ;
        RECT 812.920 3296.000 813.200 3300.000 ;
        RECT 2693.920 1966.550 2694.060 3308.550 ;
        RECT 2693.860 1966.230 2694.120 1966.550 ;
        RECT 2900.860 1966.230 2901.120 1966.550 ;
        RECT 2900.920 1965.045 2901.060 1966.230 ;
        RECT 2900.850 1964.675 2901.130 1965.045 ;
      LAYER via2 ;
        RECT 2900.850 1964.720 2901.130 1965.000 ;
      LAYER met3 ;
        RECT 2900.825 1965.010 2901.155 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2900.825 1964.710 2924.800 1965.010 ;
        RECT 2900.825 1964.695 2901.155 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 875.910 3312.520 876.230 3312.580 ;
        RECT 2887.490 3312.520 2887.810 3312.580 ;
        RECT 875.910 3312.380 2887.810 3312.520 ;
        RECT 875.910 3312.320 876.230 3312.380 ;
        RECT 2887.490 3312.320 2887.810 3312.380 ;
        RECT 2887.490 2201.060 2887.810 2201.120 ;
        RECT 2898.530 2201.060 2898.850 2201.120 ;
        RECT 2887.490 2200.920 2898.850 2201.060 ;
        RECT 2887.490 2200.860 2887.810 2200.920 ;
        RECT 2898.530 2200.860 2898.850 2200.920 ;
      LAYER via ;
        RECT 875.940 3312.320 876.200 3312.580 ;
        RECT 2887.520 3312.320 2887.780 3312.580 ;
        RECT 2887.520 2200.860 2887.780 2201.120 ;
        RECT 2898.560 2200.860 2898.820 2201.120 ;
      LAYER met2 ;
        RECT 875.940 3312.290 876.200 3312.610 ;
        RECT 2887.520 3312.290 2887.780 3312.610 ;
        RECT 876.000 3300.000 876.140 3312.290 ;
        RECT 875.940 3296.000 876.220 3300.000 ;
        RECT 2887.580 2201.150 2887.720 3312.290 ;
        RECT 2887.520 2200.830 2887.780 2201.150 ;
        RECT 2898.560 2200.830 2898.820 2201.150 ;
        RECT 2898.620 2199.645 2898.760 2200.830 ;
        RECT 2898.550 2199.275 2898.830 2199.645 ;
      LAYER via2 ;
        RECT 2898.550 2199.320 2898.830 2199.600 ;
      LAYER met3 ;
        RECT 2898.525 2199.610 2898.855 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2898.525 2199.310 2924.800 2199.610 ;
        RECT 2898.525 2199.295 2898.855 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 328.530 3306.995 328.810 3307.365 ;
        RECT 2902.230 3306.995 2902.510 3307.365 ;
        RECT 328.600 3300.000 328.740 3306.995 ;
        RECT 328.540 3296.000 328.820 3300.000 ;
        RECT 2902.300 205.205 2902.440 3306.995 ;
        RECT 2902.230 204.835 2902.510 205.205 ;
      LAYER via2 ;
        RECT 328.530 3307.040 328.810 3307.320 ;
        RECT 2902.230 3307.040 2902.510 3307.320 ;
        RECT 2902.230 204.880 2902.510 205.160 ;
      LAYER met3 ;
        RECT 328.505 3307.330 328.835 3307.345 ;
        RECT 2902.205 3307.330 2902.535 3307.345 ;
        RECT 328.505 3307.030 2902.535 3307.330 ;
        RECT 328.505 3307.015 328.835 3307.030 ;
        RECT 2902.205 3307.015 2902.535 3307.030 ;
        RECT 2902.205 205.170 2902.535 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2902.205 204.870 2924.800 205.170 ;
        RECT 2902.205 204.855 2902.535 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 960.090 3313.540 960.410 3313.600 ;
        RECT 2699.810 3313.540 2700.130 3313.600 ;
        RECT 960.090 3313.400 2700.130 3313.540 ;
        RECT 960.090 3313.340 960.410 3313.400 ;
        RECT 2699.810 3313.340 2700.130 3313.400 ;
        RECT 2699.810 2552.960 2700.130 2553.020 ;
        RECT 2898.990 2552.960 2899.310 2553.020 ;
        RECT 2699.810 2552.820 2899.310 2552.960 ;
        RECT 2699.810 2552.760 2700.130 2552.820 ;
        RECT 2898.990 2552.760 2899.310 2552.820 ;
      LAYER via ;
        RECT 960.120 3313.340 960.380 3313.600 ;
        RECT 2699.840 3313.340 2700.100 3313.600 ;
        RECT 2699.840 2552.760 2700.100 2553.020 ;
        RECT 2899.020 2552.760 2899.280 2553.020 ;
      LAYER met2 ;
        RECT 960.120 3313.310 960.380 3313.630 ;
        RECT 2699.840 3313.310 2700.100 3313.630 ;
        RECT 960.180 3300.000 960.320 3313.310 ;
        RECT 960.120 3296.000 960.400 3300.000 ;
        RECT 2699.900 2553.050 2700.040 3313.310 ;
        RECT 2699.840 2552.730 2700.100 2553.050 ;
        RECT 2899.020 2552.730 2899.280 2553.050 ;
        RECT 2899.080 2551.885 2899.220 2552.730 ;
        RECT 2899.010 2551.515 2899.290 2551.885 ;
      LAYER via2 ;
        RECT 2899.010 2551.560 2899.290 2551.840 ;
      LAYER met3 ;
        RECT 2898.985 2551.850 2899.315 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2898.985 2551.550 2924.800 2551.850 ;
        RECT 2898.985 2551.535 2899.315 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1023.110 3313.880 1023.430 3313.940 ;
        RECT 2699.350 3313.880 2699.670 3313.940 ;
        RECT 1023.110 3313.740 2699.670 3313.880 ;
        RECT 1023.110 3313.680 1023.430 3313.740 ;
        RECT 2699.350 3313.680 2699.670 3313.740 ;
        RECT 2699.350 2787.560 2699.670 2787.620 ;
        RECT 2900.370 2787.560 2900.690 2787.620 ;
        RECT 2699.350 2787.420 2900.690 2787.560 ;
        RECT 2699.350 2787.360 2699.670 2787.420 ;
        RECT 2900.370 2787.360 2900.690 2787.420 ;
      LAYER via ;
        RECT 1023.140 3313.680 1023.400 3313.940 ;
        RECT 2699.380 3313.680 2699.640 3313.940 ;
        RECT 2699.380 2787.360 2699.640 2787.620 ;
        RECT 2900.400 2787.360 2900.660 2787.620 ;
      LAYER met2 ;
        RECT 1023.140 3313.650 1023.400 3313.970 ;
        RECT 2699.380 3313.650 2699.640 3313.970 ;
        RECT 1023.200 3300.000 1023.340 3313.650 ;
        RECT 1023.140 3296.000 1023.420 3300.000 ;
        RECT 2699.440 2787.650 2699.580 3313.650 ;
        RECT 2699.380 2787.330 2699.640 2787.650 ;
        RECT 2900.400 2787.330 2900.660 2787.650 ;
        RECT 2900.460 2786.485 2900.600 2787.330 ;
        RECT 2900.390 2786.115 2900.670 2786.485 ;
      LAYER via2 ;
        RECT 2900.390 2786.160 2900.670 2786.440 ;
      LAYER met3 ;
        RECT 2900.365 2786.450 2900.695 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.365 2786.150 2924.800 2786.450 ;
        RECT 2900.365 2786.135 2900.695 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1087.970 3296.880 1088.290 3296.940 ;
        RECT 2698.890 3296.880 2699.210 3296.940 ;
        RECT 1087.970 3296.740 2699.210 3296.880 ;
        RECT 1087.970 3296.680 1088.290 3296.740 ;
        RECT 2698.890 3296.680 2699.210 3296.740 ;
        RECT 2698.890 3022.160 2699.210 3022.220 ;
        RECT 2900.370 3022.160 2900.690 3022.220 ;
        RECT 2698.890 3022.020 2900.690 3022.160 ;
        RECT 2698.890 3021.960 2699.210 3022.020 ;
        RECT 2900.370 3021.960 2900.690 3022.020 ;
      LAYER via ;
        RECT 1088.000 3296.680 1088.260 3296.940 ;
        RECT 2698.920 3296.680 2699.180 3296.940 ;
        RECT 2698.920 3021.960 2699.180 3022.220 ;
        RECT 2900.400 3021.960 2900.660 3022.220 ;
      LAYER met2 ;
        RECT 1086.620 3297.050 1086.900 3300.000 ;
        RECT 1086.620 3296.970 1088.200 3297.050 ;
        RECT 1086.620 3296.910 1088.260 3296.970 ;
        RECT 1086.620 3296.000 1086.900 3296.910 ;
        RECT 1088.000 3296.650 1088.260 3296.910 ;
        RECT 2698.920 3296.650 2699.180 3296.970 ;
        RECT 2698.980 3022.250 2699.120 3296.650 ;
        RECT 2698.920 3021.930 2699.180 3022.250 ;
        RECT 2900.400 3021.930 2900.660 3022.250 ;
        RECT 2900.460 3021.085 2900.600 3021.930 ;
        RECT 2900.390 3020.715 2900.670 3021.085 ;
      LAYER via2 ;
        RECT 2900.390 3020.760 2900.670 3021.040 ;
      LAYER met3 ;
        RECT 2900.365 3021.050 2900.695 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.365 3020.750 2924.800 3021.050 ;
        RECT 2900.365 3020.735 2900.695 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1151.450 3297.560 1151.770 3297.620 ;
        RECT 2698.430 3297.560 2698.750 3297.620 ;
        RECT 1151.450 3297.420 2698.750 3297.560 ;
        RECT 1151.450 3297.360 1151.770 3297.420 ;
        RECT 2698.430 3297.360 2698.750 3297.420 ;
        RECT 2698.430 3256.760 2698.750 3256.820 ;
        RECT 2900.370 3256.760 2900.690 3256.820 ;
        RECT 2698.430 3256.620 2900.690 3256.760 ;
        RECT 2698.430 3256.560 2698.750 3256.620 ;
        RECT 2900.370 3256.560 2900.690 3256.620 ;
      LAYER via ;
        RECT 1151.480 3297.360 1151.740 3297.620 ;
        RECT 2698.460 3297.360 2698.720 3297.620 ;
        RECT 2698.460 3256.560 2698.720 3256.820 ;
        RECT 2900.400 3256.560 2900.660 3256.820 ;
      LAYER met2 ;
        RECT 1149.640 3297.730 1149.920 3300.000 ;
        RECT 1149.640 3297.650 1151.680 3297.730 ;
        RECT 1149.640 3297.590 1151.740 3297.650 ;
        RECT 1149.640 3296.000 1149.920 3297.590 ;
        RECT 1151.480 3297.330 1151.740 3297.590 ;
        RECT 2698.460 3297.330 2698.720 3297.650 ;
        RECT 2698.520 3256.850 2698.660 3297.330 ;
        RECT 2698.460 3256.530 2698.720 3256.850 ;
        RECT 2900.400 3256.530 2900.660 3256.850 ;
        RECT 2900.460 3255.685 2900.600 3256.530 ;
        RECT 2900.390 3255.315 2900.670 3255.685 ;
      LAYER via2 ;
        RECT 2900.390 3255.360 2900.670 3255.640 ;
      LAYER met3 ;
        RECT 2900.365 3255.650 2900.695 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.365 3255.350 2924.800 3255.650 ;
        RECT 2900.365 3255.335 2900.695 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1214.010 3484.900 1214.330 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 1214.010 3484.760 2901.150 3484.900 ;
        RECT 1214.010 3484.700 1214.330 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 1214.040 3484.700 1214.300 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 1214.040 3484.670 1214.300 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 1212.660 3299.770 1212.940 3300.000 ;
        RECT 1214.100 3299.770 1214.240 3484.670 ;
        RECT 1212.660 3299.630 1214.240 3299.770 ;
        RECT 1212.660 3296.000 1212.940 3299.630 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1276.110 3502.580 1276.430 3502.640 ;
        RECT 2635.870 3502.580 2636.190 3502.640 ;
        RECT 1276.110 3502.440 2636.190 3502.580 ;
        RECT 1276.110 3502.380 1276.430 3502.440 ;
        RECT 2635.870 3502.380 2636.190 3502.440 ;
      LAYER via ;
        RECT 1276.140 3502.380 1276.400 3502.640 ;
        RECT 2635.900 3502.380 2636.160 3502.640 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3502.670 2636.100 3517.600 ;
        RECT 1276.140 3502.350 1276.400 3502.670 ;
        RECT 2635.900 3502.350 2636.160 3502.670 ;
        RECT 1276.200 3300.000 1276.340 3502.350 ;
        RECT 1276.140 3296.000 1276.420 3300.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1345.110 3504.280 1345.430 3504.340 ;
        RECT 2311.570 3504.280 2311.890 3504.340 ;
        RECT 1345.110 3504.140 2311.890 3504.280 ;
        RECT 1345.110 3504.080 1345.430 3504.140 ;
        RECT 2311.570 3504.080 2311.890 3504.140 ;
      LAYER via ;
        RECT 1345.140 3504.080 1345.400 3504.340 ;
        RECT 2311.600 3504.080 2311.860 3504.340 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3504.370 2311.800 3517.600 ;
        RECT 1345.140 3504.050 1345.400 3504.370 ;
        RECT 2311.600 3504.050 2311.860 3504.370 ;
        RECT 1345.200 3300.450 1345.340 3504.050 ;
        RECT 1341.980 3300.310 1345.340 3300.450 ;
        RECT 1339.160 3299.090 1339.440 3300.000 ;
        RECT 1341.980 3299.090 1342.120 3300.310 ;
        RECT 1339.160 3298.950 1342.120 3299.090 ;
        RECT 1339.160 3296.000 1339.440 3298.950 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1407.210 3500.540 1407.530 3500.600 ;
        RECT 1987.270 3500.540 1987.590 3500.600 ;
        RECT 1407.210 3500.400 1987.590 3500.540 ;
        RECT 1407.210 3500.340 1407.530 3500.400 ;
        RECT 1987.270 3500.340 1987.590 3500.400 ;
      LAYER via ;
        RECT 1407.240 3500.340 1407.500 3500.600 ;
        RECT 1987.300 3500.340 1987.560 3500.600 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3500.630 1987.500 3517.600 ;
        RECT 1407.240 3500.310 1407.500 3500.630 ;
        RECT 1987.300 3500.310 1987.560 3500.630 ;
        RECT 1407.300 3300.450 1407.440 3500.310 ;
        RECT 1404.540 3300.310 1407.440 3300.450 ;
        RECT 1402.180 3299.090 1402.460 3300.000 ;
        RECT 1404.540 3299.090 1404.680 3300.310 ;
        RECT 1402.180 3298.950 1404.680 3299.090 ;
        RECT 1402.180 3296.000 1402.460 3298.950 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1469.310 3498.840 1469.630 3498.900 ;
        RECT 1662.510 3498.840 1662.830 3498.900 ;
        RECT 1469.310 3498.700 1662.830 3498.840 ;
        RECT 1469.310 3498.640 1469.630 3498.700 ;
        RECT 1662.510 3498.640 1662.830 3498.700 ;
      LAYER via ;
        RECT 1469.340 3498.640 1469.600 3498.900 ;
        RECT 1662.540 3498.640 1662.800 3498.900 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3498.930 1662.740 3517.600 ;
        RECT 1469.340 3498.610 1469.600 3498.930 ;
        RECT 1662.540 3498.610 1662.800 3498.930 ;
        RECT 1465.200 3299.090 1465.480 3300.000 ;
        RECT 1469.400 3299.090 1469.540 3498.610 ;
        RECT 1465.200 3298.950 1469.540 3299.090 ;
        RECT 1465.200 3296.000 1465.480 3298.950 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1489.625 3498.005 1489.795 3499.195 ;
      LAYER mcon ;
        RECT 1489.625 3499.025 1489.795 3499.195 ;
      LAYER met1 ;
        RECT 1338.210 3499.180 1338.530 3499.240 ;
        RECT 1489.565 3499.180 1489.855 3499.225 ;
        RECT 1338.210 3499.040 1489.855 3499.180 ;
        RECT 1338.210 3498.980 1338.530 3499.040 ;
        RECT 1489.565 3498.995 1489.855 3499.040 ;
        RECT 1489.565 3498.160 1489.855 3498.205 ;
        RECT 1524.970 3498.160 1525.290 3498.220 ;
        RECT 1489.565 3498.020 1525.290 3498.160 ;
        RECT 1489.565 3497.975 1489.855 3498.020 ;
        RECT 1524.970 3497.960 1525.290 3498.020 ;
      LAYER via ;
        RECT 1338.240 3498.980 1338.500 3499.240 ;
        RECT 1525.000 3497.960 1525.260 3498.220 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3499.270 1338.440 3517.600 ;
        RECT 1338.240 3498.950 1338.500 3499.270 ;
        RECT 1525.000 3497.930 1525.260 3498.250 ;
        RECT 1525.060 3300.450 1525.200 3497.930 ;
        RECT 1525.060 3300.310 1526.580 3300.450 ;
        RECT 1526.440 3299.090 1526.580 3300.310 ;
        RECT 1528.680 3299.090 1528.960 3300.000 ;
        RECT 1526.440 3298.950 1528.960 3299.090 ;
        RECT 1528.680 3296.000 1528.960 3298.950 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2694.750 441.560 2695.070 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 2694.750 441.420 2901.150 441.560 ;
        RECT 2694.750 441.360 2695.070 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 2694.780 441.360 2695.040 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 392.020 3297.050 392.300 3300.000 ;
        RECT 392.930 3297.050 393.210 3297.165 ;
        RECT 392.020 3296.910 393.210 3297.050 ;
        RECT 392.020 3296.000 392.300 3296.910 ;
        RECT 392.930 3296.795 393.210 3296.910 ;
        RECT 2694.770 3292.035 2695.050 3292.405 ;
        RECT 2694.840 441.650 2694.980 3292.035 ;
        RECT 2694.780 441.330 2695.040 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 392.930 3296.840 393.210 3297.120 ;
        RECT 2694.770 3292.080 2695.050 3292.360 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 392.905 3297.130 393.235 3297.145 ;
        RECT 405.990 3297.130 406.370 3297.140 ;
        RECT 392.905 3296.830 406.370 3297.130 ;
        RECT 392.905 3296.815 393.235 3296.830 ;
        RECT 405.990 3296.820 406.370 3296.830 ;
        RECT 405.990 3292.370 406.370 3292.380 ;
        RECT 2694.745 3292.370 2695.075 3292.385 ;
        RECT 405.990 3292.070 2695.075 3292.370 ;
        RECT 405.990 3292.060 406.370 3292.070 ;
        RECT 2694.745 3292.055 2695.075 3292.070 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
      LAYER via3 ;
        RECT 406.020 3296.820 406.340 3297.140 ;
        RECT 406.020 3292.060 406.340 3292.380 ;
      LAYER met4 ;
        RECT 406.015 3296.815 406.345 3297.145 ;
        RECT 406.030 3292.385 406.330 3296.815 ;
        RECT 406.015 3292.055 406.345 3292.385 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3500.200 1014.230 3500.260 ;
        RECT 1587.070 3500.200 1587.390 3500.260 ;
        RECT 1013.910 3500.060 1587.390 3500.200 ;
        RECT 1013.910 3500.000 1014.230 3500.060 ;
        RECT 1587.070 3500.000 1587.390 3500.060 ;
      LAYER via ;
        RECT 1013.940 3500.000 1014.200 3500.260 ;
        RECT 1587.100 3500.000 1587.360 3500.260 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3500.290 1014.140 3517.600 ;
        RECT 1013.940 3499.970 1014.200 3500.290 ;
        RECT 1587.100 3499.970 1587.360 3500.290 ;
        RECT 1587.160 3299.090 1587.300 3499.970 ;
        RECT 1591.700 3299.090 1591.980 3300.000 ;
        RECT 1587.160 3298.950 1591.980 3299.090 ;
        RECT 1591.700 3296.000 1591.980 3298.950 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3504.620 689.470 3504.680 ;
        RECT 1649.170 3504.620 1649.490 3504.680 ;
        RECT 689.150 3504.480 1649.490 3504.620 ;
        RECT 689.150 3504.420 689.470 3504.480 ;
        RECT 1649.170 3504.420 1649.490 3504.480 ;
      LAYER via ;
        RECT 689.180 3504.420 689.440 3504.680 ;
        RECT 1649.200 3504.420 1649.460 3504.680 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3504.710 689.380 3517.600 ;
        RECT 689.180 3504.390 689.440 3504.710 ;
        RECT 1649.200 3504.390 1649.460 3504.710 ;
        RECT 1649.260 3300.450 1649.400 3504.390 ;
        RECT 1649.260 3300.310 1652.620 3300.450 ;
        RECT 1652.480 3299.090 1652.620 3300.310 ;
        RECT 1654.720 3299.090 1655.000 3300.000 ;
        RECT 1652.480 3298.950 1655.000 3299.090 ;
        RECT 1654.720 3296.000 1655.000 3298.950 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 3502.920 365.170 3502.980 ;
        RECT 1718.170 3502.920 1718.490 3502.980 ;
        RECT 364.850 3502.780 1718.490 3502.920 ;
        RECT 364.850 3502.720 365.170 3502.780 ;
        RECT 1718.170 3502.720 1718.490 3502.780 ;
      LAYER via ;
        RECT 364.880 3502.720 365.140 3502.980 ;
        RECT 1718.200 3502.720 1718.460 3502.980 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3503.010 365.080 3517.600 ;
        RECT 364.880 3502.690 365.140 3503.010 ;
        RECT 1718.200 3502.690 1718.460 3503.010 ;
        RECT 1718.260 3300.000 1718.400 3502.690 ;
        RECT 1718.200 3296.000 1718.480 3300.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.845 40.780 3517.600 ;
        RECT 40.570 3501.475 40.850 3501.845 ;
        RECT 1780.290 3501.475 1780.570 3501.845 ;
        RECT 1780.360 3299.770 1780.500 3501.475 ;
        RECT 1781.220 3299.770 1781.500 3300.000 ;
        RECT 1780.360 3299.630 1781.500 3299.770 ;
        RECT 1781.220 3296.000 1781.500 3299.630 ;
      LAYER via2 ;
        RECT 40.570 3501.520 40.850 3501.800 ;
        RECT 1780.290 3501.520 1780.570 3501.800 ;
      LAYER met3 ;
        RECT 40.545 3501.810 40.875 3501.825 ;
        RECT 1780.265 3501.810 1780.595 3501.825 ;
        RECT 40.545 3501.510 1780.595 3501.810 ;
        RECT 40.545 3501.495 40.875 3501.510 ;
        RECT 1780.265 3501.495 1780.595 3501.510 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1842.905 3295.705 1843.075 3298.255 ;
      LAYER mcon ;
        RECT 1842.905 3298.085 1843.075 3298.255 ;
      LAYER met1 ;
        RECT 1842.830 3298.240 1843.150 3298.300 ;
        RECT 1842.635 3298.100 1843.150 3298.240 ;
        RECT 1842.830 3298.040 1843.150 3298.100 ;
        RECT 43.310 3295.860 43.630 3295.920 ;
        RECT 1842.845 3295.860 1843.135 3295.905 ;
        RECT 43.310 3295.720 1843.135 3295.860 ;
        RECT 43.310 3295.660 43.630 3295.720 ;
        RECT 1842.845 3295.675 1843.135 3295.720 ;
        RECT 15.710 3267.980 16.030 3268.040 ;
        RECT 43.310 3267.980 43.630 3268.040 ;
        RECT 15.710 3267.840 43.630 3267.980 ;
        RECT 15.710 3267.780 16.030 3267.840 ;
        RECT 43.310 3267.780 43.630 3267.840 ;
      LAYER via ;
        RECT 1842.860 3298.040 1843.120 3298.300 ;
        RECT 43.340 3295.660 43.600 3295.920 ;
        RECT 15.740 3267.780 16.000 3268.040 ;
        RECT 43.340 3267.780 43.600 3268.040 ;
      LAYER met2 ;
        RECT 1844.240 3298.410 1844.520 3300.000 ;
        RECT 1842.920 3298.330 1844.520 3298.410 ;
        RECT 1842.860 3298.270 1844.520 3298.330 ;
        RECT 1842.860 3298.010 1843.120 3298.270 ;
        RECT 1844.240 3296.000 1844.520 3298.270 ;
        RECT 43.340 3295.630 43.600 3295.950 ;
        RECT 43.400 3268.070 43.540 3295.630 ;
        RECT 15.740 3267.925 16.000 3268.070 ;
        RECT 15.730 3267.555 16.010 3267.925 ;
        RECT 43.340 3267.750 43.600 3268.070 ;
      LAYER via2 ;
        RECT 15.730 3267.600 16.010 3267.880 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.705 3267.890 16.035 3267.905 ;
        RECT -4.800 3267.590 16.035 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.705 3267.575 16.035 3267.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1906.385 3295.365 1906.555 3298.255 ;
      LAYER mcon ;
        RECT 1906.385 3298.085 1906.555 3298.255 ;
      LAYER met1 ;
        RECT 1906.310 3298.240 1906.630 3298.300 ;
        RECT 1906.115 3298.100 1906.630 3298.240 ;
        RECT 1906.310 3298.040 1906.630 3298.100 ;
        RECT 43.770 3295.520 44.090 3295.580 ;
        RECT 1906.325 3295.520 1906.615 3295.565 ;
        RECT 43.770 3295.380 1906.615 3295.520 ;
        RECT 43.770 3295.320 44.090 3295.380 ;
        RECT 1906.325 3295.335 1906.615 3295.380 ;
        RECT 15.710 2980.340 16.030 2980.400 ;
        RECT 43.770 2980.340 44.090 2980.400 ;
        RECT 15.710 2980.200 44.090 2980.340 ;
        RECT 15.710 2980.140 16.030 2980.200 ;
        RECT 43.770 2980.140 44.090 2980.200 ;
      LAYER via ;
        RECT 1906.340 3298.040 1906.600 3298.300 ;
        RECT 43.800 3295.320 44.060 3295.580 ;
        RECT 15.740 2980.140 16.000 2980.400 ;
        RECT 43.800 2980.140 44.060 2980.400 ;
      LAYER met2 ;
        RECT 1907.720 3298.410 1908.000 3300.000 ;
        RECT 1906.400 3298.330 1908.000 3298.410 ;
        RECT 1906.340 3298.270 1908.000 3298.330 ;
        RECT 1906.340 3298.010 1906.600 3298.270 ;
        RECT 1907.720 3296.000 1908.000 3298.270 ;
        RECT 43.800 3295.290 44.060 3295.610 ;
        RECT 43.860 2980.430 44.000 3295.290 ;
        RECT 15.740 2980.285 16.000 2980.430 ;
        RECT 15.730 2979.915 16.010 2980.285 ;
        RECT 43.800 2980.110 44.060 2980.430 ;
      LAYER via2 ;
        RECT 15.730 2979.960 16.010 2980.240 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 15.705 2980.250 16.035 2980.265 ;
        RECT -4.800 2979.950 16.035 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 15.705 2979.935 16.035 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 44.230 3313.200 44.550 3313.260 ;
        RECT 1970.710 3313.200 1971.030 3313.260 ;
        RECT 44.230 3313.060 1971.030 3313.200 ;
        RECT 44.230 3313.000 44.550 3313.060 ;
        RECT 1970.710 3313.000 1971.030 3313.060 ;
        RECT 16.170 2694.060 16.490 2694.120 ;
        RECT 44.230 2694.060 44.550 2694.120 ;
        RECT 16.170 2693.920 44.550 2694.060 ;
        RECT 16.170 2693.860 16.490 2693.920 ;
        RECT 44.230 2693.860 44.550 2693.920 ;
      LAYER via ;
        RECT 44.260 3313.000 44.520 3313.260 ;
        RECT 1970.740 3313.000 1971.000 3313.260 ;
        RECT 16.200 2693.860 16.460 2694.120 ;
        RECT 44.260 2693.860 44.520 2694.120 ;
      LAYER met2 ;
        RECT 44.260 3312.970 44.520 3313.290 ;
        RECT 1970.740 3312.970 1971.000 3313.290 ;
        RECT 44.320 2694.150 44.460 3312.970 ;
        RECT 1970.800 3300.000 1970.940 3312.970 ;
        RECT 1970.740 3296.000 1971.020 3300.000 ;
        RECT 16.200 2693.830 16.460 2694.150 ;
        RECT 44.260 2693.830 44.520 2694.150 ;
        RECT 16.260 2693.325 16.400 2693.830 ;
        RECT 16.190 2692.955 16.470 2693.325 ;
      LAYER via2 ;
        RECT 16.190 2693.000 16.470 2693.280 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 16.165 2693.290 16.495 2693.305 ;
        RECT -4.800 2692.990 16.495 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 16.165 2692.975 16.495 2692.990 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 47.910 3312.860 48.230 3312.920 ;
        RECT 2033.730 3312.860 2034.050 3312.920 ;
        RECT 47.910 3312.720 2034.050 3312.860 ;
        RECT 47.910 3312.660 48.230 3312.720 ;
        RECT 2033.730 3312.660 2034.050 3312.720 ;
        RECT 16.170 2406.080 16.490 2406.140 ;
        RECT 47.910 2406.080 48.230 2406.140 ;
        RECT 16.170 2405.940 48.230 2406.080 ;
        RECT 16.170 2405.880 16.490 2405.940 ;
        RECT 47.910 2405.880 48.230 2405.940 ;
      LAYER via ;
        RECT 47.940 3312.660 48.200 3312.920 ;
        RECT 2033.760 3312.660 2034.020 3312.920 ;
        RECT 16.200 2405.880 16.460 2406.140 ;
        RECT 47.940 2405.880 48.200 2406.140 ;
      LAYER met2 ;
        RECT 47.940 3312.630 48.200 3312.950 ;
        RECT 2033.760 3312.630 2034.020 3312.950 ;
        RECT 48.000 2406.170 48.140 3312.630 ;
        RECT 2033.820 3300.000 2033.960 3312.630 ;
        RECT 2033.760 3296.000 2034.040 3300.000 ;
        RECT 16.200 2405.850 16.460 2406.170 ;
        RECT 47.940 2405.850 48.200 2406.170 ;
        RECT 16.260 2405.685 16.400 2405.850 ;
        RECT 16.190 2405.315 16.470 2405.685 ;
      LAYER via2 ;
        RECT 16.190 2405.360 16.470 2405.640 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 16.165 2405.650 16.495 2405.665 ;
        RECT -4.800 2405.350 16.495 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 16.165 2405.335 16.495 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1153.290 3311.160 1153.610 3311.220 ;
        RECT 2096.750 3311.160 2097.070 3311.220 ;
        RECT 1153.290 3311.020 2097.070 3311.160 ;
        RECT 1153.290 3310.960 1153.610 3311.020 ;
        RECT 2096.750 3310.960 2097.070 3311.020 ;
        RECT 16.630 3298.240 16.950 3298.300 ;
        RECT 1153.290 3298.240 1153.610 3298.300 ;
        RECT 16.630 3298.100 1153.610 3298.240 ;
        RECT 16.630 3298.040 16.950 3298.100 ;
        RECT 1153.290 3298.040 1153.610 3298.100 ;
      LAYER via ;
        RECT 1153.320 3310.960 1153.580 3311.220 ;
        RECT 2096.780 3310.960 2097.040 3311.220 ;
        RECT 16.660 3298.040 16.920 3298.300 ;
        RECT 1153.320 3298.040 1153.580 3298.300 ;
      LAYER met2 ;
        RECT 1153.320 3310.930 1153.580 3311.250 ;
        RECT 2096.780 3310.930 2097.040 3311.250 ;
        RECT 1153.380 3298.330 1153.520 3310.930 ;
        RECT 2096.840 3300.000 2096.980 3310.930 ;
        RECT 16.660 3298.010 16.920 3298.330 ;
        RECT 1153.320 3298.010 1153.580 3298.330 ;
        RECT 16.720 2118.725 16.860 3298.010 ;
        RECT 2096.780 3296.000 2097.060 3300.000 ;
        RECT 16.650 2118.355 16.930 2118.725 ;
      LAYER via2 ;
        RECT 16.650 2118.400 16.930 2118.680 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.625 2118.690 16.955 2118.705 ;
        RECT -4.800 2118.390 16.955 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.625 2118.375 16.955 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 47.450 3312.180 47.770 3312.240 ;
        RECT 2160.230 3312.180 2160.550 3312.240 ;
        RECT 47.450 3312.040 2160.550 3312.180 ;
        RECT 47.450 3311.980 47.770 3312.040 ;
        RECT 2160.230 3311.980 2160.550 3312.040 ;
        RECT 15.710 1833.520 16.030 1833.580 ;
        RECT 47.450 1833.520 47.770 1833.580 ;
        RECT 15.710 1833.380 47.770 1833.520 ;
        RECT 15.710 1833.320 16.030 1833.380 ;
        RECT 47.450 1833.320 47.770 1833.380 ;
      LAYER via ;
        RECT 47.480 3311.980 47.740 3312.240 ;
        RECT 2160.260 3311.980 2160.520 3312.240 ;
        RECT 15.740 1833.320 16.000 1833.580 ;
        RECT 47.480 1833.320 47.740 1833.580 ;
      LAYER met2 ;
        RECT 47.480 3311.950 47.740 3312.270 ;
        RECT 2160.260 3311.950 2160.520 3312.270 ;
        RECT 47.540 1833.610 47.680 3311.950 ;
        RECT 2160.320 3300.000 2160.460 3311.950 ;
        RECT 2160.260 3296.000 2160.540 3300.000 ;
        RECT 15.740 1833.290 16.000 1833.610 ;
        RECT 47.480 1833.290 47.740 1833.610 ;
        RECT 15.800 1831.085 15.940 1833.290 ;
        RECT 15.730 1830.715 16.010 1831.085 ;
      LAYER via2 ;
        RECT 15.730 1830.760 16.010 1831.040 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 15.705 1831.050 16.035 1831.065 ;
        RECT -4.800 1830.750 16.035 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 15.705 1830.735 16.035 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 455.010 3309.460 455.330 3309.520 ;
        RECT 829.450 3309.460 829.770 3309.520 ;
        RECT 455.010 3309.320 829.770 3309.460 ;
        RECT 455.010 3309.260 455.330 3309.320 ;
        RECT 829.450 3309.260 829.770 3309.320 ;
        RECT 829.450 3296.540 829.770 3296.600 ;
        RECT 2903.130 3296.540 2903.450 3296.600 ;
        RECT 829.450 3296.400 2903.450 3296.540 ;
        RECT 829.450 3296.340 829.770 3296.400 ;
        RECT 2903.130 3296.340 2903.450 3296.400 ;
      LAYER via ;
        RECT 455.040 3309.260 455.300 3309.520 ;
        RECT 829.480 3309.260 829.740 3309.520 ;
        RECT 829.480 3296.340 829.740 3296.600 ;
        RECT 2903.160 3296.340 2903.420 3296.600 ;
      LAYER met2 ;
        RECT 455.040 3309.230 455.300 3309.550 ;
        RECT 829.480 3309.230 829.740 3309.550 ;
        RECT 455.100 3300.000 455.240 3309.230 ;
        RECT 455.040 3296.000 455.320 3300.000 ;
        RECT 829.540 3296.630 829.680 3309.230 ;
        RECT 829.480 3296.310 829.740 3296.630 ;
        RECT 2903.160 3296.310 2903.420 3296.630 ;
        RECT 2903.220 674.405 2903.360 3296.310 ;
        RECT 2903.150 674.035 2903.430 674.405 ;
      LAYER via2 ;
        RECT 2903.150 674.080 2903.430 674.360 ;
      LAYER met3 ;
        RECT 2903.125 674.370 2903.455 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2903.125 674.070 2924.800 674.370 ;
        RECT 2903.125 674.055 2903.455 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 265.490 3307.760 265.810 3307.820 ;
        RECT 2223.250 3307.760 2223.570 3307.820 ;
        RECT 265.490 3307.620 2223.570 3307.760 ;
        RECT 265.490 3307.560 265.810 3307.620 ;
        RECT 2223.250 3307.560 2223.570 3307.620 ;
        RECT 15.250 1545.540 15.570 1545.600 ;
        RECT 265.490 1545.540 265.810 1545.600 ;
        RECT 15.250 1545.400 265.810 1545.540 ;
        RECT 15.250 1545.340 15.570 1545.400 ;
        RECT 265.490 1545.340 265.810 1545.400 ;
      LAYER via ;
        RECT 265.520 3307.560 265.780 3307.820 ;
        RECT 2223.280 3307.560 2223.540 3307.820 ;
        RECT 15.280 1545.340 15.540 1545.600 ;
        RECT 265.520 1545.340 265.780 1545.600 ;
      LAYER met2 ;
        RECT 265.520 3307.530 265.780 3307.850 ;
        RECT 2223.280 3307.530 2223.540 3307.850 ;
        RECT 265.580 1545.630 265.720 3307.530 ;
        RECT 2223.340 3300.000 2223.480 3307.530 ;
        RECT 2223.280 3296.000 2223.560 3300.000 ;
        RECT 15.280 1545.310 15.540 1545.630 ;
        RECT 265.520 1545.310 265.780 1545.630 ;
        RECT 15.340 1544.125 15.480 1545.310 ;
        RECT 15.270 1543.755 15.550 1544.125 ;
      LAYER via2 ;
        RECT 15.270 1543.800 15.550 1544.080 ;
      LAYER met3 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 15.245 1544.090 15.575 1544.105 ;
        RECT -4.800 1543.790 15.575 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 15.245 1543.775 15.575 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 272.390 3306.740 272.710 3306.800 ;
        RECT 2286.270 3306.740 2286.590 3306.800 ;
        RECT 272.390 3306.600 2286.590 3306.740 ;
        RECT 272.390 3306.540 272.710 3306.600 ;
        RECT 2286.270 3306.540 2286.590 3306.600 ;
        RECT 16.630 1331.680 16.950 1331.740 ;
        RECT 272.390 1331.680 272.710 1331.740 ;
        RECT 16.630 1331.540 272.710 1331.680 ;
        RECT 16.630 1331.480 16.950 1331.540 ;
        RECT 272.390 1331.480 272.710 1331.540 ;
      LAYER via ;
        RECT 272.420 3306.540 272.680 3306.800 ;
        RECT 2286.300 3306.540 2286.560 3306.800 ;
        RECT 16.660 1331.480 16.920 1331.740 ;
        RECT 272.420 1331.480 272.680 1331.740 ;
      LAYER met2 ;
        RECT 272.420 3306.510 272.680 3306.830 ;
        RECT 2286.300 3306.510 2286.560 3306.830 ;
        RECT 272.480 1331.770 272.620 3306.510 ;
        RECT 2286.360 3300.000 2286.500 3306.510 ;
        RECT 2286.300 3296.000 2286.580 3300.000 ;
        RECT 16.660 1331.450 16.920 1331.770 ;
        RECT 272.420 1331.450 272.680 1331.770 ;
        RECT 16.720 1328.565 16.860 1331.450 ;
        RECT 16.650 1328.195 16.930 1328.565 ;
      LAYER via2 ;
        RECT 16.650 1328.240 16.930 1328.520 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 16.625 1328.530 16.955 1328.545 ;
        RECT -4.800 1328.230 16.955 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 16.625 1328.215 16.955 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2347.985 3292.645 2348.155 3298.255 ;
      LAYER mcon ;
        RECT 2347.985 3298.085 2348.155 3298.255 ;
      LAYER met1 ;
        RECT 2347.910 3298.240 2348.230 3298.300 ;
        RECT 2347.715 3298.100 2348.230 3298.240 ;
        RECT 2347.910 3298.040 2348.230 3298.100 ;
        RECT 46.530 3292.800 46.850 3292.860 ;
        RECT 2347.925 3292.800 2348.215 3292.845 ;
        RECT 46.530 3292.660 2348.215 3292.800 ;
        RECT 46.530 3292.600 46.850 3292.660 ;
        RECT 2347.925 3292.615 2348.215 3292.660 ;
        RECT 16.630 1115.440 16.950 1115.500 ;
        RECT 46.530 1115.440 46.850 1115.500 ;
        RECT 16.630 1115.300 46.850 1115.440 ;
        RECT 16.630 1115.240 16.950 1115.300 ;
        RECT 46.530 1115.240 46.850 1115.300 ;
      LAYER via ;
        RECT 2347.940 3298.040 2348.200 3298.300 ;
        RECT 46.560 3292.600 46.820 3292.860 ;
        RECT 16.660 1115.240 16.920 1115.500 ;
        RECT 46.560 1115.240 46.820 1115.500 ;
      LAYER met2 ;
        RECT 2349.780 3298.410 2350.060 3300.000 ;
        RECT 2348.000 3298.330 2350.060 3298.410 ;
        RECT 2347.940 3298.270 2350.060 3298.330 ;
        RECT 2347.940 3298.010 2348.200 3298.270 ;
        RECT 2349.780 3296.000 2350.060 3298.270 ;
        RECT 46.560 3292.570 46.820 3292.890 ;
        RECT 46.620 1115.530 46.760 3292.570 ;
        RECT 16.660 1115.210 16.920 1115.530 ;
        RECT 46.560 1115.210 46.820 1115.530 ;
        RECT 16.720 1113.005 16.860 1115.210 ;
        RECT 16.650 1112.635 16.930 1113.005 ;
      LAYER via2 ;
        RECT 16.650 1112.680 16.930 1112.960 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 16.625 1112.970 16.955 1112.985 ;
        RECT -4.800 1112.670 16.955 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 16.625 1112.655 16.955 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 898.180 16.950 898.240 ;
        RECT 45.150 898.180 45.470 898.240 ;
        RECT 16.630 898.040 45.470 898.180 ;
        RECT 16.630 897.980 16.950 898.040 ;
        RECT 45.150 897.980 45.470 898.040 ;
      LAYER via ;
        RECT 16.660 897.980 16.920 898.240 ;
        RECT 45.180 897.980 45.440 898.240 ;
      LAYER met2 ;
        RECT 45.170 3309.715 45.450 3310.085 ;
        RECT 2412.790 3309.715 2413.070 3310.085 ;
        RECT 45.240 898.270 45.380 3309.715 ;
        RECT 2412.860 3300.000 2413.000 3309.715 ;
        RECT 2412.800 3296.000 2413.080 3300.000 ;
        RECT 16.660 897.950 16.920 898.270 ;
        RECT 45.180 897.950 45.440 898.270 ;
        RECT 16.720 897.445 16.860 897.950 ;
        RECT 16.650 897.075 16.930 897.445 ;
      LAYER via2 ;
        RECT 45.170 3309.760 45.450 3310.040 ;
        RECT 2412.790 3309.760 2413.070 3310.040 ;
        RECT 16.650 897.120 16.930 897.400 ;
      LAYER met3 ;
        RECT 45.145 3310.050 45.475 3310.065 ;
        RECT 2412.765 3310.050 2413.095 3310.065 ;
        RECT 45.145 3309.750 2413.095 3310.050 ;
        RECT 45.145 3309.735 45.475 3309.750 ;
        RECT 2412.765 3309.735 2413.095 3309.750 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.625 897.410 16.955 897.425 ;
        RECT -4.800 897.110 16.955 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 16.625 897.095 16.955 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2287.650 3306.740 2287.970 3306.800 ;
        RECT 2475.790 3306.740 2476.110 3306.800 ;
        RECT 2287.650 3306.600 2476.110 3306.740 ;
        RECT 2287.650 3306.540 2287.970 3306.600 ;
        RECT 2475.790 3306.540 2476.110 3306.600 ;
      LAYER via ;
        RECT 2287.680 3306.540 2287.940 3306.800 ;
        RECT 2475.820 3306.540 2476.080 3306.800 ;
      LAYER met2 ;
        RECT 2287.680 3306.510 2287.940 3306.830 ;
        RECT 2475.820 3306.510 2476.080 3306.830 ;
        RECT 2287.740 3297.165 2287.880 3306.510 ;
        RECT 2475.880 3300.000 2476.020 3306.510 ;
        RECT 2287.670 3296.795 2287.950 3297.165 ;
        RECT 2475.820 3296.000 2476.100 3300.000 ;
        RECT 18.490 3294.075 18.770 3294.445 ;
        RECT 18.560 681.885 18.700 3294.075 ;
        RECT 18.490 681.515 18.770 681.885 ;
      LAYER via2 ;
        RECT 2287.670 3296.840 2287.950 3297.120 ;
        RECT 18.490 3294.120 18.770 3294.400 ;
        RECT 18.490 681.560 18.770 681.840 ;
      LAYER met3 ;
        RECT 2280.030 3297.130 2280.410 3297.140 ;
        RECT 2287.645 3297.130 2287.975 3297.145 ;
        RECT 2280.030 3296.830 2287.975 3297.130 ;
        RECT 2280.030 3296.820 2280.410 3296.830 ;
        RECT 2287.645 3296.815 2287.975 3296.830 ;
        RECT 18.465 3294.410 18.795 3294.425 ;
        RECT 2280.030 3294.410 2280.410 3294.420 ;
        RECT 18.465 3294.110 2280.410 3294.410 ;
        RECT 18.465 3294.095 18.795 3294.110 ;
        RECT 2280.030 3294.100 2280.410 3294.110 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 18.465 681.850 18.795 681.865 ;
        RECT -4.800 681.550 18.795 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 18.465 681.535 18.795 681.550 ;
      LAYER via3 ;
        RECT 2280.060 3296.820 2280.380 3297.140 ;
        RECT 2280.060 3294.100 2280.380 3294.420 ;
      LAYER met4 ;
        RECT 2280.055 3296.815 2280.385 3297.145 ;
        RECT 2280.070 3294.425 2280.370 3296.815 ;
        RECT 2280.055 3294.095 2280.385 3294.425 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 469.100 16.950 469.160 ;
        RECT 293.090 469.100 293.410 469.160 ;
        RECT 16.630 468.960 293.410 469.100 ;
        RECT 16.630 468.900 16.950 468.960 ;
        RECT 293.090 468.900 293.410 468.960 ;
      LAYER via ;
        RECT 16.660 468.900 16.920 469.160 ;
        RECT 293.120 468.900 293.380 469.160 ;
      LAYER met2 ;
        RECT 293.110 3310.395 293.390 3310.765 ;
        RECT 2538.830 3310.395 2539.110 3310.765 ;
        RECT 293.180 469.190 293.320 3310.395 ;
        RECT 2538.900 3300.000 2539.040 3310.395 ;
        RECT 2538.840 3296.000 2539.120 3300.000 ;
        RECT 16.660 468.870 16.920 469.190 ;
        RECT 293.120 468.870 293.380 469.190 ;
        RECT 16.720 466.325 16.860 468.870 ;
        RECT 16.650 465.955 16.930 466.325 ;
      LAYER via2 ;
        RECT 293.110 3310.440 293.390 3310.720 ;
        RECT 2538.830 3310.440 2539.110 3310.720 ;
        RECT 16.650 466.000 16.930 466.280 ;
      LAYER met3 ;
        RECT 293.085 3310.730 293.415 3310.745 ;
        RECT 2538.805 3310.730 2539.135 3310.745 ;
        RECT 293.085 3310.430 2539.135 3310.730 ;
        RECT 293.085 3310.415 293.415 3310.430 ;
        RECT 2538.805 3310.415 2539.135 3310.430 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 16.625 466.290 16.955 466.305 ;
        RECT -4.800 465.990 16.955 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 16.625 465.975 16.955 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.030 3306.315 18.310 3306.685 ;
        RECT 2602.310 3306.315 2602.590 3306.685 ;
        RECT 18.100 250.765 18.240 3306.315 ;
        RECT 2602.380 3300.000 2602.520 3306.315 ;
        RECT 2602.320 3296.000 2602.600 3300.000 ;
        RECT 18.030 250.395 18.310 250.765 ;
      LAYER via2 ;
        RECT 18.030 3306.360 18.310 3306.640 ;
        RECT 2602.310 3306.360 2602.590 3306.640 ;
        RECT 18.030 250.440 18.310 250.720 ;
      LAYER met3 ;
        RECT 18.005 3306.650 18.335 3306.665 ;
        RECT 2602.285 3306.650 2602.615 3306.665 ;
        RECT 18.005 3306.350 2602.615 3306.650 ;
        RECT 18.005 3306.335 18.335 3306.350 ;
        RECT 2602.285 3306.335 2602.615 3306.350 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 18.005 250.730 18.335 250.745 ;
        RECT -4.800 250.430 18.335 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 18.005 250.415 18.335 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.110 3304.955 17.390 3305.325 ;
        RECT 2665.330 3304.955 2665.610 3305.325 ;
        RECT 17.180 35.885 17.320 3304.955 ;
        RECT 2665.400 3300.000 2665.540 3304.955 ;
        RECT 2665.340 3296.000 2665.620 3300.000 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 17.110 3305.000 17.390 3305.280 ;
        RECT 2665.330 3305.000 2665.610 3305.280 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 17.085 3305.290 17.415 3305.305 ;
        RECT 2665.305 3305.290 2665.635 3305.305 ;
        RECT 17.085 3304.990 2665.635 3305.290 ;
        RECT 17.085 3304.975 17.415 3304.990 ;
        RECT 2665.305 3304.975 2665.635 3304.990 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 518.030 3306.060 518.350 3306.120 ;
        RECT 2701.190 3306.060 2701.510 3306.120 ;
        RECT 518.030 3305.920 2701.510 3306.060 ;
        RECT 518.030 3305.860 518.350 3305.920 ;
        RECT 2701.190 3305.860 2701.510 3305.920 ;
        RECT 2701.190 910.760 2701.510 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 2701.190 910.620 2901.150 910.760 ;
        RECT 2701.190 910.560 2701.510 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 518.060 3305.860 518.320 3306.120 ;
        RECT 2701.220 3305.860 2701.480 3306.120 ;
        RECT 2701.220 910.560 2701.480 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 518.060 3305.830 518.320 3306.150 ;
        RECT 2701.220 3305.830 2701.480 3306.150 ;
        RECT 518.120 3300.000 518.260 3305.830 ;
        RECT 518.060 3296.000 518.340 3300.000 ;
        RECT 2701.280 910.850 2701.420 3305.830 ;
        RECT 2701.220 910.530 2701.480 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 582.965 3292.985 583.135 3296.555 ;
      LAYER mcon ;
        RECT 582.965 3296.385 583.135 3296.555 ;
      LAYER met1 ;
        RECT 582.890 3296.540 583.210 3296.600 ;
        RECT 582.695 3296.400 583.210 3296.540 ;
        RECT 582.890 3296.340 583.210 3296.400 ;
        RECT 582.905 3293.140 583.195 3293.185 ;
        RECT 2701.650 3293.140 2701.970 3293.200 ;
        RECT 582.905 3293.000 2701.970 3293.140 ;
        RECT 582.905 3292.955 583.195 3293.000 ;
        RECT 2701.650 3292.940 2701.970 3293.000 ;
        RECT 2701.650 1145.360 2701.970 1145.420 ;
        RECT 2898.990 1145.360 2899.310 1145.420 ;
        RECT 2701.650 1145.220 2899.310 1145.360 ;
        RECT 2701.650 1145.160 2701.970 1145.220 ;
        RECT 2898.990 1145.160 2899.310 1145.220 ;
      LAYER via ;
        RECT 582.920 3296.340 583.180 3296.600 ;
        RECT 2701.680 3292.940 2701.940 3293.200 ;
        RECT 2701.680 1145.160 2701.940 1145.420 ;
        RECT 2899.020 1145.160 2899.280 1145.420 ;
      LAYER met2 ;
        RECT 581.080 3296.370 581.360 3300.000 ;
        RECT 582.920 3296.370 583.180 3296.630 ;
        RECT 581.080 3296.310 583.180 3296.370 ;
        RECT 581.080 3296.230 583.120 3296.310 ;
        RECT 581.080 3296.000 581.360 3296.230 ;
        RECT 2701.680 3292.910 2701.940 3293.230 ;
        RECT 2701.740 1145.450 2701.880 3292.910 ;
        RECT 2701.680 1145.130 2701.940 1145.450 ;
        RECT 2899.020 1145.130 2899.280 1145.450 ;
        RECT 2899.080 1144.285 2899.220 1145.130 ;
        RECT 2899.010 1143.915 2899.290 1144.285 ;
      LAYER via2 ;
        RECT 2899.010 1143.960 2899.290 1144.240 ;
      LAYER met3 ;
        RECT 2898.985 1144.250 2899.315 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2898.985 1143.950 2924.800 1144.250 ;
        RECT 2898.985 1143.935 2899.315 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 646.445 3294.005 646.615 3296.555 ;
      LAYER mcon ;
        RECT 646.445 3296.385 646.615 3296.555 ;
      LAYER met1 ;
        RECT 646.370 3296.540 646.690 3296.600 ;
        RECT 646.175 3296.400 646.690 3296.540 ;
        RECT 646.370 3296.340 646.690 3296.400 ;
        RECT 646.385 3294.160 646.675 3294.205 ;
        RECT 2702.570 3294.160 2702.890 3294.220 ;
        RECT 646.385 3294.020 2702.890 3294.160 ;
        RECT 646.385 3293.975 646.675 3294.020 ;
        RECT 2702.570 3293.960 2702.890 3294.020 ;
        RECT 2702.570 1379.960 2702.890 1380.020 ;
        RECT 2898.990 1379.960 2899.310 1380.020 ;
        RECT 2702.570 1379.820 2899.310 1379.960 ;
        RECT 2702.570 1379.760 2702.890 1379.820 ;
        RECT 2898.990 1379.760 2899.310 1379.820 ;
      LAYER via ;
        RECT 646.400 3296.340 646.660 3296.600 ;
        RECT 2702.600 3293.960 2702.860 3294.220 ;
        RECT 2702.600 1379.760 2702.860 1380.020 ;
        RECT 2899.020 1379.760 2899.280 1380.020 ;
      LAYER met2 ;
        RECT 644.560 3296.370 644.840 3300.000 ;
        RECT 646.400 3296.370 646.660 3296.630 ;
        RECT 644.560 3296.310 646.660 3296.370 ;
        RECT 644.560 3296.230 646.600 3296.310 ;
        RECT 644.560 3296.000 644.840 3296.230 ;
        RECT 2702.600 3293.930 2702.860 3294.250 ;
        RECT 2702.660 1380.050 2702.800 3293.930 ;
        RECT 2702.600 1379.730 2702.860 1380.050 ;
        RECT 2899.020 1379.730 2899.280 1380.050 ;
        RECT 2899.080 1378.885 2899.220 1379.730 ;
        RECT 2899.010 1378.515 2899.290 1378.885 ;
      LAYER via2 ;
        RECT 2899.010 1378.560 2899.290 1378.840 ;
      LAYER met3 ;
        RECT 2898.985 1378.850 2899.315 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2898.985 1378.550 2924.800 1378.850 ;
        RECT 2898.985 1378.535 2899.315 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 707.550 3307.080 707.870 3307.140 ;
        RECT 2703.490 3307.080 2703.810 3307.140 ;
        RECT 707.550 3306.940 2703.810 3307.080 ;
        RECT 707.550 3306.880 707.870 3306.940 ;
        RECT 2703.490 3306.880 2703.810 3306.940 ;
        RECT 2703.490 1614.560 2703.810 1614.620 ;
        RECT 2898.990 1614.560 2899.310 1614.620 ;
        RECT 2703.490 1614.420 2899.310 1614.560 ;
        RECT 2703.490 1614.360 2703.810 1614.420 ;
        RECT 2898.990 1614.360 2899.310 1614.420 ;
      LAYER via ;
        RECT 707.580 3306.880 707.840 3307.140 ;
        RECT 2703.520 3306.880 2703.780 3307.140 ;
        RECT 2703.520 1614.360 2703.780 1614.620 ;
        RECT 2899.020 1614.360 2899.280 1614.620 ;
      LAYER met2 ;
        RECT 707.580 3306.850 707.840 3307.170 ;
        RECT 2703.520 3306.850 2703.780 3307.170 ;
        RECT 707.640 3300.000 707.780 3306.850 ;
        RECT 707.580 3296.000 707.860 3300.000 ;
        RECT 2703.580 1614.650 2703.720 3306.850 ;
        RECT 2703.520 1614.330 2703.780 1614.650 ;
        RECT 2899.020 1614.330 2899.280 1614.650 ;
        RECT 2899.080 1613.485 2899.220 1614.330 ;
        RECT 2899.010 1613.115 2899.290 1613.485 ;
      LAYER via2 ;
        RECT 2899.010 1613.160 2899.290 1613.440 ;
      LAYER met3 ;
        RECT 2898.985 1613.450 2899.315 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2898.985 1613.150 2924.800 1613.450 ;
        RECT 2898.985 1613.135 2899.315 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 770.570 3308.440 770.890 3308.500 ;
        RECT 2703.950 3308.440 2704.270 3308.500 ;
        RECT 770.570 3308.300 2704.270 3308.440 ;
        RECT 770.570 3308.240 770.890 3308.300 ;
        RECT 2703.950 3308.240 2704.270 3308.300 ;
        RECT 2703.950 1849.160 2704.270 1849.220 ;
        RECT 2898.990 1849.160 2899.310 1849.220 ;
        RECT 2703.950 1849.020 2899.310 1849.160 ;
        RECT 2703.950 1848.960 2704.270 1849.020 ;
        RECT 2898.990 1848.960 2899.310 1849.020 ;
      LAYER via ;
        RECT 770.600 3308.240 770.860 3308.500 ;
        RECT 2703.980 3308.240 2704.240 3308.500 ;
        RECT 2703.980 1848.960 2704.240 1849.220 ;
        RECT 2899.020 1848.960 2899.280 1849.220 ;
      LAYER met2 ;
        RECT 770.600 3308.210 770.860 3308.530 ;
        RECT 2703.980 3308.210 2704.240 3308.530 ;
        RECT 770.660 3300.000 770.800 3308.210 ;
        RECT 770.600 3296.000 770.880 3300.000 ;
        RECT 2704.040 1849.250 2704.180 3308.210 ;
        RECT 2703.980 1848.930 2704.240 1849.250 ;
        RECT 2899.020 1848.930 2899.280 1849.250 ;
        RECT 2899.080 1848.085 2899.220 1848.930 ;
        RECT 2899.010 1847.715 2899.290 1848.085 ;
      LAYER via2 ;
        RECT 2899.010 1847.760 2899.290 1848.040 ;
      LAYER met3 ;
        RECT 2898.985 1848.050 2899.315 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2898.985 1847.750 2924.800 1848.050 ;
        RECT 2898.985 1847.735 2899.315 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 834.050 3309.120 834.370 3309.180 ;
        RECT 2704.410 3309.120 2704.730 3309.180 ;
        RECT 834.050 3308.980 2704.730 3309.120 ;
        RECT 834.050 3308.920 834.370 3308.980 ;
        RECT 2704.410 3308.920 2704.730 3308.980 ;
        RECT 2704.410 2083.760 2704.730 2083.820 ;
        RECT 2898.990 2083.760 2899.310 2083.820 ;
        RECT 2704.410 2083.620 2899.310 2083.760 ;
        RECT 2704.410 2083.560 2704.730 2083.620 ;
        RECT 2898.990 2083.560 2899.310 2083.620 ;
      LAYER via ;
        RECT 834.080 3308.920 834.340 3309.180 ;
        RECT 2704.440 3308.920 2704.700 3309.180 ;
        RECT 2704.440 2083.560 2704.700 2083.820 ;
        RECT 2899.020 2083.560 2899.280 2083.820 ;
      LAYER met2 ;
        RECT 834.080 3308.890 834.340 3309.210 ;
        RECT 2704.440 3308.890 2704.700 3309.210 ;
        RECT 834.140 3300.000 834.280 3308.890 ;
        RECT 834.080 3296.000 834.360 3300.000 ;
        RECT 2704.500 2083.850 2704.640 3308.890 ;
        RECT 2704.440 2083.530 2704.700 2083.850 ;
        RECT 2899.020 2083.530 2899.280 2083.850 ;
        RECT 2899.080 2082.685 2899.220 2083.530 ;
        RECT 2899.010 2082.315 2899.290 2082.685 ;
      LAYER via2 ;
        RECT 2899.010 2082.360 2899.290 2082.640 ;
      LAYER met3 ;
        RECT 2898.985 2082.650 2899.315 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2898.985 2082.350 2924.800 2082.650 ;
        RECT 2898.985 2082.335 2899.315 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 898.525 3296.045 898.695 3296.895 ;
      LAYER mcon ;
        RECT 898.525 3296.725 898.695 3296.895 ;
      LAYER met1 ;
        RECT 898.450 3296.880 898.770 3296.940 ;
        RECT 898.255 3296.740 898.770 3296.880 ;
        RECT 898.450 3296.680 898.770 3296.740 ;
        RECT 898.465 3296.200 898.755 3296.245 ;
        RECT 2700.730 3296.200 2701.050 3296.260 ;
        RECT 898.465 3296.060 2701.050 3296.200 ;
        RECT 898.465 3296.015 898.755 3296.060 ;
        RECT 2700.730 3296.000 2701.050 3296.060 ;
        RECT 2700.730 2318.360 2701.050 2318.420 ;
        RECT 2898.990 2318.360 2899.310 2318.420 ;
        RECT 2700.730 2318.220 2899.310 2318.360 ;
        RECT 2700.730 2318.160 2701.050 2318.220 ;
        RECT 2898.990 2318.160 2899.310 2318.220 ;
      LAYER via ;
        RECT 898.480 3296.680 898.740 3296.940 ;
        RECT 2700.760 3296.000 2701.020 3296.260 ;
        RECT 2700.760 2318.160 2701.020 2318.420 ;
        RECT 2899.020 2318.160 2899.280 2318.420 ;
      LAYER met2 ;
        RECT 897.100 3297.050 897.380 3300.000 ;
        RECT 897.100 3296.970 898.680 3297.050 ;
        RECT 897.100 3296.910 898.740 3296.970 ;
        RECT 897.100 3296.000 897.380 3296.910 ;
        RECT 898.480 3296.650 898.740 3296.910 ;
        RECT 2700.760 3295.970 2701.020 3296.290 ;
        RECT 2700.820 2318.450 2700.960 3295.970 ;
        RECT 2700.760 2318.130 2701.020 2318.450 ;
        RECT 2899.020 2318.130 2899.280 2318.450 ;
        RECT 2899.080 2317.285 2899.220 2318.130 ;
        RECT 2899.010 2316.915 2899.290 2317.285 ;
      LAYER via2 ;
        RECT 2899.010 2316.960 2899.290 2317.240 ;
      LAYER met3 ;
        RECT 2898.985 2317.250 2899.315 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2898.985 2316.950 2924.800 2317.250 ;
        RECT 2898.985 2316.935 2899.315 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 349.690 3307.675 349.970 3308.045 ;
        RECT 2901.310 3307.675 2901.590 3308.045 ;
        RECT 349.760 3300.000 349.900 3307.675 ;
        RECT 349.700 3296.000 349.980 3300.000 ;
        RECT 2901.380 146.725 2901.520 3307.675 ;
        RECT 2901.310 146.355 2901.590 146.725 ;
      LAYER via2 ;
        RECT 349.690 3307.720 349.970 3308.000 ;
        RECT 2901.310 3307.720 2901.590 3308.000 ;
        RECT 2901.310 146.400 2901.590 146.680 ;
      LAYER met3 ;
        RECT 349.665 3308.010 349.995 3308.025 ;
        RECT 2901.285 3308.010 2901.615 3308.025 ;
        RECT 349.665 3307.710 2901.615 3308.010 ;
        RECT 349.665 3307.695 349.995 3307.710 ;
        RECT 2901.285 3307.695 2901.615 3307.710 ;
        RECT 2901.285 146.690 2901.615 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2901.285 146.390 2924.800 146.690 ;
        RECT 2901.285 146.375 2901.615 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 981.250 3310.140 981.570 3310.200 ;
        RECT 2700.270 3310.140 2700.590 3310.200 ;
        RECT 981.250 3310.000 2700.590 3310.140 ;
        RECT 981.250 3309.940 981.570 3310.000 ;
        RECT 2700.270 3309.940 2700.590 3310.000 ;
        RECT 2700.270 2497.540 2700.590 2497.600 ;
        RECT 2899.910 2497.540 2900.230 2497.600 ;
        RECT 2700.270 2497.400 2900.230 2497.540 ;
        RECT 2700.270 2497.340 2700.590 2497.400 ;
        RECT 2899.910 2497.340 2900.230 2497.400 ;
      LAYER via ;
        RECT 981.280 3309.940 981.540 3310.200 ;
        RECT 2700.300 3309.940 2700.560 3310.200 ;
        RECT 2700.300 2497.340 2700.560 2497.600 ;
        RECT 2899.940 2497.340 2900.200 2497.600 ;
      LAYER met2 ;
        RECT 981.280 3309.910 981.540 3310.230 ;
        RECT 2700.300 3309.910 2700.560 3310.230 ;
        RECT 981.340 3300.000 981.480 3309.910 ;
        RECT 981.280 3296.000 981.560 3300.000 ;
        RECT 2700.360 2497.630 2700.500 3309.910 ;
        RECT 2700.300 2497.310 2700.560 2497.630 ;
        RECT 2899.940 2497.310 2900.200 2497.630 ;
        RECT 2900.000 2493.405 2900.140 2497.310 ;
        RECT 2899.930 2493.035 2900.210 2493.405 ;
      LAYER via2 ;
        RECT 2899.930 2493.080 2900.210 2493.360 ;
      LAYER met3 ;
        RECT 2899.905 2493.370 2900.235 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2899.905 2493.070 2924.800 2493.370 ;
        RECT 2899.905 2493.055 2900.235 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1908.225 3295.365 1908.395 3298.255 ;
      LAYER mcon ;
        RECT 1908.225 3298.085 1908.395 3298.255 ;
      LAYER met1 ;
        RECT 1044.270 3311.500 1044.590 3311.560 ;
        RECT 1908.150 3311.500 1908.470 3311.560 ;
        RECT 1044.270 3311.360 1908.470 3311.500 ;
        RECT 1044.270 3311.300 1044.590 3311.360 ;
        RECT 1908.150 3311.300 1908.470 3311.360 ;
        RECT 1908.150 3298.240 1908.470 3298.300 ;
        RECT 1907.955 3298.100 1908.470 3298.240 ;
        RECT 1908.150 3298.040 1908.470 3298.100 ;
        RECT 1908.165 3295.520 1908.455 3295.565 ;
        RECT 2900.830 3295.520 2901.150 3295.580 ;
        RECT 1908.165 3295.380 2901.150 3295.520 ;
        RECT 1908.165 3295.335 1908.455 3295.380 ;
        RECT 2900.830 3295.320 2901.150 3295.380 ;
      LAYER via ;
        RECT 1044.300 3311.300 1044.560 3311.560 ;
        RECT 1908.180 3311.300 1908.440 3311.560 ;
        RECT 1908.180 3298.040 1908.440 3298.300 ;
        RECT 2900.860 3295.320 2901.120 3295.580 ;
      LAYER met2 ;
        RECT 1044.300 3311.270 1044.560 3311.590 ;
        RECT 1908.180 3311.270 1908.440 3311.590 ;
        RECT 1044.360 3300.000 1044.500 3311.270 ;
        RECT 1044.300 3296.000 1044.580 3300.000 ;
        RECT 1908.240 3298.330 1908.380 3311.270 ;
        RECT 1908.180 3298.010 1908.440 3298.330 ;
        RECT 2900.860 3295.290 2901.120 3295.610 ;
        RECT 2900.920 2728.005 2901.060 3295.290 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
      LAYER met3 ;
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1109.130 3297.220 1109.450 3297.280 ;
        RECT 2709.010 3297.220 2709.330 3297.280 ;
        RECT 1109.130 3297.080 2709.330 3297.220 ;
        RECT 1109.130 3297.020 1109.450 3297.080 ;
        RECT 2709.010 3297.020 2709.330 3297.080 ;
        RECT 2709.010 2966.740 2709.330 2966.800 ;
        RECT 2900.370 2966.740 2900.690 2966.800 ;
        RECT 2709.010 2966.600 2900.690 2966.740 ;
        RECT 2709.010 2966.540 2709.330 2966.600 ;
        RECT 2900.370 2966.540 2900.690 2966.600 ;
      LAYER via ;
        RECT 1109.160 3297.020 1109.420 3297.280 ;
        RECT 2709.040 3297.020 2709.300 3297.280 ;
        RECT 2709.040 2966.540 2709.300 2966.800 ;
        RECT 2900.400 2966.540 2900.660 2966.800 ;
      LAYER met2 ;
        RECT 1107.780 3297.050 1108.060 3300.000 ;
        RECT 1109.160 3297.050 1109.420 3297.310 ;
        RECT 1107.780 3296.990 1109.420 3297.050 ;
        RECT 2709.040 3296.990 2709.300 3297.310 ;
        RECT 1107.780 3296.910 1109.360 3296.990 ;
        RECT 1107.780 3296.000 1108.060 3296.910 ;
        RECT 2709.100 2966.830 2709.240 3296.990 ;
        RECT 2709.040 2966.510 2709.300 2966.830 ;
        RECT 2900.400 2966.510 2900.660 2966.830 ;
        RECT 2900.460 2962.605 2900.600 2966.510 ;
        RECT 2900.390 2962.235 2900.670 2962.605 ;
      LAYER via2 ;
        RECT 2900.390 2962.280 2900.670 2962.560 ;
      LAYER met3 ;
        RECT 2900.365 2962.570 2900.695 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.365 2962.270 2924.800 2962.570 ;
        RECT 2900.365 2962.255 2900.695 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1172.610 3297.900 1172.930 3297.960 ;
        RECT 2709.470 3297.900 2709.790 3297.960 ;
        RECT 1172.610 3297.760 2709.790 3297.900 ;
        RECT 1172.610 3297.700 1172.930 3297.760 ;
        RECT 2709.470 3297.700 2709.790 3297.760 ;
        RECT 2709.470 3201.340 2709.790 3201.400 ;
        RECT 2900.370 3201.340 2900.690 3201.400 ;
        RECT 2709.470 3201.200 2900.690 3201.340 ;
        RECT 2709.470 3201.140 2709.790 3201.200 ;
        RECT 2900.370 3201.140 2900.690 3201.200 ;
      LAYER via ;
        RECT 1172.640 3297.700 1172.900 3297.960 ;
        RECT 2709.500 3297.700 2709.760 3297.960 ;
        RECT 2709.500 3201.140 2709.760 3201.400 ;
        RECT 2900.400 3201.140 2900.660 3201.400 ;
      LAYER met2 ;
        RECT 1170.800 3297.730 1171.080 3300.000 ;
        RECT 1172.640 3297.730 1172.900 3297.990 ;
        RECT 1170.800 3297.670 1172.900 3297.730 ;
        RECT 2709.500 3297.670 2709.760 3297.990 ;
        RECT 1170.800 3297.590 1172.840 3297.670 ;
        RECT 1170.800 3296.000 1171.080 3297.590 ;
        RECT 2709.560 3201.430 2709.700 3297.670 ;
        RECT 2709.500 3201.110 2709.760 3201.430 ;
        RECT 2900.400 3201.110 2900.660 3201.430 ;
        RECT 2900.460 3197.205 2900.600 3201.110 ;
        RECT 2900.390 3196.835 2900.670 3197.205 ;
      LAYER via2 ;
        RECT 2900.390 3196.880 2900.670 3197.160 ;
      LAYER met3 ;
        RECT 2900.365 3197.170 2900.695 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.365 3196.870 2924.800 3197.170 ;
        RECT 2900.365 3196.855 2900.695 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1234.710 3429.480 1235.030 3429.540 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 1234.710 3429.340 2901.150 3429.480 ;
        RECT 1234.710 3429.280 1235.030 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 1234.740 3429.280 1235.000 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 1234.740 3429.250 1235.000 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 1233.820 3299.770 1234.100 3300.000 ;
        RECT 1234.800 3299.770 1234.940 3429.250 ;
        RECT 1233.820 3299.630 1234.940 3299.770 ;
        RECT 1233.820 3296.000 1234.100 3299.630 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1296.810 3502.240 1297.130 3502.300 ;
        RECT 2717.290 3502.240 2717.610 3502.300 ;
        RECT 1296.810 3502.100 2717.610 3502.240 ;
        RECT 1296.810 3502.040 1297.130 3502.100 ;
        RECT 2717.290 3502.040 2717.610 3502.100 ;
      LAYER via ;
        RECT 1296.840 3502.040 1297.100 3502.300 ;
        RECT 2717.320 3502.040 2717.580 3502.300 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3502.330 2717.520 3517.600 ;
        RECT 1296.840 3502.010 1297.100 3502.330 ;
        RECT 2717.320 3502.010 2717.580 3502.330 ;
        RECT 1296.900 3300.000 1297.040 3502.010 ;
        RECT 1296.840 3296.000 1297.120 3300.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1365.810 3503.940 1366.130 3504.000 ;
        RECT 2392.530 3503.940 2392.850 3504.000 ;
        RECT 1365.810 3503.800 2392.850 3503.940 ;
        RECT 1365.810 3503.740 1366.130 3503.800 ;
        RECT 2392.530 3503.740 2392.850 3503.800 ;
      LAYER via ;
        RECT 1365.840 3503.740 1366.100 3504.000 ;
        RECT 2392.560 3503.740 2392.820 3504.000 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3504.030 2392.760 3517.600 ;
        RECT 1365.840 3503.710 1366.100 3504.030 ;
        RECT 2392.560 3503.710 2392.820 3504.030 ;
        RECT 1365.900 3300.450 1366.040 3503.710 ;
        RECT 1363.140 3300.310 1366.040 3300.450 ;
        RECT 1360.320 3299.090 1360.600 3300.000 ;
        RECT 1363.140 3299.090 1363.280 3300.310 ;
        RECT 1360.320 3298.950 1363.280 3299.090 ;
        RECT 1360.320 3296.000 1360.600 3298.950 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1427.910 3500.880 1428.230 3500.940 ;
        RECT 2068.230 3500.880 2068.550 3500.940 ;
        RECT 1427.910 3500.740 2068.550 3500.880 ;
        RECT 1427.910 3500.680 1428.230 3500.740 ;
        RECT 2068.230 3500.680 2068.550 3500.740 ;
      LAYER via ;
        RECT 1427.940 3500.680 1428.200 3500.940 ;
        RECT 2068.260 3500.680 2068.520 3500.940 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3500.970 2068.460 3517.600 ;
        RECT 1427.940 3500.650 1428.200 3500.970 ;
        RECT 2068.260 3500.650 2068.520 3500.970 ;
        RECT 1423.340 3299.090 1423.620 3300.000 ;
        RECT 1428.000 3299.090 1428.140 3500.650 ;
        RECT 1423.340 3298.950 1428.140 3299.090 ;
        RECT 1423.340 3296.000 1423.620 3298.950 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1500.205 3497.665 1500.375 3499.195 ;
        RECT 1525.505 3497.665 1525.675 3499.535 ;
      LAYER mcon ;
        RECT 1525.505 3499.365 1525.675 3499.535 ;
        RECT 1500.205 3499.025 1500.375 3499.195 ;
      LAYER met1 ;
        RECT 1525.445 3499.520 1525.735 3499.565 ;
        RECT 1743.930 3499.520 1744.250 3499.580 ;
        RECT 1525.445 3499.380 1744.250 3499.520 ;
        RECT 1525.445 3499.335 1525.735 3499.380 ;
        RECT 1743.930 3499.320 1744.250 3499.380 ;
        RECT 1490.010 3499.180 1490.330 3499.240 ;
        RECT 1500.145 3499.180 1500.435 3499.225 ;
        RECT 1490.010 3499.040 1500.435 3499.180 ;
        RECT 1490.010 3498.980 1490.330 3499.040 ;
        RECT 1500.145 3498.995 1500.435 3499.040 ;
        RECT 1500.145 3497.820 1500.435 3497.865 ;
        RECT 1525.445 3497.820 1525.735 3497.865 ;
        RECT 1500.145 3497.680 1525.735 3497.820 ;
        RECT 1500.145 3497.635 1500.435 3497.680 ;
        RECT 1525.445 3497.635 1525.735 3497.680 ;
      LAYER via ;
        RECT 1743.960 3499.320 1744.220 3499.580 ;
        RECT 1490.040 3498.980 1490.300 3499.240 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3499.610 1744.160 3517.600 ;
        RECT 1743.960 3499.290 1744.220 3499.610 ;
        RECT 1490.040 3498.950 1490.300 3499.270 ;
        RECT 1486.360 3299.090 1486.640 3300.000 ;
        RECT 1490.100 3299.090 1490.240 3498.950 ;
        RECT 1486.360 3298.950 1490.240 3299.090 ;
        RECT 1486.360 3296.000 1486.640 3298.950 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.170 3498.500 1419.490 3498.560 ;
        RECT 1545.670 3498.500 1545.990 3498.560 ;
        RECT 1419.170 3498.360 1545.990 3498.500 ;
        RECT 1419.170 3498.300 1419.490 3498.360 ;
        RECT 1545.670 3498.300 1545.990 3498.360 ;
      LAYER via ;
        RECT 1419.200 3498.300 1419.460 3498.560 ;
        RECT 1545.700 3498.300 1545.960 3498.560 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3498.590 1419.400 3517.600 ;
        RECT 1419.200 3498.270 1419.460 3498.590 ;
        RECT 1545.700 3498.270 1545.960 3498.590 ;
        RECT 1545.760 3299.090 1545.900 3498.270 ;
        RECT 1549.840 3299.090 1550.120 3300.000 ;
        RECT 1545.760 3298.950 1550.120 3299.090 ;
        RECT 1549.840 3296.000 1550.120 3298.950 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 412.690 3308.100 413.010 3308.160 ;
        RECT 778.390 3308.100 778.710 3308.160 ;
        RECT 412.690 3307.960 778.710 3308.100 ;
        RECT 412.690 3307.900 413.010 3307.960 ;
        RECT 778.390 3307.900 778.710 3307.960 ;
      LAYER via ;
        RECT 412.720 3307.900 412.980 3308.160 ;
        RECT 778.420 3307.900 778.680 3308.160 ;
      LAYER met2 ;
        RECT 412.720 3307.870 412.980 3308.190 ;
        RECT 778.420 3307.870 778.680 3308.190 ;
        RECT 412.780 3300.000 412.920 3307.870 ;
        RECT 412.720 3296.000 413.000 3300.000 ;
        RECT 778.480 3297.165 778.620 3307.870 ;
        RECT 778.410 3296.795 778.690 3297.165 ;
        RECT 2901.770 3295.435 2902.050 3295.805 ;
        RECT 2901.840 381.325 2901.980 3295.435 ;
        RECT 2901.770 380.955 2902.050 381.325 ;
      LAYER via2 ;
        RECT 778.410 3296.840 778.690 3297.120 ;
        RECT 2901.770 3295.480 2902.050 3295.760 ;
        RECT 2901.770 381.000 2902.050 381.280 ;
      LAYER met3 ;
        RECT 778.385 3297.130 778.715 3297.145 ;
        RECT 778.385 3296.815 778.930 3297.130 ;
        RECT 778.630 3295.770 778.930 3296.815 ;
        RECT 2901.745 3295.770 2902.075 3295.785 ;
        RECT 778.630 3295.470 2902.075 3295.770 ;
        RECT 2901.745 3295.455 2902.075 3295.470 ;
        RECT 2901.745 381.290 2902.075 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2901.745 380.990 2924.800 381.290 ;
        RECT 2901.745 380.975 2902.075 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1094.870 3499.860 1095.190 3499.920 ;
        RECT 1607.770 3499.860 1608.090 3499.920 ;
        RECT 1094.870 3499.720 1608.090 3499.860 ;
        RECT 1094.870 3499.660 1095.190 3499.720 ;
        RECT 1607.770 3499.660 1608.090 3499.720 ;
      LAYER via ;
        RECT 1094.900 3499.660 1095.160 3499.920 ;
        RECT 1607.800 3499.660 1608.060 3499.920 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3499.950 1095.100 3517.600 ;
        RECT 1094.900 3499.630 1095.160 3499.950 ;
        RECT 1607.800 3499.630 1608.060 3499.950 ;
        RECT 1607.860 3300.450 1608.000 3499.630 ;
        RECT 1607.860 3300.310 1610.300 3300.450 ;
        RECT 1610.160 3299.090 1610.300 3300.310 ;
        RECT 1612.860 3299.090 1613.140 3300.000 ;
        RECT 1610.160 3298.950 1613.140 3299.090 ;
        RECT 1612.860 3296.000 1613.140 3298.950 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 770.570 3504.960 770.890 3505.020 ;
        RECT 1669.870 3504.960 1670.190 3505.020 ;
        RECT 770.570 3504.820 1670.190 3504.960 ;
        RECT 770.570 3504.760 770.890 3504.820 ;
        RECT 1669.870 3504.760 1670.190 3504.820 ;
      LAYER via ;
        RECT 770.600 3504.760 770.860 3505.020 ;
        RECT 1669.900 3504.760 1670.160 3505.020 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3505.050 770.800 3517.600 ;
        RECT 770.600 3504.730 770.860 3505.050 ;
        RECT 1669.900 3504.730 1670.160 3505.050 ;
        RECT 1669.960 3300.450 1670.100 3504.730 ;
        RECT 1669.960 3300.310 1673.780 3300.450 ;
        RECT 1673.640 3299.090 1673.780 3300.310 ;
        RECT 1675.880 3299.090 1676.160 3300.000 ;
        RECT 1673.640 3298.950 1676.160 3299.090 ;
        RECT 1675.880 3296.000 1676.160 3298.950 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3503.260 446.130 3503.320 ;
        RECT 1739.330 3503.260 1739.650 3503.320 ;
        RECT 445.810 3503.120 1739.650 3503.260 ;
        RECT 445.810 3503.060 446.130 3503.120 ;
        RECT 1739.330 3503.060 1739.650 3503.120 ;
      LAYER via ;
        RECT 445.840 3503.060 446.100 3503.320 ;
        RECT 1739.360 3503.060 1739.620 3503.320 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3503.350 446.040 3517.600 ;
        RECT 445.840 3503.030 446.100 3503.350 ;
        RECT 1739.360 3503.030 1739.620 3503.350 ;
        RECT 1738.900 3299.770 1739.180 3300.000 ;
        RECT 1739.420 3299.770 1739.560 3503.030 ;
        RECT 1738.900 3299.630 1739.560 3299.770 ;
        RECT 1738.900 3296.000 1739.180 3299.630 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3501.560 121.830 3501.620 ;
        RECT 1800.970 3501.560 1801.290 3501.620 ;
        RECT 121.510 3501.420 1801.290 3501.560 ;
        RECT 121.510 3501.360 121.830 3501.420 ;
        RECT 1800.970 3501.360 1801.290 3501.420 ;
      LAYER via ;
        RECT 121.540 3501.360 121.800 3501.620 ;
        RECT 1801.000 3501.360 1801.260 3501.620 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3501.650 121.740 3517.600 ;
        RECT 121.540 3501.330 121.800 3501.650 ;
        RECT 1801.000 3501.330 1801.260 3501.650 ;
        RECT 1801.060 3299.770 1801.200 3501.330 ;
        RECT 1802.380 3299.770 1802.660 3300.000 ;
        RECT 1801.060 3299.630 1802.660 3299.770 ;
        RECT 1802.380 3296.000 1802.660 3299.630 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 1863.070 3339.720 1863.390 3339.780 ;
        RECT 17.090 3339.580 1863.390 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 1863.070 3339.520 1863.390 3339.580 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 1863.100 3339.520 1863.360 3339.780 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 1863.100 3339.490 1863.360 3339.810 ;
        RECT 1863.160 3299.090 1863.300 3339.490 ;
        RECT 1865.400 3299.090 1865.680 3300.000 ;
        RECT 1863.160 3298.950 1865.680 3299.090 ;
        RECT 1865.400 3296.000 1865.680 3298.950 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1926.625 3295.025 1926.795 3298.255 ;
      LAYER mcon ;
        RECT 1926.625 3298.085 1926.795 3298.255 ;
      LAYER met1 ;
        RECT 1926.550 3298.240 1926.870 3298.300 ;
        RECT 1926.355 3298.100 1926.870 3298.240 ;
        RECT 1926.550 3298.040 1926.870 3298.100 ;
        RECT 25.370 3295.180 25.690 3295.240 ;
        RECT 1926.565 3295.180 1926.855 3295.225 ;
        RECT 25.370 3295.040 1926.855 3295.180 ;
        RECT 25.370 3294.980 25.690 3295.040 ;
        RECT 1926.565 3294.995 1926.855 3295.040 ;
        RECT 13.870 3052.420 14.190 3052.480 ;
        RECT 25.370 3052.420 25.690 3052.480 ;
        RECT 13.870 3052.280 25.690 3052.420 ;
        RECT 13.870 3052.220 14.190 3052.280 ;
        RECT 25.370 3052.220 25.690 3052.280 ;
      LAYER via ;
        RECT 1926.580 3298.040 1926.840 3298.300 ;
        RECT 25.400 3294.980 25.660 3295.240 ;
        RECT 13.900 3052.220 14.160 3052.480 ;
        RECT 25.400 3052.220 25.660 3052.480 ;
      LAYER met2 ;
        RECT 1928.420 3298.410 1928.700 3300.000 ;
        RECT 1926.640 3298.330 1928.700 3298.410 ;
        RECT 1926.580 3298.270 1928.700 3298.330 ;
        RECT 1926.580 3298.010 1926.840 3298.270 ;
        RECT 1928.420 3296.000 1928.700 3298.270 ;
        RECT 25.400 3294.950 25.660 3295.270 ;
        RECT 25.460 3052.510 25.600 3294.950 ;
        RECT 13.900 3052.365 14.160 3052.510 ;
        RECT 13.890 3051.995 14.170 3052.365 ;
        RECT 25.400 3052.190 25.660 3052.510 ;
      LAYER via2 ;
        RECT 13.890 3052.040 14.170 3052.320 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 13.865 3052.330 14.195 3052.345 ;
        RECT -4.800 3052.030 14.195 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 13.865 3052.015 14.195 3052.030 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1169.390 3311.840 1169.710 3311.900 ;
        RECT 1991.870 3311.840 1992.190 3311.900 ;
        RECT 1169.390 3311.700 1992.190 3311.840 ;
        RECT 1169.390 3311.640 1169.710 3311.700 ;
        RECT 1991.870 3311.640 1992.190 3311.700 ;
        RECT 16.170 3297.900 16.490 3297.960 ;
        RECT 1169.390 3297.900 1169.710 3297.960 ;
        RECT 16.170 3297.760 1169.710 3297.900 ;
        RECT 16.170 3297.700 16.490 3297.760 ;
        RECT 1169.390 3297.700 1169.710 3297.760 ;
      LAYER via ;
        RECT 1169.420 3311.640 1169.680 3311.900 ;
        RECT 1991.900 3311.640 1992.160 3311.900 ;
        RECT 16.200 3297.700 16.460 3297.960 ;
        RECT 1169.420 3297.700 1169.680 3297.960 ;
      LAYER met2 ;
        RECT 1169.420 3311.610 1169.680 3311.930 ;
        RECT 1991.900 3311.610 1992.160 3311.930 ;
        RECT 1169.480 3297.990 1169.620 3311.610 ;
        RECT 1991.960 3300.000 1992.100 3311.610 ;
        RECT 16.200 3297.670 16.460 3297.990 ;
        RECT 1169.420 3297.670 1169.680 3297.990 ;
        RECT 16.260 2765.405 16.400 3297.670 ;
        RECT 1991.900 3296.000 1992.180 3300.000 ;
        RECT 16.190 2765.035 16.470 2765.405 ;
      LAYER via2 ;
        RECT 16.190 2765.080 16.470 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 16.165 2765.370 16.495 2765.385 ;
        RECT -4.800 2765.070 16.495 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 16.165 2765.055 16.495 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2053.585 3294.345 2053.755 3298.255 ;
      LAYER mcon ;
        RECT 2053.585 3298.085 2053.755 3298.255 ;
      LAYER met1 ;
        RECT 2053.510 3298.240 2053.830 3298.300 ;
        RECT 2053.315 3298.100 2053.830 3298.240 ;
        RECT 2053.510 3298.040 2053.830 3298.100 ;
        RECT 24.910 3294.500 25.230 3294.560 ;
        RECT 2053.525 3294.500 2053.815 3294.545 ;
        RECT 24.910 3294.360 2053.815 3294.500 ;
        RECT 24.910 3294.300 25.230 3294.360 ;
        RECT 2053.525 3294.315 2053.815 3294.360 ;
        RECT 13.870 2483.600 14.190 2483.660 ;
        RECT 24.910 2483.600 25.230 2483.660 ;
        RECT 13.870 2483.460 25.230 2483.600 ;
        RECT 13.870 2483.400 14.190 2483.460 ;
        RECT 24.910 2483.400 25.230 2483.460 ;
      LAYER via ;
        RECT 2053.540 3298.040 2053.800 3298.300 ;
        RECT 24.940 3294.300 25.200 3294.560 ;
        RECT 13.900 2483.400 14.160 2483.660 ;
        RECT 24.940 2483.400 25.200 2483.660 ;
      LAYER met2 ;
        RECT 2054.920 3298.410 2055.200 3300.000 ;
        RECT 2053.600 3298.330 2055.200 3298.410 ;
        RECT 2053.540 3298.270 2055.200 3298.330 ;
        RECT 2053.540 3298.010 2053.800 3298.270 ;
        RECT 2054.920 3296.000 2055.200 3298.270 ;
        RECT 24.940 3294.270 25.200 3294.590 ;
        RECT 25.000 2483.690 25.140 3294.270 ;
        RECT 13.900 2483.370 14.160 2483.690 ;
        RECT 24.940 2483.370 25.200 2483.690 ;
        RECT 13.960 2477.765 14.100 2483.370 ;
        RECT 13.890 2477.395 14.170 2477.765 ;
      LAYER via2 ;
        RECT 13.890 2477.440 14.170 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 13.865 2477.730 14.195 2477.745 ;
        RECT -4.800 2477.430 14.195 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 13.865 2477.415 14.195 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2116.145 3293.325 2116.315 3298.255 ;
      LAYER mcon ;
        RECT 2116.145 3298.085 2116.315 3298.255 ;
      LAYER met1 ;
        RECT 2116.070 3298.240 2116.390 3298.300 ;
        RECT 2115.875 3298.100 2116.390 3298.240 ;
        RECT 2116.070 3298.040 2116.390 3298.100 ;
        RECT 24.450 3293.480 24.770 3293.540 ;
        RECT 2116.085 3293.480 2116.375 3293.525 ;
        RECT 24.450 3293.340 2116.375 3293.480 ;
        RECT 24.450 3293.280 24.770 3293.340 ;
        RECT 2116.085 3293.295 2116.375 3293.340 ;
        RECT 13.870 2193.920 14.190 2193.980 ;
        RECT 24.450 2193.920 24.770 2193.980 ;
        RECT 13.870 2193.780 24.770 2193.920 ;
        RECT 13.870 2193.720 14.190 2193.780 ;
        RECT 24.450 2193.720 24.770 2193.780 ;
      LAYER via ;
        RECT 2116.100 3298.040 2116.360 3298.300 ;
        RECT 24.480 3293.280 24.740 3293.540 ;
        RECT 13.900 2193.720 14.160 2193.980 ;
        RECT 24.480 2193.720 24.740 2193.980 ;
      LAYER met2 ;
        RECT 2117.940 3298.410 2118.220 3300.000 ;
        RECT 2116.160 3298.330 2118.220 3298.410 ;
        RECT 2116.100 3298.270 2118.220 3298.330 ;
        RECT 2116.100 3298.010 2116.360 3298.270 ;
        RECT 2117.940 3296.000 2118.220 3298.270 ;
        RECT 24.480 3293.250 24.740 3293.570 ;
        RECT 24.540 2194.010 24.680 3293.250 ;
        RECT 13.900 2193.690 14.160 2194.010 ;
        RECT 24.480 2193.690 24.740 2194.010 ;
        RECT 13.960 2190.125 14.100 2193.690 ;
        RECT 13.890 2189.755 14.170 2190.125 ;
      LAYER via2 ;
        RECT 13.890 2189.800 14.170 2190.080 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 13.865 2190.090 14.195 2190.105 ;
        RECT -4.800 2189.790 14.195 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 13.865 2189.775 14.195 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 3306.400 20.630 3306.460 ;
        RECT 2180.930 3306.400 2181.250 3306.460 ;
        RECT 20.310 3306.260 2181.250 3306.400 ;
        RECT 20.310 3306.200 20.630 3306.260 ;
        RECT 2180.930 3306.200 2181.250 3306.260 ;
      LAYER via ;
        RECT 20.340 3306.200 20.600 3306.460 ;
        RECT 2180.960 3306.200 2181.220 3306.460 ;
      LAYER met2 ;
        RECT 20.340 3306.170 20.600 3306.490 ;
        RECT 2180.960 3306.170 2181.220 3306.490 ;
        RECT 20.400 1903.165 20.540 3306.170 ;
        RECT 2181.020 3300.000 2181.160 3306.170 ;
        RECT 2180.960 3296.000 2181.240 3300.000 ;
        RECT 20.330 1902.795 20.610 1903.165 ;
      LAYER via2 ;
        RECT 20.330 1902.840 20.610 1903.120 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 20.305 1903.130 20.635 1903.145 ;
        RECT -4.800 1902.830 20.635 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 20.305 1902.815 20.635 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 476.170 3311.840 476.490 3311.900 ;
        RECT 1162.950 3311.840 1163.270 3311.900 ;
        RECT 476.170 3311.700 1163.270 3311.840 ;
        RECT 476.170 3311.640 476.490 3311.700 ;
        RECT 1162.950 3311.640 1163.270 3311.700 ;
      LAYER via ;
        RECT 476.200 3311.640 476.460 3311.900 ;
        RECT 1162.980 3311.640 1163.240 3311.900 ;
      LAYER met2 ;
        RECT 476.200 3311.610 476.460 3311.930 ;
        RECT 1162.980 3311.610 1163.240 3311.930 ;
        RECT 476.260 3300.000 476.400 3311.610 ;
        RECT 1163.040 3301.245 1163.180 3311.610 ;
        RECT 1162.970 3300.875 1163.250 3301.245 ;
        RECT 2902.690 3300.875 2902.970 3301.245 ;
        RECT 476.200 3296.000 476.480 3300.000 ;
        RECT 2902.760 615.925 2902.900 3300.875 ;
        RECT 2902.690 615.555 2902.970 615.925 ;
      LAYER via2 ;
        RECT 1162.970 3300.920 1163.250 3301.200 ;
        RECT 2902.690 3300.920 2902.970 3301.200 ;
        RECT 2902.690 615.600 2902.970 615.880 ;
      LAYER met3 ;
        RECT 1162.945 3301.210 1163.275 3301.225 ;
        RECT 2902.665 3301.210 2902.995 3301.225 ;
        RECT 1162.945 3300.910 2902.995 3301.210 ;
        RECT 1162.945 3300.895 1163.275 3300.910 ;
        RECT 2902.665 3300.895 2902.995 3300.910 ;
        RECT 2902.665 615.890 2902.995 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2902.665 615.590 2924.800 615.890 ;
        RECT 2902.665 615.575 2902.995 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1069.110 3310.820 1069.430 3310.880 ;
        RECT 2244.410 3310.820 2244.730 3310.880 ;
        RECT 1069.110 3310.680 2244.730 3310.820 ;
        RECT 1069.110 3310.620 1069.430 3310.680 ;
        RECT 2244.410 3310.620 2244.730 3310.680 ;
        RECT 19.390 3305.040 19.710 3305.100 ;
        RECT 1069.110 3305.040 1069.430 3305.100 ;
        RECT 19.390 3304.900 1069.430 3305.040 ;
        RECT 19.390 3304.840 19.710 3304.900 ;
        RECT 1069.110 3304.840 1069.430 3304.900 ;
      LAYER via ;
        RECT 1069.140 3310.620 1069.400 3310.880 ;
        RECT 2244.440 3310.620 2244.700 3310.880 ;
        RECT 19.420 3304.840 19.680 3305.100 ;
        RECT 1069.140 3304.840 1069.400 3305.100 ;
      LAYER met2 ;
        RECT 1069.140 3310.590 1069.400 3310.910 ;
        RECT 2244.440 3310.590 2244.700 3310.910 ;
        RECT 1069.200 3305.130 1069.340 3310.590 ;
        RECT 19.420 3304.810 19.680 3305.130 ;
        RECT 1069.140 3304.810 1069.400 3305.130 ;
        RECT 19.480 1615.525 19.620 3304.810 ;
        RECT 2244.500 3300.000 2244.640 3310.590 ;
        RECT 2244.440 3296.000 2244.720 3300.000 ;
        RECT 19.410 1615.155 19.690 1615.525 ;
      LAYER via2 ;
        RECT 19.410 1615.200 19.690 1615.480 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 19.385 1615.490 19.715 1615.505 ;
        RECT -4.800 1615.190 19.715 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 19.385 1615.175 19.715 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 46.990 3305.720 47.310 3305.780 ;
        RECT 2307.430 3305.720 2307.750 3305.780 ;
        RECT 46.990 3305.580 2307.750 3305.720 ;
        RECT 46.990 3305.520 47.310 3305.580 ;
        RECT 2307.430 3305.520 2307.750 3305.580 ;
        RECT 16.630 1400.700 16.950 1400.760 ;
        RECT 46.990 1400.700 47.310 1400.760 ;
        RECT 16.630 1400.560 47.310 1400.700 ;
        RECT 16.630 1400.500 16.950 1400.560 ;
        RECT 46.990 1400.500 47.310 1400.560 ;
      LAYER via ;
        RECT 47.020 3305.520 47.280 3305.780 ;
        RECT 2307.460 3305.520 2307.720 3305.780 ;
        RECT 16.660 1400.500 16.920 1400.760 ;
        RECT 47.020 1400.500 47.280 1400.760 ;
      LAYER met2 ;
        RECT 47.020 3305.490 47.280 3305.810 ;
        RECT 2307.460 3305.490 2307.720 3305.810 ;
        RECT 47.080 1400.790 47.220 3305.490 ;
        RECT 2307.520 3300.000 2307.660 3305.490 ;
        RECT 2307.460 3296.000 2307.740 3300.000 ;
        RECT 16.660 1400.645 16.920 1400.790 ;
        RECT 16.650 1400.275 16.930 1400.645 ;
        RECT 47.020 1400.470 47.280 1400.790 ;
      LAYER via2 ;
        RECT 16.650 1400.320 16.930 1400.600 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 16.625 1400.610 16.955 1400.625 ;
        RECT -4.800 1400.310 16.955 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 16.625 1400.295 16.955 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 293.550 3300.960 293.870 3301.020 ;
        RECT 2370.450 3300.960 2370.770 3301.020 ;
        RECT 293.550 3300.820 2370.770 3300.960 ;
        RECT 293.550 3300.760 293.870 3300.820 ;
        RECT 2370.450 3300.760 2370.770 3300.820 ;
        RECT 16.630 1186.840 16.950 1186.900 ;
        RECT 293.550 1186.840 293.870 1186.900 ;
        RECT 16.630 1186.700 293.870 1186.840 ;
        RECT 16.630 1186.640 16.950 1186.700 ;
        RECT 293.550 1186.640 293.870 1186.700 ;
      LAYER via ;
        RECT 293.580 3300.760 293.840 3301.020 ;
        RECT 2370.480 3300.760 2370.740 3301.020 ;
        RECT 16.660 1186.640 16.920 1186.900 ;
        RECT 293.580 1186.640 293.840 1186.900 ;
      LAYER met2 ;
        RECT 293.580 3300.730 293.840 3301.050 ;
        RECT 2370.480 3300.730 2370.740 3301.050 ;
        RECT 293.640 1186.930 293.780 3300.730 ;
        RECT 2370.540 3300.000 2370.680 3300.730 ;
        RECT 2370.480 3296.000 2370.760 3300.000 ;
        RECT 16.660 1186.610 16.920 1186.930 ;
        RECT 293.580 1186.610 293.840 1186.930 ;
        RECT 16.720 1185.085 16.860 1186.610 ;
        RECT 16.650 1184.715 16.930 1185.085 ;
      LAYER via2 ;
        RECT 16.650 1184.760 16.930 1185.040 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 16.625 1185.050 16.955 1185.065 ;
        RECT -4.800 1184.750 16.955 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 16.625 1184.735 16.955 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 45.610 3305.380 45.930 3305.440 ;
        RECT 2433.930 3305.380 2434.250 3305.440 ;
        RECT 45.610 3305.240 2434.250 3305.380 ;
        RECT 45.610 3305.180 45.930 3305.240 ;
        RECT 2433.930 3305.180 2434.250 3305.240 ;
        RECT 16.630 972.640 16.950 972.700 ;
        RECT 45.610 972.640 45.930 972.700 ;
        RECT 16.630 972.500 45.930 972.640 ;
        RECT 16.630 972.440 16.950 972.500 ;
        RECT 45.610 972.440 45.930 972.500 ;
      LAYER via ;
        RECT 45.640 3305.180 45.900 3305.440 ;
        RECT 2433.960 3305.180 2434.220 3305.440 ;
        RECT 16.660 972.440 16.920 972.700 ;
        RECT 45.640 972.440 45.900 972.700 ;
      LAYER met2 ;
        RECT 45.640 3305.150 45.900 3305.470 ;
        RECT 2433.960 3305.150 2434.220 3305.470 ;
        RECT 45.700 972.730 45.840 3305.150 ;
        RECT 2434.020 3300.000 2434.160 3305.150 ;
        RECT 2433.960 3296.000 2434.240 3300.000 ;
        RECT 16.660 972.410 16.920 972.730 ;
        RECT 45.640 972.410 45.900 972.730 ;
        RECT 16.720 969.525 16.860 972.410 ;
        RECT 16.650 969.155 16.930 969.525 ;
      LAYER via2 ;
        RECT 16.650 969.200 16.930 969.480 ;
      LAYER met3 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 16.625 969.490 16.955 969.505 ;
        RECT -4.800 969.190 16.955 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 16.625 969.175 16.955 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.870 3309.035 20.150 3309.405 ;
        RECT 2496.970 3309.035 2497.250 3309.405 ;
        RECT 19.940 753.965 20.080 3309.035 ;
        RECT 2497.040 3300.000 2497.180 3309.035 ;
        RECT 2496.980 3296.000 2497.260 3300.000 ;
        RECT 19.870 753.595 20.150 753.965 ;
      LAYER via2 ;
        RECT 19.870 3309.080 20.150 3309.360 ;
        RECT 2496.970 3309.080 2497.250 3309.360 ;
        RECT 19.870 753.640 20.150 753.920 ;
      LAYER met3 ;
        RECT 19.845 3309.370 20.175 3309.385 ;
        RECT 2496.945 3309.370 2497.275 3309.385 ;
        RECT 19.845 3309.070 2497.275 3309.370 ;
        RECT 19.845 3309.055 20.175 3309.070 ;
        RECT 2496.945 3309.055 2497.275 3309.070 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 19.845 753.930 20.175 753.945 ;
        RECT -4.800 753.630 20.175 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 19.845 753.615 20.175 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.950 3308.355 19.230 3308.725 ;
        RECT 2559.990 3308.355 2560.270 3308.725 ;
        RECT 19.020 538.405 19.160 3308.355 ;
        RECT 2560.060 3300.000 2560.200 3308.355 ;
        RECT 2560.000 3296.000 2560.280 3300.000 ;
        RECT 18.950 538.035 19.230 538.405 ;
      LAYER via2 ;
        RECT 18.950 3308.400 19.230 3308.680 ;
        RECT 2559.990 3308.400 2560.270 3308.680 ;
        RECT 18.950 538.080 19.230 538.360 ;
      LAYER met3 ;
        RECT 18.925 3308.690 19.255 3308.705 ;
        RECT 2559.965 3308.690 2560.295 3308.705 ;
        RECT 18.925 3308.390 2560.295 3308.690 ;
        RECT 18.925 3308.375 19.255 3308.390 ;
        RECT 2559.965 3308.375 2560.295 3308.390 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 18.925 538.370 19.255 538.385 ;
        RECT -4.800 538.070 19.255 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 18.925 538.055 19.255 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 322.900 14.190 322.960 ;
        RECT 23.990 322.900 24.310 322.960 ;
        RECT 13.870 322.760 24.310 322.900 ;
        RECT 13.870 322.700 14.190 322.760 ;
        RECT 23.990 322.700 24.310 322.760 ;
      LAYER via ;
        RECT 13.900 322.700 14.160 322.960 ;
        RECT 24.020 322.700 24.280 322.960 ;
      LAYER met2 ;
        RECT 24.010 3305.635 24.290 3306.005 ;
        RECT 2623.010 3305.635 2623.290 3306.005 ;
        RECT 24.080 322.990 24.220 3305.635 ;
        RECT 2623.080 3300.000 2623.220 3305.635 ;
        RECT 2623.020 3296.000 2623.300 3300.000 ;
        RECT 13.900 322.845 14.160 322.990 ;
        RECT 13.890 322.475 14.170 322.845 ;
        RECT 24.020 322.670 24.280 322.990 ;
      LAYER via2 ;
        RECT 24.010 3305.680 24.290 3305.960 ;
        RECT 2623.010 3305.680 2623.290 3305.960 ;
        RECT 13.890 322.520 14.170 322.800 ;
      LAYER met3 ;
        RECT 23.985 3305.970 24.315 3305.985 ;
        RECT 2622.985 3305.970 2623.315 3305.985 ;
        RECT 23.985 3305.670 2623.315 3305.970 ;
        RECT 23.985 3305.655 24.315 3305.670 ;
        RECT 2622.985 3305.655 2623.315 3305.670 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 13.865 322.810 14.195 322.825 ;
        RECT -4.800 322.510 14.195 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 13.865 322.495 14.195 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 110.400 14.650 110.460 ;
        RECT 2690.150 110.400 2690.470 110.460 ;
        RECT 14.330 110.260 2690.470 110.400 ;
        RECT 14.330 110.200 14.650 110.260 ;
        RECT 2690.150 110.200 2690.470 110.260 ;
      LAYER via ;
        RECT 14.360 110.200 14.620 110.460 ;
        RECT 2690.180 110.200 2690.440 110.460 ;
      LAYER met2 ;
        RECT 2686.500 3296.370 2686.780 3300.000 ;
        RECT 2686.500 3296.230 2690.380 3296.370 ;
        RECT 2686.500 3296.000 2686.780 3296.230 ;
        RECT 2690.240 110.490 2690.380 3296.230 ;
        RECT 14.360 110.170 14.620 110.490 ;
        RECT 2690.180 110.170 2690.440 110.490 ;
        RECT 14.420 107.285 14.560 110.170 ;
        RECT 14.350 106.915 14.630 107.285 ;
      LAYER via2 ;
        RECT 14.350 106.960 14.630 107.240 ;
      LAYER met3 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 14.325 107.250 14.655 107.265 ;
        RECT -4.800 106.950 14.655 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 14.325 106.935 14.655 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 539.190 3309.800 539.510 3309.860 ;
        RECT 848.770 3309.800 849.090 3309.860 ;
        RECT 539.190 3309.660 849.090 3309.800 ;
        RECT 539.190 3309.600 539.510 3309.660 ;
        RECT 848.770 3309.600 849.090 3309.660 ;
        RECT 848.770 3301.980 849.090 3302.040 ;
        RECT 2903.590 3301.980 2903.910 3302.040 ;
        RECT 848.770 3301.840 2903.910 3301.980 ;
        RECT 848.770 3301.780 849.090 3301.840 ;
        RECT 2903.590 3301.780 2903.910 3301.840 ;
      LAYER via ;
        RECT 539.220 3309.600 539.480 3309.860 ;
        RECT 848.800 3309.600 849.060 3309.860 ;
        RECT 848.800 3301.780 849.060 3302.040 ;
        RECT 2903.620 3301.780 2903.880 3302.040 ;
      LAYER met2 ;
        RECT 539.220 3309.570 539.480 3309.890 ;
        RECT 848.800 3309.570 849.060 3309.890 ;
        RECT 539.280 3300.000 539.420 3309.570 ;
        RECT 848.860 3302.070 849.000 3309.570 ;
        RECT 848.800 3301.750 849.060 3302.070 ;
        RECT 2903.620 3301.750 2903.880 3302.070 ;
        RECT 539.220 3296.000 539.500 3300.000 ;
        RECT 2903.680 850.525 2903.820 3301.750 ;
        RECT 2903.610 850.155 2903.890 850.525 ;
      LAYER via2 ;
        RECT 2903.610 850.200 2903.890 850.480 ;
      LAYER met3 ;
        RECT 2903.585 850.490 2903.915 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2903.585 850.190 2924.800 850.490 ;
        RECT 2903.585 850.175 2903.915 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 602.210 3308.780 602.530 3308.840 ;
        RECT 793.570 3308.780 793.890 3308.840 ;
        RECT 602.210 3308.640 793.890 3308.780 ;
        RECT 602.210 3308.580 602.530 3308.640 ;
        RECT 793.570 3308.580 793.890 3308.640 ;
        RECT 793.570 3301.640 793.890 3301.700 ;
        RECT 2904.510 3301.640 2904.830 3301.700 ;
        RECT 793.570 3301.500 2904.830 3301.640 ;
        RECT 793.570 3301.440 793.890 3301.500 ;
        RECT 2904.510 3301.440 2904.830 3301.500 ;
      LAYER via ;
        RECT 602.240 3308.580 602.500 3308.840 ;
        RECT 793.600 3308.580 793.860 3308.840 ;
        RECT 793.600 3301.440 793.860 3301.700 ;
        RECT 2904.540 3301.440 2904.800 3301.700 ;
      LAYER met2 ;
        RECT 602.240 3308.550 602.500 3308.870 ;
        RECT 793.600 3308.550 793.860 3308.870 ;
        RECT 602.300 3300.000 602.440 3308.550 ;
        RECT 793.660 3301.730 793.800 3308.550 ;
        RECT 793.600 3301.410 793.860 3301.730 ;
        RECT 2904.540 3301.410 2904.800 3301.730 ;
        RECT 602.240 3296.000 602.520 3300.000 ;
        RECT 2904.600 1085.125 2904.740 3301.410 ;
        RECT 2904.530 1084.755 2904.810 1085.125 ;
      LAYER via2 ;
        RECT 2904.530 1084.800 2904.810 1085.080 ;
      LAYER met3 ;
        RECT 2904.505 1085.090 2904.835 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2904.505 1084.790 2924.800 1085.090 ;
        RECT 2904.505 1084.775 2904.835 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 665.230 3301.300 665.550 3301.360 ;
        RECT 2702.110 3301.300 2702.430 3301.360 ;
        RECT 665.230 3301.160 2702.430 3301.300 ;
        RECT 665.230 3301.100 665.550 3301.160 ;
        RECT 2702.110 3301.100 2702.430 3301.160 ;
        RECT 2702.110 1324.540 2702.430 1324.600 ;
        RECT 2899.910 1324.540 2900.230 1324.600 ;
        RECT 2702.110 1324.400 2900.230 1324.540 ;
        RECT 2702.110 1324.340 2702.430 1324.400 ;
        RECT 2899.910 1324.340 2900.230 1324.400 ;
      LAYER via ;
        RECT 665.260 3301.100 665.520 3301.360 ;
        RECT 2702.140 3301.100 2702.400 3301.360 ;
        RECT 2702.140 1324.340 2702.400 1324.600 ;
        RECT 2899.940 1324.340 2900.200 1324.600 ;
      LAYER met2 ;
        RECT 665.260 3301.070 665.520 3301.390 ;
        RECT 2702.140 3301.070 2702.400 3301.390 ;
        RECT 665.320 3300.000 665.460 3301.070 ;
        RECT 665.260 3296.000 665.540 3300.000 ;
        RECT 2702.200 1324.630 2702.340 3301.070 ;
        RECT 2702.140 1324.310 2702.400 1324.630 ;
        RECT 2899.940 1324.310 2900.200 1324.630 ;
        RECT 2900.000 1319.725 2900.140 1324.310 ;
        RECT 2899.930 1319.355 2900.210 1319.725 ;
      LAYER via2 ;
        RECT 2899.930 1319.400 2900.210 1319.680 ;
      LAYER met3 ;
        RECT 2899.905 1319.690 2900.235 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2899.905 1319.390 2924.800 1319.690 ;
        RECT 2899.905 1319.375 2900.235 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 728.710 3307.420 729.030 3307.480 ;
        RECT 2703.030 3307.420 2703.350 3307.480 ;
        RECT 728.710 3307.280 2703.350 3307.420 ;
        RECT 728.710 3307.220 729.030 3307.280 ;
        RECT 2703.030 3307.220 2703.350 3307.280 ;
        RECT 2703.030 1559.140 2703.350 1559.200 ;
        RECT 2899.910 1559.140 2900.230 1559.200 ;
        RECT 2703.030 1559.000 2900.230 1559.140 ;
        RECT 2703.030 1558.940 2703.350 1559.000 ;
        RECT 2899.910 1558.940 2900.230 1559.000 ;
      LAYER via ;
        RECT 728.740 3307.220 729.000 3307.480 ;
        RECT 2703.060 3307.220 2703.320 3307.480 ;
        RECT 2703.060 1558.940 2703.320 1559.200 ;
        RECT 2899.940 1558.940 2900.200 1559.200 ;
      LAYER met2 ;
        RECT 728.740 3307.190 729.000 3307.510 ;
        RECT 2703.060 3307.190 2703.320 3307.510 ;
        RECT 728.800 3300.000 728.940 3307.190 ;
        RECT 728.740 3296.000 729.020 3300.000 ;
        RECT 2703.120 1559.230 2703.260 3307.190 ;
        RECT 2703.060 1558.910 2703.320 1559.230 ;
        RECT 2899.940 1558.910 2900.200 1559.230 ;
        RECT 2900.000 1554.325 2900.140 1558.910 ;
        RECT 2899.930 1553.955 2900.210 1554.325 ;
      LAYER via2 ;
        RECT 2899.930 1554.000 2900.210 1554.280 ;
      LAYER met3 ;
        RECT 2899.905 1554.290 2900.235 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2899.905 1553.990 2924.800 1554.290 ;
        RECT 2899.905 1553.975 2900.235 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 791.730 3308.100 792.050 3308.160 ;
        RECT 2742.590 3308.100 2742.910 3308.160 ;
        RECT 791.730 3307.960 2742.910 3308.100 ;
        RECT 791.730 3307.900 792.050 3307.960 ;
        RECT 2742.590 3307.900 2742.910 3307.960 ;
        RECT 2742.590 1793.740 2742.910 1793.800 ;
        RECT 2899.910 1793.740 2900.230 1793.800 ;
        RECT 2742.590 1793.600 2900.230 1793.740 ;
        RECT 2742.590 1793.540 2742.910 1793.600 ;
        RECT 2899.910 1793.540 2900.230 1793.600 ;
      LAYER via ;
        RECT 791.760 3307.900 792.020 3308.160 ;
        RECT 2742.620 3307.900 2742.880 3308.160 ;
        RECT 2742.620 1793.540 2742.880 1793.800 ;
        RECT 2899.940 1793.540 2900.200 1793.800 ;
      LAYER met2 ;
        RECT 791.760 3307.870 792.020 3308.190 ;
        RECT 2742.620 3307.870 2742.880 3308.190 ;
        RECT 791.820 3300.000 791.960 3307.870 ;
        RECT 791.760 3296.000 792.040 3300.000 ;
        RECT 2742.680 1793.830 2742.820 3307.870 ;
        RECT 2742.620 1793.510 2742.880 1793.830 ;
        RECT 2899.940 1793.510 2900.200 1793.830 ;
        RECT 2900.000 1789.605 2900.140 1793.510 ;
        RECT 2899.930 1789.235 2900.210 1789.605 ;
      LAYER via2 ;
        RECT 2899.930 1789.280 2900.210 1789.560 ;
      LAYER met3 ;
        RECT 2899.905 1789.570 2900.235 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2899.905 1789.270 2924.800 1789.570 ;
        RECT 2899.905 1789.255 2900.235 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 854.750 3309.460 855.070 3309.520 ;
        RECT 2708.090 3309.460 2708.410 3309.520 ;
        RECT 854.750 3309.320 2708.410 3309.460 ;
        RECT 854.750 3309.260 855.070 3309.320 ;
        RECT 2708.090 3309.260 2708.410 3309.320 ;
        RECT 2708.090 2028.340 2708.410 2028.400 ;
        RECT 2899.910 2028.340 2900.230 2028.400 ;
        RECT 2708.090 2028.200 2900.230 2028.340 ;
        RECT 2708.090 2028.140 2708.410 2028.200 ;
        RECT 2899.910 2028.140 2900.230 2028.200 ;
      LAYER via ;
        RECT 854.780 3309.260 855.040 3309.520 ;
        RECT 2708.120 3309.260 2708.380 3309.520 ;
        RECT 2708.120 2028.140 2708.380 2028.400 ;
        RECT 2899.940 2028.140 2900.200 2028.400 ;
      LAYER met2 ;
        RECT 854.780 3309.230 855.040 3309.550 ;
        RECT 2708.120 3309.230 2708.380 3309.550 ;
        RECT 854.840 3300.000 854.980 3309.230 ;
        RECT 854.780 3296.000 855.060 3300.000 ;
        RECT 2708.180 2028.430 2708.320 3309.230 ;
        RECT 2708.120 2028.110 2708.380 2028.430 ;
        RECT 2899.940 2028.110 2900.200 2028.430 ;
        RECT 2900.000 2024.205 2900.140 2028.110 ;
        RECT 2899.930 2023.835 2900.210 2024.205 ;
      LAYER via2 ;
        RECT 2899.930 2023.880 2900.210 2024.160 ;
      LAYER met3 ;
        RECT 2899.905 2024.170 2900.235 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2899.905 2023.870 2924.800 2024.170 ;
        RECT 2899.905 2023.855 2900.235 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 918.230 3309.800 918.550 3309.860 ;
        RECT 2708.550 3309.800 2708.870 3309.860 ;
        RECT 918.230 3309.660 2708.870 3309.800 ;
        RECT 918.230 3309.600 918.550 3309.660 ;
        RECT 2708.550 3309.600 2708.870 3309.660 ;
        RECT 2708.550 2262.940 2708.870 2263.000 ;
        RECT 2899.910 2262.940 2900.230 2263.000 ;
        RECT 2708.550 2262.800 2900.230 2262.940 ;
        RECT 2708.550 2262.740 2708.870 2262.800 ;
        RECT 2899.910 2262.740 2900.230 2262.800 ;
      LAYER via ;
        RECT 918.260 3309.600 918.520 3309.860 ;
        RECT 2708.580 3309.600 2708.840 3309.860 ;
        RECT 2708.580 2262.740 2708.840 2263.000 ;
        RECT 2899.940 2262.740 2900.200 2263.000 ;
      LAYER met2 ;
        RECT 918.260 3309.570 918.520 3309.890 ;
        RECT 2708.580 3309.570 2708.840 3309.890 ;
        RECT 918.320 3300.000 918.460 3309.570 ;
        RECT 918.260 3296.000 918.540 3300.000 ;
        RECT 2708.640 2263.030 2708.780 3309.570 ;
        RECT 2708.580 2262.710 2708.840 2263.030 ;
        RECT 2899.940 2262.710 2900.200 2263.030 ;
        RECT 2900.000 2258.805 2900.140 2262.710 ;
        RECT 2899.930 2258.435 2900.210 2258.805 ;
      LAYER via2 ;
        RECT 2899.930 2258.480 2900.210 2258.760 ;
      LAYER met3 ;
        RECT 2899.905 2258.770 2900.235 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2899.905 2258.470 2924.800 2258.770 ;
        RECT 2899.905 2258.455 2900.235 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 633.030 17.580 633.350 17.640 ;
        RECT 814.730 17.580 815.050 17.640 ;
        RECT 633.030 17.440 815.050 17.580 ;
        RECT 633.030 17.380 633.350 17.440 ;
        RECT 814.730 17.380 815.050 17.440 ;
      LAYER via ;
        RECT 633.060 17.380 633.320 17.640 ;
        RECT 814.760 17.380 815.020 17.640 ;
      LAYER met2 ;
        RECT 818.900 300.290 819.180 304.000 ;
        RECT 814.820 300.150 819.180 300.290 ;
        RECT 814.820 17.670 814.960 300.150 ;
        RECT 818.900 300.000 819.180 300.150 ;
        RECT 633.060 17.350 633.320 17.670 ;
        RECT 814.760 17.350 815.020 17.670 ;
        RECT 633.120 2.400 633.260 17.350 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2288.110 286.860 2288.430 286.920 ;
        RECT 2415.530 286.860 2415.850 286.920 ;
        RECT 2288.110 286.720 2415.850 286.860 ;
        RECT 2288.110 286.660 2288.430 286.720 ;
        RECT 2415.530 286.660 2415.850 286.720 ;
      LAYER via ;
        RECT 2288.140 286.660 2288.400 286.920 ;
        RECT 2415.560 286.660 2415.820 286.920 ;
      LAYER met2 ;
        RECT 2288.140 300.000 2288.420 304.000 ;
        RECT 2288.200 286.950 2288.340 300.000 ;
        RECT 2288.140 286.630 2288.400 286.950 ;
        RECT 2415.560 286.630 2415.820 286.950 ;
        RECT 2415.620 3.130 2415.760 286.630 ;
        RECT 2415.620 2.990 2417.600 3.130 ;
        RECT 2417.460 2.400 2417.600 2.990 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2302.830 289.580 2303.150 289.640 ;
        RECT 2429.790 289.580 2430.110 289.640 ;
        RECT 2302.830 289.440 2430.110 289.580 ;
        RECT 2302.830 289.380 2303.150 289.440 ;
        RECT 2429.790 289.380 2430.110 289.440 ;
        RECT 2429.790 2.960 2430.110 3.020 ;
        RECT 2434.850 2.960 2435.170 3.020 ;
        RECT 2429.790 2.820 2435.170 2.960 ;
        RECT 2429.790 2.760 2430.110 2.820 ;
        RECT 2434.850 2.760 2435.170 2.820 ;
      LAYER via ;
        RECT 2302.860 289.380 2303.120 289.640 ;
        RECT 2429.820 289.380 2430.080 289.640 ;
        RECT 2429.820 2.760 2430.080 3.020 ;
        RECT 2434.880 2.760 2435.140 3.020 ;
      LAYER met2 ;
        RECT 2302.860 300.000 2303.140 304.000 ;
        RECT 2302.920 289.670 2303.060 300.000 ;
        RECT 2302.860 289.350 2303.120 289.670 ;
        RECT 2429.820 289.350 2430.080 289.670 ;
        RECT 2429.880 3.050 2430.020 289.350 ;
        RECT 2429.820 2.730 2430.080 3.050 ;
        RECT 2434.880 2.730 2435.140 3.050 ;
        RECT 2434.940 2.400 2435.080 2.730 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2317.550 286.520 2317.870 286.580 ;
        RECT 2450.490 286.520 2450.810 286.580 ;
        RECT 2317.550 286.380 2450.810 286.520 ;
        RECT 2317.550 286.320 2317.870 286.380 ;
        RECT 2450.490 286.320 2450.810 286.380 ;
      LAYER via ;
        RECT 2317.580 286.320 2317.840 286.580 ;
        RECT 2450.520 286.320 2450.780 286.580 ;
      LAYER met2 ;
        RECT 2317.580 300.000 2317.860 304.000 ;
        RECT 2317.640 286.610 2317.780 300.000 ;
        RECT 2317.580 286.290 2317.840 286.610 ;
        RECT 2450.520 286.290 2450.780 286.610 ;
        RECT 2450.580 16.730 2450.720 286.290 ;
        RECT 2450.580 16.590 2453.020 16.730 ;
        RECT 2452.880 2.400 2453.020 16.590 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2332.270 288.560 2332.590 288.620 ;
        RECT 2471.190 288.560 2471.510 288.620 ;
        RECT 2332.270 288.420 2471.510 288.560 ;
        RECT 2332.270 288.360 2332.590 288.420 ;
        RECT 2471.190 288.360 2471.510 288.420 ;
      LAYER via ;
        RECT 2332.300 288.360 2332.560 288.620 ;
        RECT 2471.220 288.360 2471.480 288.620 ;
      LAYER met2 ;
        RECT 2332.300 300.000 2332.580 304.000 ;
        RECT 2332.360 288.650 2332.500 300.000 ;
        RECT 2332.300 288.330 2332.560 288.650 ;
        RECT 2471.220 288.330 2471.480 288.650 ;
        RECT 2471.280 17.410 2471.420 288.330 ;
        RECT 2470.820 17.270 2471.420 17.410 ;
        RECT 2470.820 2.400 2470.960 17.270 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2484.530 288.560 2484.850 288.620 ;
        RECT 2471.740 288.420 2484.850 288.560 ;
        RECT 2346.990 288.220 2347.310 288.280 ;
        RECT 2471.740 288.220 2471.880 288.420 ;
        RECT 2484.530 288.360 2484.850 288.420 ;
        RECT 2346.990 288.080 2471.880 288.220 ;
        RECT 2346.990 288.020 2347.310 288.080 ;
      LAYER via ;
        RECT 2347.020 288.020 2347.280 288.280 ;
        RECT 2484.560 288.360 2484.820 288.620 ;
      LAYER met2 ;
        RECT 2347.020 300.000 2347.300 304.000 ;
        RECT 2347.080 288.310 2347.220 300.000 ;
        RECT 2484.560 288.330 2484.820 288.650 ;
        RECT 2347.020 287.990 2347.280 288.310 ;
        RECT 2484.620 16.730 2484.760 288.330 ;
        RECT 2484.620 16.590 2488.900 16.730 ;
        RECT 2488.760 2.400 2488.900 16.590 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2361.710 287.200 2362.030 287.260 ;
        RECT 2505.230 287.200 2505.550 287.260 ;
        RECT 2361.710 287.060 2505.550 287.200 ;
        RECT 2361.710 287.000 2362.030 287.060 ;
        RECT 2505.230 287.000 2505.550 287.060 ;
        RECT 2505.230 2.960 2505.550 3.020 ;
        RECT 2506.150 2.960 2506.470 3.020 ;
        RECT 2505.230 2.820 2506.470 2.960 ;
        RECT 2505.230 2.760 2505.550 2.820 ;
        RECT 2506.150 2.760 2506.470 2.820 ;
      LAYER via ;
        RECT 2361.740 287.000 2362.000 287.260 ;
        RECT 2505.260 287.000 2505.520 287.260 ;
        RECT 2505.260 2.760 2505.520 3.020 ;
        RECT 2506.180 2.760 2506.440 3.020 ;
      LAYER met2 ;
        RECT 2361.740 300.000 2362.020 304.000 ;
        RECT 2361.800 287.290 2361.940 300.000 ;
        RECT 2361.740 286.970 2362.000 287.290 ;
        RECT 2505.260 286.970 2505.520 287.290 ;
        RECT 2505.320 3.050 2505.460 286.970 ;
        RECT 2505.260 2.730 2505.520 3.050 ;
        RECT 2506.180 2.730 2506.440 3.050 ;
        RECT 2506.240 2.400 2506.380 2.730 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2376.430 287.880 2376.750 287.940 ;
        RECT 2518.570 287.880 2518.890 287.940 ;
        RECT 2376.430 287.740 2518.890 287.880 ;
        RECT 2376.430 287.680 2376.750 287.740 ;
        RECT 2518.570 287.680 2518.890 287.740 ;
        RECT 2518.570 2.960 2518.890 3.020 ;
        RECT 2524.090 2.960 2524.410 3.020 ;
        RECT 2518.570 2.820 2524.410 2.960 ;
        RECT 2518.570 2.760 2518.890 2.820 ;
        RECT 2524.090 2.760 2524.410 2.820 ;
      LAYER via ;
        RECT 2376.460 287.680 2376.720 287.940 ;
        RECT 2518.600 287.680 2518.860 287.940 ;
        RECT 2518.600 2.760 2518.860 3.020 ;
        RECT 2524.120 2.760 2524.380 3.020 ;
      LAYER met2 ;
        RECT 2376.460 300.000 2376.740 304.000 ;
        RECT 2376.520 287.970 2376.660 300.000 ;
        RECT 2376.460 287.650 2376.720 287.970 ;
        RECT 2518.600 287.650 2518.860 287.970 ;
        RECT 2518.660 3.050 2518.800 287.650 ;
        RECT 2518.600 2.730 2518.860 3.050 ;
        RECT 2524.120 2.730 2524.380 3.050 ;
        RECT 2524.180 2.400 2524.320 2.730 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2391.150 287.540 2391.470 287.600 ;
        RECT 2539.730 287.540 2540.050 287.600 ;
        RECT 2391.150 287.400 2540.050 287.540 ;
        RECT 2391.150 287.340 2391.470 287.400 ;
        RECT 2539.730 287.340 2540.050 287.400 ;
        RECT 2539.730 2.960 2540.050 3.020 ;
        RECT 2542.030 2.960 2542.350 3.020 ;
        RECT 2539.730 2.820 2542.350 2.960 ;
        RECT 2539.730 2.760 2540.050 2.820 ;
        RECT 2542.030 2.760 2542.350 2.820 ;
      LAYER via ;
        RECT 2391.180 287.340 2391.440 287.600 ;
        RECT 2539.760 287.340 2540.020 287.600 ;
        RECT 2539.760 2.760 2540.020 3.020 ;
        RECT 2542.060 2.760 2542.320 3.020 ;
      LAYER met2 ;
        RECT 2391.180 300.000 2391.460 304.000 ;
        RECT 2391.240 287.630 2391.380 300.000 ;
        RECT 2391.180 287.310 2391.440 287.630 ;
        RECT 2539.760 287.310 2540.020 287.630 ;
        RECT 2539.820 3.050 2539.960 287.310 ;
        RECT 2539.760 2.730 2540.020 3.050 ;
        RECT 2542.060 2.730 2542.320 3.050 ;
        RECT 2542.120 2.400 2542.260 2.730 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2405.870 286.180 2406.190 286.240 ;
        RECT 2560.430 286.180 2560.750 286.240 ;
        RECT 2405.870 286.040 2560.750 286.180 ;
        RECT 2405.870 285.980 2406.190 286.040 ;
        RECT 2560.430 285.980 2560.750 286.040 ;
      LAYER via ;
        RECT 2405.900 285.980 2406.160 286.240 ;
        RECT 2560.460 285.980 2560.720 286.240 ;
      LAYER met2 ;
        RECT 2405.900 300.000 2406.180 304.000 ;
        RECT 2405.960 286.270 2406.100 300.000 ;
        RECT 2405.900 285.950 2406.160 286.270 ;
        RECT 2560.460 285.950 2560.720 286.270 ;
        RECT 2560.520 3.130 2560.660 285.950 ;
        RECT 2560.060 2.990 2560.660 3.130 ;
        RECT 2560.060 2.400 2560.200 2.990 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2420.590 286.860 2420.910 286.920 ;
        RECT 2573.770 286.860 2574.090 286.920 ;
        RECT 2420.590 286.720 2574.090 286.860 ;
        RECT 2420.590 286.660 2420.910 286.720 ;
        RECT 2573.770 286.660 2574.090 286.720 ;
        RECT 2573.770 2.960 2574.090 3.020 ;
        RECT 2577.910 2.960 2578.230 3.020 ;
        RECT 2573.770 2.820 2578.230 2.960 ;
        RECT 2573.770 2.760 2574.090 2.820 ;
        RECT 2577.910 2.760 2578.230 2.820 ;
      LAYER via ;
        RECT 2420.620 286.660 2420.880 286.920 ;
        RECT 2573.800 286.660 2574.060 286.920 ;
        RECT 2573.800 2.760 2574.060 3.020 ;
        RECT 2577.940 2.760 2578.200 3.020 ;
      LAYER met2 ;
        RECT 2420.620 300.000 2420.900 304.000 ;
        RECT 2420.680 286.950 2420.820 300.000 ;
        RECT 2420.620 286.630 2420.880 286.950 ;
        RECT 2573.800 286.630 2574.060 286.950 ;
        RECT 2573.860 3.050 2574.000 286.630 ;
        RECT 2573.800 2.730 2574.060 3.050 ;
        RECT 2577.940 2.730 2578.200 3.050 ;
        RECT 2578.000 2.400 2578.140 2.730 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 960.165 144.925 960.335 193.035 ;
        RECT 961.085 48.365 961.255 96.475 ;
      LAYER mcon ;
        RECT 960.165 192.865 960.335 193.035 ;
        RECT 961.085 96.305 961.255 96.475 ;
      LAYER met1 ;
        RECT 960.105 193.020 960.395 193.065 ;
        RECT 960.550 193.020 960.870 193.080 ;
        RECT 960.105 192.880 960.870 193.020 ;
        RECT 960.105 192.835 960.395 192.880 ;
        RECT 960.550 192.820 960.870 192.880 ;
        RECT 960.090 145.080 960.410 145.140 ;
        RECT 959.895 144.940 960.410 145.080 ;
        RECT 960.090 144.880 960.410 144.940 ;
        RECT 961.010 96.460 961.330 96.520 ;
        RECT 960.815 96.320 961.330 96.460 ;
        RECT 961.010 96.260 961.330 96.320 ;
        RECT 961.025 48.520 961.315 48.565 ;
        RECT 961.470 48.520 961.790 48.580 ;
        RECT 961.025 48.380 961.790 48.520 ;
        RECT 961.025 48.335 961.315 48.380 ;
        RECT 961.470 48.320 961.790 48.380 ;
        RECT 811.510 17.240 811.830 17.300 ;
        RECT 961.470 17.240 961.790 17.300 ;
        RECT 811.510 17.100 961.790 17.240 ;
        RECT 811.510 17.040 811.830 17.100 ;
        RECT 961.470 17.040 961.790 17.100 ;
      LAYER via ;
        RECT 960.580 192.820 960.840 193.080 ;
        RECT 960.120 144.880 960.380 145.140 ;
        RECT 961.040 96.260 961.300 96.520 ;
        RECT 961.500 48.320 961.760 48.580 ;
        RECT 811.540 17.040 811.800 17.300 ;
        RECT 961.500 17.040 961.760 17.300 ;
      LAYER met2 ;
        RECT 965.640 300.970 965.920 304.000 ;
        RECT 961.560 300.830 965.920 300.970 ;
        RECT 961.560 277.850 961.700 300.830 ;
        RECT 965.640 300.000 965.920 300.830 ;
        RECT 960.640 277.710 961.700 277.850 ;
        RECT 960.640 193.110 960.780 277.710 ;
        RECT 960.580 192.790 960.840 193.110 ;
        RECT 960.120 144.850 960.380 145.170 ;
        RECT 960.180 110.570 960.320 144.850 ;
        RECT 960.180 110.430 961.240 110.570 ;
        RECT 961.100 96.550 961.240 110.430 ;
        RECT 961.040 96.230 961.300 96.550 ;
        RECT 961.500 48.290 961.760 48.610 ;
        RECT 961.560 17.330 961.700 48.290 ;
        RECT 811.540 17.010 811.800 17.330 ;
        RECT 961.500 17.010 961.760 17.330 ;
        RECT 811.600 2.400 811.740 17.010 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2435.310 24.040 2435.630 24.100 ;
        RECT 2595.390 24.040 2595.710 24.100 ;
        RECT 2435.310 23.900 2595.710 24.040 ;
        RECT 2435.310 23.840 2435.630 23.900 ;
        RECT 2595.390 23.840 2595.710 23.900 ;
      LAYER via ;
        RECT 2435.340 23.840 2435.600 24.100 ;
        RECT 2595.420 23.840 2595.680 24.100 ;
      LAYER met2 ;
        RECT 2435.340 300.000 2435.620 304.000 ;
        RECT 2435.400 24.130 2435.540 300.000 ;
        RECT 2435.340 23.810 2435.600 24.130 ;
        RECT 2595.420 23.810 2595.680 24.130 ;
        RECT 2595.480 2.400 2595.620 23.810 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2450.030 285.500 2450.350 285.560 ;
        RECT 2608.270 285.500 2608.590 285.560 ;
        RECT 2450.030 285.360 2608.590 285.500 ;
        RECT 2450.030 285.300 2450.350 285.360 ;
        RECT 2608.270 285.300 2608.590 285.360 ;
        RECT 2608.270 2.960 2608.590 3.020 ;
        RECT 2613.330 2.960 2613.650 3.020 ;
        RECT 2608.270 2.820 2613.650 2.960 ;
        RECT 2608.270 2.760 2608.590 2.820 ;
        RECT 2613.330 2.760 2613.650 2.820 ;
      LAYER via ;
        RECT 2450.060 285.300 2450.320 285.560 ;
        RECT 2608.300 285.300 2608.560 285.560 ;
        RECT 2608.300 2.760 2608.560 3.020 ;
        RECT 2613.360 2.760 2613.620 3.020 ;
      LAYER met2 ;
        RECT 2450.060 300.000 2450.340 304.000 ;
        RECT 2450.120 285.590 2450.260 300.000 ;
        RECT 2450.060 285.270 2450.320 285.590 ;
        RECT 2608.300 285.270 2608.560 285.590 ;
        RECT 2608.360 3.050 2608.500 285.270 ;
        RECT 2608.300 2.730 2608.560 3.050 ;
        RECT 2613.360 2.730 2613.620 3.050 ;
        RECT 2613.420 2.400 2613.560 2.730 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2464.290 286.520 2464.610 286.580 ;
        RECT 2628.970 286.520 2629.290 286.580 ;
        RECT 2464.290 286.380 2629.290 286.520 ;
        RECT 2464.290 286.320 2464.610 286.380 ;
        RECT 2628.970 286.320 2629.290 286.380 ;
        RECT 2628.970 2.960 2629.290 3.020 ;
        RECT 2631.270 2.960 2631.590 3.020 ;
        RECT 2628.970 2.820 2631.590 2.960 ;
        RECT 2628.970 2.760 2629.290 2.820 ;
        RECT 2631.270 2.760 2631.590 2.820 ;
      LAYER via ;
        RECT 2464.320 286.320 2464.580 286.580 ;
        RECT 2629.000 286.320 2629.260 286.580 ;
        RECT 2629.000 2.760 2629.260 3.020 ;
        RECT 2631.300 2.760 2631.560 3.020 ;
      LAYER met2 ;
        RECT 2464.320 300.000 2464.600 304.000 ;
        RECT 2464.380 286.610 2464.520 300.000 ;
        RECT 2464.320 286.290 2464.580 286.610 ;
        RECT 2629.000 286.290 2629.260 286.610 ;
        RECT 2629.060 3.050 2629.200 286.290 ;
        RECT 2629.000 2.730 2629.260 3.050 ;
        RECT 2631.300 2.730 2631.560 3.050 ;
        RECT 2631.360 2.400 2631.500 2.730 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2479.010 285.160 2479.330 285.220 ;
        RECT 2643.690 285.160 2644.010 285.220 ;
        RECT 2479.010 285.020 2644.010 285.160 ;
        RECT 2479.010 284.960 2479.330 285.020 ;
        RECT 2643.690 284.960 2644.010 285.020 ;
      LAYER via ;
        RECT 2479.040 284.960 2479.300 285.220 ;
        RECT 2643.720 284.960 2643.980 285.220 ;
      LAYER met2 ;
        RECT 2479.040 300.000 2479.320 304.000 ;
        RECT 2479.100 285.250 2479.240 300.000 ;
        RECT 2479.040 284.930 2479.300 285.250 ;
        RECT 2643.720 284.930 2643.980 285.250 ;
        RECT 2643.780 16.730 2643.920 284.930 ;
        RECT 2643.780 16.590 2649.440 16.730 ;
        RECT 2649.300 2.400 2649.440 16.590 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2663.470 289.240 2663.790 289.300 ;
        RECT 2650.220 289.100 2663.790 289.240 ;
        RECT 2493.730 288.900 2494.050 288.960 ;
        RECT 2650.220 288.900 2650.360 289.100 ;
        RECT 2663.470 289.040 2663.790 289.100 ;
        RECT 2493.730 288.760 2650.360 288.900 ;
        RECT 2493.730 288.700 2494.050 288.760 ;
      LAYER via ;
        RECT 2493.760 288.700 2494.020 288.960 ;
        RECT 2663.500 289.040 2663.760 289.300 ;
      LAYER met2 ;
        RECT 2493.760 300.000 2494.040 304.000 ;
        RECT 2493.820 288.990 2493.960 300.000 ;
        RECT 2663.500 289.010 2663.760 289.330 ;
        RECT 2493.760 288.670 2494.020 288.990 ;
        RECT 2663.560 14.010 2663.700 289.010 ;
        RECT 2663.560 13.870 2667.380 14.010 ;
        RECT 2667.240 2.400 2667.380 13.870 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2511.210 26.080 2511.530 26.140 ;
        RECT 2684.630 26.080 2684.950 26.140 ;
        RECT 2511.210 25.940 2684.950 26.080 ;
        RECT 2511.210 25.880 2511.530 25.940 ;
        RECT 2684.630 25.880 2684.950 25.940 ;
      LAYER via ;
        RECT 2511.240 25.880 2511.500 26.140 ;
        RECT 2684.660 25.880 2684.920 26.140 ;
      LAYER met2 ;
        RECT 2508.480 300.290 2508.760 304.000 ;
        RECT 2508.480 300.150 2511.440 300.290 ;
        RECT 2508.480 300.000 2508.760 300.150 ;
        RECT 2511.300 26.170 2511.440 300.150 ;
        RECT 2511.240 25.850 2511.500 26.170 ;
        RECT 2684.660 25.850 2684.920 26.170 ;
        RECT 2684.720 2.400 2684.860 25.850 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2525.010 25.740 2525.330 25.800 ;
        RECT 2702.570 25.740 2702.890 25.800 ;
        RECT 2525.010 25.600 2702.890 25.740 ;
        RECT 2525.010 25.540 2525.330 25.600 ;
        RECT 2702.570 25.540 2702.890 25.600 ;
      LAYER via ;
        RECT 2525.040 25.540 2525.300 25.800 ;
        RECT 2702.600 25.540 2702.860 25.800 ;
      LAYER met2 ;
        RECT 2523.200 300.290 2523.480 304.000 ;
        RECT 2523.200 300.150 2525.240 300.290 ;
        RECT 2523.200 300.000 2523.480 300.150 ;
        RECT 2525.100 25.830 2525.240 300.150 ;
        RECT 2525.040 25.510 2525.300 25.830 ;
        RECT 2702.600 25.510 2702.860 25.830 ;
        RECT 2702.660 2.400 2702.800 25.510 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2537.890 287.200 2538.210 287.260 ;
        RECT 2718.670 287.200 2718.990 287.260 ;
        RECT 2537.890 287.060 2718.990 287.200 ;
        RECT 2537.890 287.000 2538.210 287.060 ;
        RECT 2718.670 287.000 2718.990 287.060 ;
        RECT 2718.670 2.960 2718.990 3.020 ;
        RECT 2720.510 2.960 2720.830 3.020 ;
        RECT 2718.670 2.820 2720.830 2.960 ;
        RECT 2718.670 2.760 2718.990 2.820 ;
        RECT 2720.510 2.760 2720.830 2.820 ;
      LAYER via ;
        RECT 2537.920 287.000 2538.180 287.260 ;
        RECT 2718.700 287.000 2718.960 287.260 ;
        RECT 2718.700 2.760 2718.960 3.020 ;
        RECT 2720.540 2.760 2720.800 3.020 ;
      LAYER met2 ;
        RECT 2537.920 300.000 2538.200 304.000 ;
        RECT 2537.980 287.290 2538.120 300.000 ;
        RECT 2537.920 286.970 2538.180 287.290 ;
        RECT 2718.700 286.970 2718.960 287.290 ;
        RECT 2718.760 3.050 2718.900 286.970 ;
        RECT 2718.700 2.730 2718.960 3.050 ;
        RECT 2720.540 2.730 2720.800 3.050 ;
        RECT 2720.600 2.400 2720.740 2.730 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2552.610 25.400 2552.930 25.460 ;
        RECT 2738.450 25.400 2738.770 25.460 ;
        RECT 2552.610 25.260 2738.770 25.400 ;
        RECT 2552.610 25.200 2552.930 25.260 ;
        RECT 2738.450 25.200 2738.770 25.260 ;
      LAYER via ;
        RECT 2552.640 25.200 2552.900 25.460 ;
        RECT 2738.480 25.200 2738.740 25.460 ;
      LAYER met2 ;
        RECT 2552.640 300.000 2552.920 304.000 ;
        RECT 2552.700 25.490 2552.840 300.000 ;
        RECT 2552.640 25.170 2552.900 25.490 ;
        RECT 2738.480 25.170 2738.740 25.490 ;
        RECT 2738.540 2.400 2738.680 25.170 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2567.330 288.220 2567.650 288.280 ;
        RECT 2572.850 288.220 2573.170 288.280 ;
        RECT 2567.330 288.080 2573.170 288.220 ;
        RECT 2567.330 288.020 2567.650 288.080 ;
        RECT 2572.850 288.020 2573.170 288.080 ;
        RECT 2572.850 25.060 2573.170 25.120 ;
        RECT 2755.930 25.060 2756.250 25.120 ;
        RECT 2572.850 24.920 2756.250 25.060 ;
        RECT 2572.850 24.860 2573.170 24.920 ;
        RECT 2755.930 24.860 2756.250 24.920 ;
      LAYER via ;
        RECT 2567.360 288.020 2567.620 288.280 ;
        RECT 2572.880 288.020 2573.140 288.280 ;
        RECT 2572.880 24.860 2573.140 25.120 ;
        RECT 2755.960 24.860 2756.220 25.120 ;
      LAYER met2 ;
        RECT 2567.360 300.000 2567.640 304.000 ;
        RECT 2567.420 288.310 2567.560 300.000 ;
        RECT 2567.360 287.990 2567.620 288.310 ;
        RECT 2572.880 287.990 2573.140 288.310 ;
        RECT 2572.940 25.150 2573.080 287.990 ;
        RECT 2572.880 24.830 2573.140 25.150 ;
        RECT 2755.960 24.830 2756.220 25.150 ;
        RECT 2756.020 2.400 2756.160 24.830 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 980.330 17.920 980.650 17.980 ;
        RECT 956.040 17.780 980.650 17.920 ;
        RECT 829.450 17.580 829.770 17.640 ;
        RECT 956.040 17.580 956.180 17.780 ;
        RECT 980.330 17.720 980.650 17.780 ;
        RECT 829.450 17.440 956.180 17.580 ;
        RECT 829.450 17.380 829.770 17.440 ;
      LAYER via ;
        RECT 829.480 17.380 829.740 17.640 ;
        RECT 980.360 17.720 980.620 17.980 ;
      LAYER met2 ;
        RECT 980.360 300.000 980.640 304.000 ;
        RECT 980.420 18.010 980.560 300.000 ;
        RECT 980.360 17.690 980.620 18.010 ;
        RECT 829.480 17.350 829.740 17.670 ;
        RECT 829.540 2.400 829.680 17.350 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2582.050 286.860 2582.370 286.920 ;
        RECT 2774.330 286.860 2774.650 286.920 ;
        RECT 2582.050 286.720 2774.650 286.860 ;
        RECT 2582.050 286.660 2582.370 286.720 ;
        RECT 2774.330 286.660 2774.650 286.720 ;
      LAYER via ;
        RECT 2582.080 286.660 2582.340 286.920 ;
        RECT 2774.360 286.660 2774.620 286.920 ;
      LAYER met2 ;
        RECT 2582.080 300.000 2582.360 304.000 ;
        RECT 2582.140 286.950 2582.280 300.000 ;
        RECT 2582.080 286.630 2582.340 286.950 ;
        RECT 2774.360 286.630 2774.620 286.950 ;
        RECT 2774.420 17.410 2774.560 286.630 ;
        RECT 2773.960 17.270 2774.560 17.410 ;
        RECT 2773.960 2.400 2774.100 17.270 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2596.770 289.240 2597.090 289.300 ;
        RECT 2600.910 289.240 2601.230 289.300 ;
        RECT 2596.770 289.100 2601.230 289.240 ;
        RECT 2596.770 289.040 2597.090 289.100 ;
        RECT 2600.910 289.040 2601.230 289.100 ;
        RECT 2600.910 24.720 2601.230 24.780 ;
        RECT 2791.810 24.720 2792.130 24.780 ;
        RECT 2600.910 24.580 2792.130 24.720 ;
        RECT 2600.910 24.520 2601.230 24.580 ;
        RECT 2791.810 24.520 2792.130 24.580 ;
      LAYER via ;
        RECT 2596.800 289.040 2597.060 289.300 ;
        RECT 2600.940 289.040 2601.200 289.300 ;
        RECT 2600.940 24.520 2601.200 24.780 ;
        RECT 2791.840 24.520 2792.100 24.780 ;
      LAYER met2 ;
        RECT 2596.800 300.000 2597.080 304.000 ;
        RECT 2596.860 289.330 2597.000 300.000 ;
        RECT 2596.800 289.010 2597.060 289.330 ;
        RECT 2600.940 289.010 2601.200 289.330 ;
        RECT 2601.000 24.810 2601.140 289.010 ;
        RECT 2600.940 24.490 2601.200 24.810 ;
        RECT 2791.840 24.490 2792.100 24.810 ;
        RECT 2791.900 2.400 2792.040 24.490 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2614.710 24.380 2615.030 24.440 ;
        RECT 2809.750 24.380 2810.070 24.440 ;
        RECT 2614.710 24.240 2810.070 24.380 ;
        RECT 2614.710 24.180 2615.030 24.240 ;
        RECT 2809.750 24.180 2810.070 24.240 ;
      LAYER via ;
        RECT 2614.740 24.180 2615.000 24.440 ;
        RECT 2809.780 24.180 2810.040 24.440 ;
      LAYER met2 ;
        RECT 2611.520 300.290 2611.800 304.000 ;
        RECT 2611.520 300.150 2614.940 300.290 ;
        RECT 2611.520 300.000 2611.800 300.150 ;
        RECT 2614.800 24.470 2614.940 300.150 ;
        RECT 2614.740 24.150 2615.000 24.470 ;
        RECT 2809.780 24.150 2810.040 24.470 ;
        RECT 2809.840 2.400 2809.980 24.150 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2626.210 286.180 2626.530 286.240 ;
        RECT 2822.170 286.180 2822.490 286.240 ;
        RECT 2626.210 286.040 2822.490 286.180 ;
        RECT 2626.210 285.980 2626.530 286.040 ;
        RECT 2822.170 285.980 2822.490 286.040 ;
      LAYER via ;
        RECT 2626.240 285.980 2626.500 286.240 ;
        RECT 2822.200 285.980 2822.460 286.240 ;
      LAYER met2 ;
        RECT 2626.240 300.000 2626.520 304.000 ;
        RECT 2626.300 286.270 2626.440 300.000 ;
        RECT 2626.240 285.950 2626.500 286.270 ;
        RECT 2822.200 285.950 2822.460 286.270 ;
        RECT 2822.260 17.410 2822.400 285.950 ;
        RECT 2822.260 17.270 2827.920 17.410 ;
        RECT 2827.780 2.400 2827.920 17.270 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2640.930 286.520 2641.250 286.580 ;
        RECT 2832.290 286.520 2832.610 286.580 ;
        RECT 2640.930 286.380 2832.610 286.520 ;
        RECT 2640.930 286.320 2641.250 286.380 ;
        RECT 2832.290 286.320 2832.610 286.380 ;
        RECT 2832.290 20.640 2832.610 20.700 ;
        RECT 2845.170 20.640 2845.490 20.700 ;
        RECT 2832.290 20.500 2845.490 20.640 ;
        RECT 2832.290 20.440 2832.610 20.500 ;
        RECT 2845.170 20.440 2845.490 20.500 ;
      LAYER via ;
        RECT 2640.960 286.320 2641.220 286.580 ;
        RECT 2832.320 286.320 2832.580 286.580 ;
        RECT 2832.320 20.440 2832.580 20.700 ;
        RECT 2845.200 20.440 2845.460 20.700 ;
      LAYER met2 ;
        RECT 2640.960 300.000 2641.240 304.000 ;
        RECT 2641.020 286.610 2641.160 300.000 ;
        RECT 2640.960 286.290 2641.220 286.610 ;
        RECT 2832.320 286.290 2832.580 286.610 ;
        RECT 2832.380 20.730 2832.520 286.290 ;
        RECT 2832.320 20.410 2832.580 20.730 ;
        RECT 2845.200 20.410 2845.460 20.730 ;
        RECT 2845.260 2.400 2845.400 20.410 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2655.650 24.040 2655.970 24.100 ;
        RECT 2863.110 24.040 2863.430 24.100 ;
        RECT 2655.650 23.900 2863.430 24.040 ;
        RECT 2655.650 23.840 2655.970 23.900 ;
        RECT 2863.110 23.840 2863.430 23.900 ;
      LAYER via ;
        RECT 2655.680 23.840 2655.940 24.100 ;
        RECT 2863.140 23.840 2863.400 24.100 ;
      LAYER met2 ;
        RECT 2655.680 300.000 2655.960 304.000 ;
        RECT 2655.740 24.130 2655.880 300.000 ;
        RECT 2655.680 23.810 2655.940 24.130 ;
        RECT 2863.140 23.810 2863.400 24.130 ;
        RECT 2863.200 2.400 2863.340 23.810 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2670.370 288.900 2670.690 288.960 ;
        RECT 2676.810 288.900 2677.130 288.960 ;
        RECT 2670.370 288.760 2677.130 288.900 ;
        RECT 2670.370 288.700 2670.690 288.760 ;
        RECT 2676.810 288.700 2677.130 288.760 ;
        RECT 2676.810 17.920 2677.130 17.980 ;
        RECT 2881.050 17.920 2881.370 17.980 ;
        RECT 2676.810 17.780 2881.370 17.920 ;
        RECT 2676.810 17.720 2677.130 17.780 ;
        RECT 2881.050 17.720 2881.370 17.780 ;
      LAYER via ;
        RECT 2670.400 288.700 2670.660 288.960 ;
        RECT 2676.840 288.700 2677.100 288.960 ;
        RECT 2676.840 17.720 2677.100 17.980 ;
        RECT 2881.080 17.720 2881.340 17.980 ;
      LAYER met2 ;
        RECT 2670.400 300.000 2670.680 304.000 ;
        RECT 2670.460 288.990 2670.600 300.000 ;
        RECT 2670.400 288.670 2670.660 288.990 ;
        RECT 2676.840 288.670 2677.100 288.990 ;
        RECT 2676.900 18.010 2677.040 288.670 ;
        RECT 2676.840 17.690 2677.100 18.010 ;
        RECT 2881.080 17.690 2881.340 18.010 ;
        RECT 2881.140 2.400 2881.280 17.690 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2685.090 289.240 2685.410 289.300 ;
        RECT 2690.610 289.240 2690.930 289.300 ;
        RECT 2685.090 289.100 2690.930 289.240 ;
        RECT 2685.090 289.040 2685.410 289.100 ;
        RECT 2690.610 289.040 2690.930 289.100 ;
        RECT 2690.610 17.240 2690.930 17.300 ;
        RECT 2898.990 17.240 2899.310 17.300 ;
        RECT 2690.610 17.100 2899.310 17.240 ;
        RECT 2690.610 17.040 2690.930 17.100 ;
        RECT 2898.990 17.040 2899.310 17.100 ;
      LAYER via ;
        RECT 2685.120 289.040 2685.380 289.300 ;
        RECT 2690.640 289.040 2690.900 289.300 ;
        RECT 2690.640 17.040 2690.900 17.300 ;
        RECT 2899.020 17.040 2899.280 17.300 ;
      LAYER met2 ;
        RECT 2685.120 300.000 2685.400 304.000 ;
        RECT 2685.180 289.330 2685.320 300.000 ;
        RECT 2685.120 289.010 2685.380 289.330 ;
        RECT 2690.640 289.010 2690.900 289.330 ;
        RECT 2690.700 17.330 2690.840 289.010 ;
        RECT 2690.640 17.010 2690.900 17.330 ;
        RECT 2899.020 17.010 2899.280 17.330 ;
        RECT 2899.080 2.400 2899.220 17.010 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 955.565 17.765 955.735 19.635 ;
      LAYER mcon ;
        RECT 955.565 19.465 955.735 19.635 ;
      LAYER met1 ;
        RECT 955.505 19.620 955.795 19.665 ;
        RECT 994.130 19.620 994.450 19.680 ;
        RECT 955.505 19.480 994.450 19.620 ;
        RECT 955.505 19.435 955.795 19.480 ;
        RECT 994.130 19.420 994.450 19.480 ;
        RECT 846.930 17.920 847.250 17.980 ;
        RECT 955.505 17.920 955.795 17.965 ;
        RECT 846.930 17.780 955.795 17.920 ;
        RECT 846.930 17.720 847.250 17.780 ;
        RECT 955.505 17.735 955.795 17.780 ;
      LAYER via ;
        RECT 994.160 19.420 994.420 19.680 ;
        RECT 846.960 17.720 847.220 17.980 ;
      LAYER met2 ;
        RECT 995.080 300.290 995.360 304.000 ;
        RECT 994.220 300.150 995.360 300.290 ;
        RECT 994.220 19.710 994.360 300.150 ;
        RECT 995.080 300.000 995.360 300.150 ;
        RECT 994.160 19.390 994.420 19.710 ;
        RECT 846.960 17.690 847.220 18.010 ;
        RECT 847.020 2.400 847.160 17.690 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 864.870 18.940 865.190 19.000 ;
        RECT 1008.390 18.940 1008.710 19.000 ;
        RECT 864.870 18.800 1008.710 18.940 ;
        RECT 864.870 18.740 865.190 18.800 ;
        RECT 1008.390 18.740 1008.710 18.800 ;
      LAYER via ;
        RECT 864.900 18.740 865.160 19.000 ;
        RECT 1008.420 18.740 1008.680 19.000 ;
      LAYER met2 ;
        RECT 1009.800 300.290 1010.080 304.000 ;
        RECT 1007.560 300.150 1010.080 300.290 ;
        RECT 1007.560 21.490 1007.700 300.150 ;
        RECT 1009.800 300.000 1010.080 300.150 ;
        RECT 1007.560 21.350 1008.620 21.490 ;
        RECT 1008.480 19.030 1008.620 21.350 ;
        RECT 864.900 18.710 865.160 19.030 ;
        RECT 1008.420 18.710 1008.680 19.030 ;
        RECT 864.960 2.400 865.100 18.710 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.350 18.600 882.670 18.660 ;
        RECT 1021.270 18.600 1021.590 18.660 ;
        RECT 882.350 18.460 1021.590 18.600 ;
        RECT 882.350 18.400 882.670 18.460 ;
        RECT 1021.270 18.400 1021.590 18.460 ;
      LAYER via ;
        RECT 882.380 18.400 882.640 18.660 ;
        RECT 1021.300 18.400 1021.560 18.660 ;
      LAYER met2 ;
        RECT 1024.520 300.290 1024.800 304.000 ;
        RECT 1021.360 300.150 1024.800 300.290 ;
        RECT 1021.360 18.690 1021.500 300.150 ;
        RECT 1024.520 300.000 1024.800 300.150 ;
        RECT 882.380 18.370 882.640 18.690 ;
        RECT 1021.300 18.370 1021.560 18.690 ;
        RECT 882.440 9.250 882.580 18.370 ;
        RECT 882.440 9.110 883.040 9.250 ;
        RECT 882.900 2.400 883.040 9.110 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 900.750 19.280 901.070 19.340 ;
        RECT 1035.070 19.280 1035.390 19.340 ;
        RECT 900.750 19.140 1035.390 19.280 ;
        RECT 900.750 19.080 901.070 19.140 ;
        RECT 1035.070 19.080 1035.390 19.140 ;
      LAYER via ;
        RECT 900.780 19.080 901.040 19.340 ;
        RECT 1035.100 19.080 1035.360 19.340 ;
      LAYER met2 ;
        RECT 1039.240 300.290 1039.520 304.000 ;
        RECT 1035.160 300.150 1039.520 300.290 ;
        RECT 1035.160 19.370 1035.300 300.150 ;
        RECT 1039.240 300.000 1039.520 300.150 ;
        RECT 900.780 19.050 901.040 19.370 ;
        RECT 1035.100 19.050 1035.360 19.370 ;
        RECT 900.840 2.400 900.980 19.050 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 918.690 19.960 919.010 20.020 ;
        RECT 1049.330 19.960 1049.650 20.020 ;
        RECT 918.690 19.820 1049.650 19.960 ;
        RECT 918.690 19.760 919.010 19.820 ;
        RECT 1049.330 19.760 1049.650 19.820 ;
      LAYER via ;
        RECT 918.720 19.760 918.980 20.020 ;
        RECT 1049.360 19.760 1049.620 20.020 ;
      LAYER met2 ;
        RECT 1053.960 300.290 1054.240 304.000 ;
        RECT 1049.420 300.150 1054.240 300.290 ;
        RECT 1049.420 20.050 1049.560 300.150 ;
        RECT 1053.960 300.000 1054.240 300.150 ;
        RECT 918.720 19.730 918.980 20.050 ;
        RECT 1049.360 19.730 1049.620 20.050 ;
        RECT 918.780 2.400 918.920 19.730 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1062.745 89.845 1062.915 137.955 ;
      LAYER mcon ;
        RECT 1062.745 137.785 1062.915 137.955 ;
      LAYER met1 ;
        RECT 1063.130 241.640 1063.450 241.700 ;
        RECT 1067.270 241.640 1067.590 241.700 ;
        RECT 1063.130 241.500 1067.590 241.640 ;
        RECT 1063.130 241.440 1063.450 241.500 ;
        RECT 1067.270 241.440 1067.590 241.500 ;
        RECT 1062.670 206.960 1062.990 207.020 ;
        RECT 1063.590 206.960 1063.910 207.020 ;
        RECT 1062.670 206.820 1063.910 206.960 ;
        RECT 1062.670 206.760 1062.990 206.820 ;
        RECT 1063.590 206.760 1063.910 206.820 ;
        RECT 1062.670 137.940 1062.990 138.000 ;
        RECT 1062.475 137.800 1062.990 137.940 ;
        RECT 1062.670 137.740 1062.990 137.800 ;
        RECT 1062.685 90.000 1062.975 90.045 ;
        RECT 1063.130 90.000 1063.450 90.060 ;
        RECT 1062.685 89.860 1063.450 90.000 ;
        RECT 1062.685 89.815 1062.975 89.860 ;
        RECT 1063.130 89.800 1063.450 89.860 ;
        RECT 936.170 18.260 936.490 18.320 ;
        RECT 1063.590 18.260 1063.910 18.320 ;
        RECT 936.170 18.120 1063.910 18.260 ;
        RECT 936.170 18.060 936.490 18.120 ;
        RECT 1063.590 18.060 1063.910 18.120 ;
      LAYER via ;
        RECT 1063.160 241.440 1063.420 241.700 ;
        RECT 1067.300 241.440 1067.560 241.700 ;
        RECT 1062.700 206.760 1062.960 207.020 ;
        RECT 1063.620 206.760 1063.880 207.020 ;
        RECT 1062.700 137.740 1062.960 138.000 ;
        RECT 1063.160 89.800 1063.420 90.060 ;
        RECT 936.200 18.060 936.460 18.320 ;
        RECT 1063.620 18.060 1063.880 18.320 ;
      LAYER met2 ;
        RECT 1068.680 300.290 1068.960 304.000 ;
        RECT 1067.360 300.150 1068.960 300.290 ;
        RECT 1067.360 241.730 1067.500 300.150 ;
        RECT 1068.680 300.000 1068.960 300.150 ;
        RECT 1063.160 241.410 1063.420 241.730 ;
        RECT 1067.300 241.410 1067.560 241.730 ;
        RECT 1063.220 207.130 1063.360 241.410 ;
        RECT 1062.760 207.050 1063.360 207.130 ;
        RECT 1062.700 206.990 1063.360 207.050 ;
        RECT 1062.700 206.730 1062.960 206.990 ;
        RECT 1063.620 206.730 1063.880 207.050 ;
        RECT 1063.680 169.050 1063.820 206.730 ;
        RECT 1062.760 168.910 1063.820 169.050 ;
        RECT 1062.760 138.030 1062.900 168.910 ;
        RECT 1062.700 137.710 1062.960 138.030 ;
        RECT 1063.160 89.770 1063.420 90.090 ;
        RECT 1063.220 62.290 1063.360 89.770 ;
        RECT 1063.220 62.150 1063.820 62.290 ;
        RECT 1063.680 18.350 1063.820 62.150 ;
        RECT 936.200 18.030 936.460 18.350 ;
        RECT 1063.620 18.030 1063.880 18.350 ;
        RECT 936.260 2.400 936.400 18.030 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1003.865 19.465 1004.035 20.315 ;
      LAYER mcon ;
        RECT 1003.865 20.145 1004.035 20.315 ;
      LAYER met1 ;
        RECT 954.110 20.300 954.430 20.360 ;
        RECT 1003.805 20.300 1004.095 20.345 ;
        RECT 954.110 20.160 1004.095 20.300 ;
        RECT 954.110 20.100 954.430 20.160 ;
        RECT 1003.805 20.115 1004.095 20.160 ;
        RECT 1003.805 19.620 1004.095 19.665 ;
        RECT 1083.370 19.620 1083.690 19.680 ;
        RECT 1003.805 19.480 1083.690 19.620 ;
        RECT 1003.805 19.435 1004.095 19.480 ;
        RECT 1083.370 19.420 1083.690 19.480 ;
      LAYER via ;
        RECT 954.140 20.100 954.400 20.360 ;
        RECT 1083.400 19.420 1083.660 19.680 ;
      LAYER met2 ;
        RECT 1083.400 300.000 1083.680 304.000 ;
        RECT 954.140 20.070 954.400 20.390 ;
        RECT 954.200 2.400 954.340 20.070 ;
        RECT 1083.460 19.710 1083.600 300.000 ;
        RECT 1083.400 19.390 1083.660 19.710 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.050 17.240 972.370 17.300 ;
        RECT 1097.630 17.240 1097.950 17.300 ;
        RECT 972.050 17.100 1097.950 17.240 ;
        RECT 972.050 17.040 972.370 17.100 ;
        RECT 1097.630 17.040 1097.950 17.100 ;
      LAYER via ;
        RECT 972.080 17.040 972.340 17.300 ;
        RECT 1097.660 17.040 1097.920 17.300 ;
      LAYER met2 ;
        RECT 1098.120 300.290 1098.400 304.000 ;
        RECT 1097.720 300.150 1098.400 300.290 ;
        RECT 1097.720 17.330 1097.860 300.150 ;
        RECT 1098.120 300.000 1098.400 300.150 ;
        RECT 972.080 17.010 972.340 17.330 ;
        RECT 1097.660 17.010 1097.920 17.330 ;
        RECT 972.140 2.400 972.280 17.010 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 828.070 279.380 828.390 279.440 ;
        RECT 831.750 279.380 832.070 279.440 ;
        RECT 828.070 279.240 832.070 279.380 ;
        RECT 828.070 279.180 828.390 279.240 ;
        RECT 831.750 279.180 832.070 279.240 ;
        RECT 650.970 19.280 651.290 19.340 ;
        RECT 828.070 19.280 828.390 19.340 ;
        RECT 650.970 19.140 828.390 19.280 ;
        RECT 650.970 19.080 651.290 19.140 ;
        RECT 828.070 19.080 828.390 19.140 ;
      LAYER via ;
        RECT 828.100 279.180 828.360 279.440 ;
        RECT 831.780 279.180 832.040 279.440 ;
        RECT 651.000 19.080 651.260 19.340 ;
        RECT 828.100 19.080 828.360 19.340 ;
      LAYER met2 ;
        RECT 833.620 300.290 833.900 304.000 ;
        RECT 831.840 300.150 833.900 300.290 ;
        RECT 831.840 279.470 831.980 300.150 ;
        RECT 833.620 300.000 833.900 300.150 ;
        RECT 828.100 279.150 828.360 279.470 ;
        RECT 831.780 279.150 832.040 279.470 ;
        RECT 828.160 19.370 828.300 279.150 ;
        RECT 651.000 19.050 651.260 19.370 ;
        RECT 828.100 19.050 828.360 19.370 ;
        RECT 651.060 2.400 651.200 19.050 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 993.210 286.180 993.530 286.240 ;
        RECT 1112.810 286.180 1113.130 286.240 ;
        RECT 993.210 286.040 1113.130 286.180 ;
        RECT 993.210 285.980 993.530 286.040 ;
        RECT 1112.810 285.980 1113.130 286.040 ;
        RECT 989.990 14.860 990.310 14.920 ;
        RECT 993.210 14.860 993.530 14.920 ;
        RECT 989.990 14.720 993.530 14.860 ;
        RECT 989.990 14.660 990.310 14.720 ;
        RECT 993.210 14.660 993.530 14.720 ;
      LAYER via ;
        RECT 993.240 285.980 993.500 286.240 ;
        RECT 1112.840 285.980 1113.100 286.240 ;
        RECT 990.020 14.660 990.280 14.920 ;
        RECT 993.240 14.660 993.500 14.920 ;
      LAYER met2 ;
        RECT 1112.840 300.000 1113.120 304.000 ;
        RECT 1112.900 286.270 1113.040 300.000 ;
        RECT 993.240 285.950 993.500 286.270 ;
        RECT 1112.840 285.950 1113.100 286.270 ;
        RECT 993.300 14.950 993.440 285.950 ;
        RECT 990.020 14.630 990.280 14.950 ;
        RECT 993.240 14.630 993.500 14.950 ;
        RECT 990.080 2.400 990.220 14.630 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1013.450 284.820 1013.770 284.880 ;
        RECT 1127.530 284.820 1127.850 284.880 ;
        RECT 1013.450 284.680 1127.850 284.820 ;
        RECT 1013.450 284.620 1013.770 284.680 ;
        RECT 1127.530 284.620 1127.850 284.680 ;
        RECT 1007.470 20.640 1007.790 20.700 ;
        RECT 1013.450 20.640 1013.770 20.700 ;
        RECT 1007.470 20.500 1013.770 20.640 ;
        RECT 1007.470 20.440 1007.790 20.500 ;
        RECT 1013.450 20.440 1013.770 20.500 ;
      LAYER via ;
        RECT 1013.480 284.620 1013.740 284.880 ;
        RECT 1127.560 284.620 1127.820 284.880 ;
        RECT 1007.500 20.440 1007.760 20.700 ;
        RECT 1013.480 20.440 1013.740 20.700 ;
      LAYER met2 ;
        RECT 1127.560 300.000 1127.840 304.000 ;
        RECT 1127.620 284.910 1127.760 300.000 ;
        RECT 1013.480 284.590 1013.740 284.910 ;
        RECT 1127.560 284.590 1127.820 284.910 ;
        RECT 1013.540 20.730 1013.680 284.590 ;
        RECT 1007.500 20.410 1007.760 20.730 ;
        RECT 1013.480 20.410 1013.740 20.730 ;
        RECT 1007.560 2.400 1007.700 20.410 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1027.710 286.860 1028.030 286.920 ;
        RECT 1142.250 286.860 1142.570 286.920 ;
        RECT 1027.710 286.720 1142.570 286.860 ;
        RECT 1027.710 286.660 1028.030 286.720 ;
        RECT 1142.250 286.660 1142.570 286.720 ;
        RECT 1025.410 20.640 1025.730 20.700 ;
        RECT 1027.710 20.640 1028.030 20.700 ;
        RECT 1025.410 20.500 1028.030 20.640 ;
        RECT 1025.410 20.440 1025.730 20.500 ;
        RECT 1027.710 20.440 1028.030 20.500 ;
      LAYER via ;
        RECT 1027.740 286.660 1028.000 286.920 ;
        RECT 1142.280 286.660 1142.540 286.920 ;
        RECT 1025.440 20.440 1025.700 20.700 ;
        RECT 1027.740 20.440 1028.000 20.700 ;
      LAYER met2 ;
        RECT 1142.280 300.000 1142.560 304.000 ;
        RECT 1142.340 286.950 1142.480 300.000 ;
        RECT 1027.740 286.630 1028.000 286.950 ;
        RECT 1142.280 286.630 1142.540 286.950 ;
        RECT 1027.800 20.730 1027.940 286.630 ;
        RECT 1025.440 20.410 1025.700 20.730 ;
        RECT 1027.740 20.410 1028.000 20.730 ;
        RECT 1025.500 2.400 1025.640 20.410 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1048.410 284.140 1048.730 284.200 ;
        RECT 1156.970 284.140 1157.290 284.200 ;
        RECT 1048.410 284.000 1157.290 284.140 ;
        RECT 1048.410 283.940 1048.730 284.000 ;
        RECT 1156.970 283.940 1157.290 284.000 ;
        RECT 1043.350 20.640 1043.670 20.700 ;
        RECT 1048.410 20.640 1048.730 20.700 ;
        RECT 1043.350 20.500 1048.730 20.640 ;
        RECT 1043.350 20.440 1043.670 20.500 ;
        RECT 1048.410 20.440 1048.730 20.500 ;
      LAYER via ;
        RECT 1048.440 283.940 1048.700 284.200 ;
        RECT 1157.000 283.940 1157.260 284.200 ;
        RECT 1043.380 20.440 1043.640 20.700 ;
        RECT 1048.440 20.440 1048.700 20.700 ;
      LAYER met2 ;
        RECT 1157.000 300.000 1157.280 304.000 ;
        RECT 1157.060 284.230 1157.200 300.000 ;
        RECT 1048.440 283.910 1048.700 284.230 ;
        RECT 1157.000 283.910 1157.260 284.230 ;
        RECT 1048.500 20.730 1048.640 283.910 ;
        RECT 1043.380 20.410 1043.640 20.730 ;
        RECT 1048.440 20.410 1048.700 20.730 ;
        RECT 1043.440 2.400 1043.580 20.410 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1062.285 2.805 1062.455 48.195 ;
      LAYER mcon ;
        RECT 1062.285 48.025 1062.455 48.195 ;
      LAYER met1 ;
        RECT 1062.210 283.800 1062.530 283.860 ;
        RECT 1171.690 283.800 1172.010 283.860 ;
        RECT 1062.210 283.660 1172.010 283.800 ;
        RECT 1062.210 283.600 1062.530 283.660 ;
        RECT 1171.690 283.600 1172.010 283.660 ;
        RECT 1062.210 48.180 1062.530 48.240 ;
        RECT 1062.015 48.040 1062.530 48.180 ;
        RECT 1062.210 47.980 1062.530 48.040 ;
        RECT 1061.290 2.960 1061.610 3.020 ;
        RECT 1062.225 2.960 1062.515 3.005 ;
        RECT 1061.290 2.820 1062.515 2.960 ;
        RECT 1061.290 2.760 1061.610 2.820 ;
        RECT 1062.225 2.775 1062.515 2.820 ;
      LAYER via ;
        RECT 1062.240 283.600 1062.500 283.860 ;
        RECT 1171.720 283.600 1171.980 283.860 ;
        RECT 1062.240 47.980 1062.500 48.240 ;
        RECT 1061.320 2.760 1061.580 3.020 ;
      LAYER met2 ;
        RECT 1171.720 300.000 1172.000 304.000 ;
        RECT 1171.780 283.890 1171.920 300.000 ;
        RECT 1062.240 283.570 1062.500 283.890 ;
        RECT 1171.720 283.570 1171.980 283.890 ;
        RECT 1062.300 48.270 1062.440 283.570 ;
        RECT 1062.240 47.950 1062.500 48.270 ;
        RECT 1061.320 2.730 1061.580 3.050 ;
        RECT 1061.380 2.400 1061.520 2.730 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1082.910 283.120 1083.230 283.180 ;
        RECT 1185.030 283.120 1185.350 283.180 ;
        RECT 1082.910 282.980 1185.350 283.120 ;
        RECT 1082.910 282.920 1083.230 282.980 ;
        RECT 1185.030 282.920 1185.350 282.980 ;
        RECT 1079.230 17.580 1079.550 17.640 ;
        RECT 1082.910 17.580 1083.230 17.640 ;
        RECT 1079.230 17.440 1083.230 17.580 ;
        RECT 1079.230 17.380 1079.550 17.440 ;
        RECT 1082.910 17.380 1083.230 17.440 ;
      LAYER via ;
        RECT 1082.940 282.920 1083.200 283.180 ;
        RECT 1185.060 282.920 1185.320 283.180 ;
        RECT 1079.260 17.380 1079.520 17.640 ;
        RECT 1082.940 17.380 1083.200 17.640 ;
      LAYER met2 ;
        RECT 1186.440 300.290 1186.720 304.000 ;
        RECT 1185.120 300.150 1186.720 300.290 ;
        RECT 1185.120 283.210 1185.260 300.150 ;
        RECT 1186.440 300.000 1186.720 300.150 ;
        RECT 1082.940 282.890 1083.200 283.210 ;
        RECT 1185.060 282.890 1185.320 283.210 ;
        RECT 1083.000 17.670 1083.140 282.890 ;
        RECT 1079.260 17.350 1079.520 17.670 ;
        RECT 1082.940 17.350 1083.200 17.670 ;
        RECT 1079.320 2.400 1079.460 17.350 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.250 287.540 1096.570 287.600 ;
        RECT 1201.130 287.540 1201.450 287.600 ;
        RECT 1096.250 287.400 1201.450 287.540 ;
        RECT 1096.250 287.340 1096.570 287.400 ;
        RECT 1201.130 287.340 1201.450 287.400 ;
      LAYER via ;
        RECT 1096.280 287.340 1096.540 287.600 ;
        RECT 1201.160 287.340 1201.420 287.600 ;
      LAYER met2 ;
        RECT 1201.160 300.000 1201.440 304.000 ;
        RECT 1201.220 287.630 1201.360 300.000 ;
        RECT 1096.280 287.310 1096.540 287.630 ;
        RECT 1201.160 287.310 1201.420 287.630 ;
        RECT 1096.340 17.410 1096.480 287.310 ;
        RECT 1096.340 17.270 1096.940 17.410 ;
        RECT 1096.800 2.400 1096.940 17.270 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1117.410 286.180 1117.730 286.240 ;
        RECT 1215.390 286.180 1215.710 286.240 ;
        RECT 1117.410 286.040 1215.710 286.180 ;
        RECT 1117.410 285.980 1117.730 286.040 ;
        RECT 1215.390 285.980 1215.710 286.040 ;
        RECT 1114.650 17.580 1114.970 17.640 ;
        RECT 1117.410 17.580 1117.730 17.640 ;
        RECT 1114.650 17.440 1117.730 17.580 ;
        RECT 1114.650 17.380 1114.970 17.440 ;
        RECT 1117.410 17.380 1117.730 17.440 ;
      LAYER via ;
        RECT 1117.440 285.980 1117.700 286.240 ;
        RECT 1215.420 285.980 1215.680 286.240 ;
        RECT 1114.680 17.380 1114.940 17.640 ;
        RECT 1117.440 17.380 1117.700 17.640 ;
      LAYER met2 ;
        RECT 1215.420 300.000 1215.700 304.000 ;
        RECT 1215.480 286.270 1215.620 300.000 ;
        RECT 1117.440 285.950 1117.700 286.270 ;
        RECT 1215.420 285.950 1215.680 286.270 ;
        RECT 1117.500 17.670 1117.640 285.950 ;
        RECT 1114.680 17.350 1114.940 17.670 ;
        RECT 1117.440 17.350 1117.700 17.670 ;
        RECT 1114.740 2.400 1114.880 17.350 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1138.110 284.820 1138.430 284.880 ;
        RECT 1230.110 284.820 1230.430 284.880 ;
        RECT 1138.110 284.680 1230.430 284.820 ;
        RECT 1138.110 284.620 1138.430 284.680 ;
        RECT 1230.110 284.620 1230.430 284.680 ;
        RECT 1132.590 17.580 1132.910 17.640 ;
        RECT 1138.110 17.580 1138.430 17.640 ;
        RECT 1132.590 17.440 1138.430 17.580 ;
        RECT 1132.590 17.380 1132.910 17.440 ;
        RECT 1138.110 17.380 1138.430 17.440 ;
      LAYER via ;
        RECT 1138.140 284.620 1138.400 284.880 ;
        RECT 1230.140 284.620 1230.400 284.880 ;
        RECT 1132.620 17.380 1132.880 17.640 ;
        RECT 1138.140 17.380 1138.400 17.640 ;
      LAYER met2 ;
        RECT 1230.140 300.000 1230.420 304.000 ;
        RECT 1230.200 284.910 1230.340 300.000 ;
        RECT 1138.140 284.590 1138.400 284.910 ;
        RECT 1230.140 284.590 1230.400 284.910 ;
        RECT 1138.200 17.670 1138.340 284.590 ;
        RECT 1132.620 17.350 1132.880 17.670 ;
        RECT 1138.140 17.350 1138.400 17.670 ;
        RECT 1132.680 2.400 1132.820 17.350 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1152.370 287.200 1152.690 287.260 ;
        RECT 1244.830 287.200 1245.150 287.260 ;
        RECT 1152.370 287.060 1245.150 287.200 ;
        RECT 1152.370 287.000 1152.690 287.060 ;
        RECT 1244.830 287.000 1245.150 287.060 ;
      LAYER via ;
        RECT 1152.400 287.000 1152.660 287.260 ;
        RECT 1244.860 287.000 1245.120 287.260 ;
      LAYER met2 ;
        RECT 1244.860 300.000 1245.140 304.000 ;
        RECT 1244.920 287.290 1245.060 300.000 ;
        RECT 1152.400 286.970 1152.660 287.290 ;
        RECT 1244.860 286.970 1245.120 287.290 ;
        RECT 1152.460 286.010 1152.600 286.970 ;
        RECT 1152.000 285.870 1152.600 286.010 ;
        RECT 1152.000 17.410 1152.140 285.870 ;
        RECT 1150.620 17.270 1152.140 17.410 ;
        RECT 1150.620 2.400 1150.760 17.270 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 841.870 286.520 842.190 286.580 ;
        RECT 846.470 286.520 846.790 286.580 ;
        RECT 841.870 286.380 846.790 286.520 ;
        RECT 841.870 286.320 842.190 286.380 ;
        RECT 846.470 286.320 846.790 286.380 ;
        RECT 668.910 18.940 669.230 19.000 ;
        RECT 841.870 18.940 842.190 19.000 ;
        RECT 668.910 18.800 842.190 18.940 ;
        RECT 668.910 18.740 669.230 18.800 ;
        RECT 841.870 18.740 842.190 18.800 ;
      LAYER via ;
        RECT 841.900 286.320 842.160 286.580 ;
        RECT 846.500 286.320 846.760 286.580 ;
        RECT 668.940 18.740 669.200 19.000 ;
        RECT 841.900 18.740 842.160 19.000 ;
      LAYER met2 ;
        RECT 848.340 300.290 848.620 304.000 ;
        RECT 846.560 300.150 848.620 300.290 ;
        RECT 846.560 286.610 846.700 300.150 ;
        RECT 848.340 300.000 848.620 300.150 ;
        RECT 841.900 286.290 842.160 286.610 ;
        RECT 846.500 286.290 846.760 286.610 ;
        RECT 841.960 19.030 842.100 286.290 ;
        RECT 668.940 18.710 669.200 19.030 ;
        RECT 841.900 18.710 842.160 19.030 ;
        RECT 669.000 2.400 669.140 18.710 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1172.610 284.140 1172.930 284.200 ;
        RECT 1259.550 284.140 1259.870 284.200 ;
        RECT 1172.610 284.000 1259.870 284.140 ;
        RECT 1172.610 283.940 1172.930 284.000 ;
        RECT 1259.550 283.940 1259.870 284.000 ;
        RECT 1168.470 17.580 1168.790 17.640 ;
        RECT 1172.610 17.580 1172.930 17.640 ;
        RECT 1168.470 17.440 1172.930 17.580 ;
        RECT 1168.470 17.380 1168.790 17.440 ;
        RECT 1172.610 17.380 1172.930 17.440 ;
      LAYER via ;
        RECT 1172.640 283.940 1172.900 284.200 ;
        RECT 1259.580 283.940 1259.840 284.200 ;
        RECT 1168.500 17.380 1168.760 17.640 ;
        RECT 1172.640 17.380 1172.900 17.640 ;
      LAYER met2 ;
        RECT 1259.580 300.000 1259.860 304.000 ;
        RECT 1259.640 284.230 1259.780 300.000 ;
        RECT 1172.640 283.910 1172.900 284.230 ;
        RECT 1259.580 283.910 1259.840 284.230 ;
        RECT 1172.700 17.670 1172.840 283.910 ;
        RECT 1168.500 17.350 1168.760 17.670 ;
        RECT 1172.640 17.350 1172.900 17.670 ;
        RECT 1168.560 2.400 1168.700 17.350 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1185.950 287.880 1186.270 287.940 ;
        RECT 1274.270 287.880 1274.590 287.940 ;
        RECT 1185.950 287.740 1274.590 287.880 ;
        RECT 1185.950 287.680 1186.270 287.740 ;
        RECT 1274.270 287.680 1274.590 287.740 ;
      LAYER via ;
        RECT 1185.980 287.680 1186.240 287.940 ;
        RECT 1274.300 287.680 1274.560 287.940 ;
      LAYER met2 ;
        RECT 1274.300 300.000 1274.580 304.000 ;
        RECT 1274.360 287.970 1274.500 300.000 ;
        RECT 1185.980 287.650 1186.240 287.970 ;
        RECT 1274.300 287.650 1274.560 287.970 ;
        RECT 1186.040 2.400 1186.180 287.650 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1207.110 287.540 1207.430 287.600 ;
        RECT 1288.990 287.540 1289.310 287.600 ;
        RECT 1207.110 287.400 1289.310 287.540 ;
        RECT 1207.110 287.340 1207.430 287.400 ;
        RECT 1288.990 287.340 1289.310 287.400 ;
        RECT 1203.890 17.580 1204.210 17.640 ;
        RECT 1207.110 17.580 1207.430 17.640 ;
        RECT 1203.890 17.440 1207.430 17.580 ;
        RECT 1203.890 17.380 1204.210 17.440 ;
        RECT 1207.110 17.380 1207.430 17.440 ;
      LAYER via ;
        RECT 1207.140 287.340 1207.400 287.600 ;
        RECT 1289.020 287.340 1289.280 287.600 ;
        RECT 1203.920 17.380 1204.180 17.640 ;
        RECT 1207.140 17.380 1207.400 17.640 ;
      LAYER met2 ;
        RECT 1289.020 300.000 1289.300 304.000 ;
        RECT 1289.080 287.630 1289.220 300.000 ;
        RECT 1207.140 287.310 1207.400 287.630 ;
        RECT 1289.020 287.310 1289.280 287.630 ;
        RECT 1207.200 17.670 1207.340 287.310 ;
        RECT 1203.920 17.350 1204.180 17.670 ;
        RECT 1207.140 17.350 1207.400 17.670 ;
        RECT 1203.980 2.400 1204.120 17.350 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1227.350 284.480 1227.670 284.540 ;
        RECT 1301.870 284.480 1302.190 284.540 ;
        RECT 1227.350 284.340 1302.190 284.480 ;
        RECT 1227.350 284.280 1227.670 284.340 ;
        RECT 1301.870 284.280 1302.190 284.340 ;
        RECT 1221.830 17.580 1222.150 17.640 ;
        RECT 1227.350 17.580 1227.670 17.640 ;
        RECT 1221.830 17.440 1227.670 17.580 ;
        RECT 1221.830 17.380 1222.150 17.440 ;
        RECT 1227.350 17.380 1227.670 17.440 ;
      LAYER via ;
        RECT 1227.380 284.280 1227.640 284.540 ;
        RECT 1301.900 284.280 1302.160 284.540 ;
        RECT 1221.860 17.380 1222.120 17.640 ;
        RECT 1227.380 17.380 1227.640 17.640 ;
      LAYER met2 ;
        RECT 1303.740 300.290 1304.020 304.000 ;
        RECT 1301.960 300.150 1304.020 300.290 ;
        RECT 1301.960 284.570 1302.100 300.150 ;
        RECT 1303.740 300.000 1304.020 300.150 ;
        RECT 1227.380 284.250 1227.640 284.570 ;
        RECT 1301.900 284.250 1302.160 284.570 ;
        RECT 1227.440 17.670 1227.580 284.250 ;
        RECT 1221.860 17.350 1222.120 17.670 ;
        RECT 1227.380 17.350 1227.640 17.670 ;
        RECT 1221.920 2.400 1222.060 17.350 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1241.610 286.520 1241.930 286.580 ;
        RECT 1318.430 286.520 1318.750 286.580 ;
        RECT 1241.610 286.380 1318.750 286.520 ;
        RECT 1241.610 286.320 1241.930 286.380 ;
        RECT 1318.430 286.320 1318.750 286.380 ;
      LAYER via ;
        RECT 1241.640 286.320 1241.900 286.580 ;
        RECT 1318.460 286.320 1318.720 286.580 ;
      LAYER met2 ;
        RECT 1318.460 300.000 1318.740 304.000 ;
        RECT 1318.520 286.610 1318.660 300.000 ;
        RECT 1241.640 286.290 1241.900 286.610 ;
        RECT 1318.460 286.290 1318.720 286.610 ;
        RECT 1241.700 17.410 1241.840 286.290 ;
        RECT 1239.860 17.270 1241.840 17.410 ;
        RECT 1239.860 2.400 1240.000 17.270 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1262.310 288.220 1262.630 288.280 ;
        RECT 1333.150 288.220 1333.470 288.280 ;
        RECT 1262.310 288.080 1333.470 288.220 ;
        RECT 1262.310 288.020 1262.630 288.080 ;
        RECT 1333.150 288.020 1333.470 288.080 ;
        RECT 1257.250 17.580 1257.570 17.640 ;
        RECT 1262.310 17.580 1262.630 17.640 ;
        RECT 1257.250 17.440 1262.630 17.580 ;
        RECT 1257.250 17.380 1257.570 17.440 ;
        RECT 1262.310 17.380 1262.630 17.440 ;
      LAYER via ;
        RECT 1262.340 288.020 1262.600 288.280 ;
        RECT 1333.180 288.020 1333.440 288.280 ;
        RECT 1257.280 17.380 1257.540 17.640 ;
        RECT 1262.340 17.380 1262.600 17.640 ;
      LAYER met2 ;
        RECT 1333.180 300.000 1333.460 304.000 ;
        RECT 1333.240 288.310 1333.380 300.000 ;
        RECT 1262.340 287.990 1262.600 288.310 ;
        RECT 1333.180 287.990 1333.440 288.310 ;
        RECT 1262.400 17.670 1262.540 287.990 ;
        RECT 1257.280 17.350 1257.540 17.670 ;
        RECT 1262.340 17.350 1262.600 17.670 ;
        RECT 1257.340 2.400 1257.480 17.350 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1276.110 288.560 1276.430 288.620 ;
        RECT 1347.870 288.560 1348.190 288.620 ;
        RECT 1276.110 288.420 1348.190 288.560 ;
        RECT 1276.110 288.360 1276.430 288.420 ;
        RECT 1347.870 288.360 1348.190 288.420 ;
      LAYER via ;
        RECT 1276.140 288.360 1276.400 288.620 ;
        RECT 1347.900 288.360 1348.160 288.620 ;
      LAYER met2 ;
        RECT 1347.900 300.000 1348.180 304.000 ;
        RECT 1347.960 288.650 1348.100 300.000 ;
        RECT 1276.140 288.330 1276.400 288.650 ;
        RECT 1347.900 288.330 1348.160 288.650 ;
        RECT 1276.200 17.410 1276.340 288.330 ;
        RECT 1275.280 17.270 1276.340 17.410 ;
        RECT 1275.280 2.400 1275.420 17.270 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1296.810 289.240 1297.130 289.300 ;
        RECT 1362.590 289.240 1362.910 289.300 ;
        RECT 1296.810 289.100 1362.910 289.240 ;
        RECT 1296.810 289.040 1297.130 289.100 ;
        RECT 1362.590 289.040 1362.910 289.100 ;
        RECT 1293.130 15.540 1293.450 15.600 ;
        RECT 1296.810 15.540 1297.130 15.600 ;
        RECT 1293.130 15.400 1297.130 15.540 ;
        RECT 1293.130 15.340 1293.450 15.400 ;
        RECT 1296.810 15.340 1297.130 15.400 ;
      LAYER via ;
        RECT 1296.840 289.040 1297.100 289.300 ;
        RECT 1362.620 289.040 1362.880 289.300 ;
        RECT 1293.160 15.340 1293.420 15.600 ;
        RECT 1296.840 15.340 1297.100 15.600 ;
      LAYER met2 ;
        RECT 1362.620 300.000 1362.900 304.000 ;
        RECT 1362.680 289.330 1362.820 300.000 ;
        RECT 1296.840 289.010 1297.100 289.330 ;
        RECT 1362.620 289.010 1362.880 289.330 ;
        RECT 1296.900 15.630 1297.040 289.010 ;
        RECT 1293.160 15.310 1293.420 15.630 ;
        RECT 1296.840 15.310 1297.100 15.630 ;
        RECT 1293.220 2.400 1293.360 15.310 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1317.510 289.580 1317.830 289.640 ;
        RECT 1377.310 289.580 1377.630 289.640 ;
        RECT 1317.510 289.440 1377.630 289.580 ;
        RECT 1317.510 289.380 1317.830 289.440 ;
        RECT 1377.310 289.380 1377.630 289.440 ;
        RECT 1311.070 17.580 1311.390 17.640 ;
        RECT 1317.510 17.580 1317.830 17.640 ;
        RECT 1311.070 17.440 1317.830 17.580 ;
        RECT 1311.070 17.380 1311.390 17.440 ;
        RECT 1317.510 17.380 1317.830 17.440 ;
      LAYER via ;
        RECT 1317.540 289.380 1317.800 289.640 ;
        RECT 1377.340 289.380 1377.600 289.640 ;
        RECT 1311.100 17.380 1311.360 17.640 ;
        RECT 1317.540 17.380 1317.800 17.640 ;
      LAYER met2 ;
        RECT 1377.340 300.000 1377.620 304.000 ;
        RECT 1377.400 289.670 1377.540 300.000 ;
        RECT 1317.540 289.350 1317.800 289.670 ;
        RECT 1377.340 289.350 1377.600 289.670 ;
        RECT 1317.600 17.670 1317.740 289.350 ;
        RECT 1311.100 17.350 1311.360 17.670 ;
        RECT 1317.540 17.350 1317.800 17.670 ;
        RECT 1311.160 2.400 1311.300 17.350 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1331.310 287.200 1331.630 287.260 ;
        RECT 1392.030 287.200 1392.350 287.260 ;
        RECT 1331.310 287.060 1392.350 287.200 ;
        RECT 1331.310 287.000 1331.630 287.060 ;
        RECT 1392.030 287.000 1392.350 287.060 ;
        RECT 1329.010 17.580 1329.330 17.640 ;
        RECT 1331.310 17.580 1331.630 17.640 ;
        RECT 1329.010 17.440 1331.630 17.580 ;
        RECT 1329.010 17.380 1329.330 17.440 ;
        RECT 1331.310 17.380 1331.630 17.440 ;
      LAYER via ;
        RECT 1331.340 287.000 1331.600 287.260 ;
        RECT 1392.060 287.000 1392.320 287.260 ;
        RECT 1329.040 17.380 1329.300 17.640 ;
        RECT 1331.340 17.380 1331.600 17.640 ;
      LAYER met2 ;
        RECT 1392.060 300.000 1392.340 304.000 ;
        RECT 1392.120 287.290 1392.260 300.000 ;
        RECT 1331.340 286.970 1331.600 287.290 ;
        RECT 1392.060 286.970 1392.320 287.290 ;
        RECT 1331.400 17.670 1331.540 286.970 ;
        RECT 1329.040 17.350 1329.300 17.670 ;
        RECT 1331.340 17.350 1331.600 17.670 ;
        RECT 1329.100 2.400 1329.240 17.350 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 831.365 16.405 831.535 18.615 ;
      LAYER mcon ;
        RECT 831.365 18.445 831.535 18.615 ;
      LAYER met1 ;
        RECT 686.390 18.600 686.710 18.660 ;
        RECT 831.305 18.600 831.595 18.645 ;
        RECT 686.390 18.460 831.595 18.600 ;
        RECT 686.390 18.400 686.710 18.460 ;
        RECT 831.305 18.415 831.595 18.460 ;
        RECT 831.305 16.560 831.595 16.605 ;
        RECT 863.490 16.560 863.810 16.620 ;
        RECT 831.305 16.420 863.810 16.560 ;
        RECT 831.305 16.375 831.595 16.420 ;
        RECT 863.490 16.360 863.810 16.420 ;
      LAYER via ;
        RECT 686.420 18.400 686.680 18.660 ;
        RECT 863.520 16.360 863.780 16.620 ;
      LAYER met2 ;
        RECT 863.060 300.290 863.340 304.000 ;
        RECT 863.060 300.150 863.720 300.290 ;
        RECT 863.060 300.000 863.340 300.150 ;
        RECT 686.420 18.370 686.680 18.690 ;
        RECT 686.480 2.400 686.620 18.370 ;
        RECT 863.580 16.650 863.720 300.150 ;
        RECT 863.520 16.330 863.780 16.650 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1352.010 285.160 1352.330 285.220 ;
        RECT 1406.750 285.160 1407.070 285.220 ;
        RECT 1352.010 285.020 1407.070 285.160 ;
        RECT 1352.010 284.960 1352.330 285.020 ;
        RECT 1406.750 284.960 1407.070 285.020 ;
        RECT 1346.490 17.580 1346.810 17.640 ;
        RECT 1352.010 17.580 1352.330 17.640 ;
        RECT 1346.490 17.440 1352.330 17.580 ;
        RECT 1346.490 17.380 1346.810 17.440 ;
        RECT 1352.010 17.380 1352.330 17.440 ;
      LAYER via ;
        RECT 1352.040 284.960 1352.300 285.220 ;
        RECT 1406.780 284.960 1407.040 285.220 ;
        RECT 1346.520 17.380 1346.780 17.640 ;
        RECT 1352.040 17.380 1352.300 17.640 ;
      LAYER met2 ;
        RECT 1406.780 300.000 1407.060 304.000 ;
        RECT 1406.840 285.250 1406.980 300.000 ;
        RECT 1352.040 284.930 1352.300 285.250 ;
        RECT 1406.780 284.930 1407.040 285.250 ;
        RECT 1352.100 17.670 1352.240 284.930 ;
        RECT 1346.520 17.350 1346.780 17.670 ;
        RECT 1352.040 17.350 1352.300 17.670 ;
        RECT 1346.580 2.400 1346.720 17.350 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1365.810 287.880 1366.130 287.940 ;
        RECT 1421.470 287.880 1421.790 287.940 ;
        RECT 1365.810 287.740 1421.790 287.880 ;
        RECT 1365.810 287.680 1366.130 287.740 ;
        RECT 1421.470 287.680 1421.790 287.740 ;
      LAYER via ;
        RECT 1365.840 287.680 1366.100 287.940 ;
        RECT 1421.500 287.680 1421.760 287.940 ;
      LAYER met2 ;
        RECT 1421.500 300.000 1421.780 304.000 ;
        RECT 1421.560 287.970 1421.700 300.000 ;
        RECT 1365.840 287.650 1366.100 287.970 ;
        RECT 1421.500 287.650 1421.760 287.970 ;
        RECT 1365.900 17.410 1366.040 287.650 ;
        RECT 1364.520 17.270 1366.040 17.410 ;
        RECT 1364.520 2.400 1364.660 17.270 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1386.510 287.540 1386.830 287.600 ;
        RECT 1436.190 287.540 1436.510 287.600 ;
        RECT 1386.510 287.400 1436.510 287.540 ;
        RECT 1386.510 287.340 1386.830 287.400 ;
        RECT 1436.190 287.340 1436.510 287.400 ;
        RECT 1382.370 17.580 1382.690 17.640 ;
        RECT 1386.510 17.580 1386.830 17.640 ;
        RECT 1382.370 17.440 1386.830 17.580 ;
        RECT 1382.370 17.380 1382.690 17.440 ;
        RECT 1386.510 17.380 1386.830 17.440 ;
      LAYER via ;
        RECT 1386.540 287.340 1386.800 287.600 ;
        RECT 1436.220 287.340 1436.480 287.600 ;
        RECT 1382.400 17.380 1382.660 17.640 ;
        RECT 1386.540 17.380 1386.800 17.640 ;
      LAYER met2 ;
        RECT 1436.220 300.000 1436.500 304.000 ;
        RECT 1436.280 287.630 1436.420 300.000 ;
        RECT 1386.540 287.310 1386.800 287.630 ;
        RECT 1436.220 287.310 1436.480 287.630 ;
        RECT 1386.600 17.670 1386.740 287.310 ;
        RECT 1382.400 17.350 1382.660 17.670 ;
        RECT 1386.540 17.350 1386.800 17.670 ;
        RECT 1382.460 2.400 1382.600 17.350 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1399.850 286.180 1400.170 286.240 ;
        RECT 1450.910 286.180 1451.230 286.240 ;
        RECT 1399.850 286.040 1451.230 286.180 ;
        RECT 1399.850 285.980 1400.170 286.040 ;
        RECT 1450.910 285.980 1451.230 286.040 ;
      LAYER via ;
        RECT 1399.880 285.980 1400.140 286.240 ;
        RECT 1450.940 285.980 1451.200 286.240 ;
      LAYER met2 ;
        RECT 1450.940 300.000 1451.220 304.000 ;
        RECT 1451.000 286.270 1451.140 300.000 ;
        RECT 1399.880 285.950 1400.140 286.270 ;
        RECT 1450.940 285.950 1451.200 286.270 ;
        RECT 1399.940 17.410 1400.080 285.950 ;
        RECT 1399.940 17.270 1400.540 17.410 ;
        RECT 1400.400 2.400 1400.540 17.270 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1421.010 288.560 1421.330 288.620 ;
        RECT 1465.170 288.560 1465.490 288.620 ;
        RECT 1421.010 288.420 1465.490 288.560 ;
        RECT 1421.010 288.360 1421.330 288.420 ;
        RECT 1465.170 288.360 1465.490 288.420 ;
        RECT 1418.250 17.580 1418.570 17.640 ;
        RECT 1421.010 17.580 1421.330 17.640 ;
        RECT 1418.250 17.440 1421.330 17.580 ;
        RECT 1418.250 17.380 1418.570 17.440 ;
        RECT 1421.010 17.380 1421.330 17.440 ;
      LAYER via ;
        RECT 1421.040 288.360 1421.300 288.620 ;
        RECT 1465.200 288.360 1465.460 288.620 ;
        RECT 1418.280 17.380 1418.540 17.640 ;
        RECT 1421.040 17.380 1421.300 17.640 ;
      LAYER met2 ;
        RECT 1465.200 300.000 1465.480 304.000 ;
        RECT 1465.260 288.650 1465.400 300.000 ;
        RECT 1421.040 288.330 1421.300 288.650 ;
        RECT 1465.200 288.330 1465.460 288.650 ;
        RECT 1421.100 17.670 1421.240 288.330 ;
        RECT 1418.280 17.350 1418.540 17.670 ;
        RECT 1421.040 17.350 1421.300 17.670 ;
        RECT 1418.340 2.400 1418.480 17.350 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1441.710 284.820 1442.030 284.880 ;
        RECT 1479.890 284.820 1480.210 284.880 ;
        RECT 1441.710 284.680 1480.210 284.820 ;
        RECT 1441.710 284.620 1442.030 284.680 ;
        RECT 1479.890 284.620 1480.210 284.680 ;
        RECT 1435.730 17.920 1436.050 17.980 ;
        RECT 1441.710 17.920 1442.030 17.980 ;
        RECT 1435.730 17.780 1442.030 17.920 ;
        RECT 1435.730 17.720 1436.050 17.780 ;
        RECT 1441.710 17.720 1442.030 17.780 ;
      LAYER via ;
        RECT 1441.740 284.620 1442.000 284.880 ;
        RECT 1479.920 284.620 1480.180 284.880 ;
        RECT 1435.760 17.720 1436.020 17.980 ;
        RECT 1441.740 17.720 1442.000 17.980 ;
      LAYER met2 ;
        RECT 1479.920 300.000 1480.200 304.000 ;
        RECT 1479.980 284.910 1480.120 300.000 ;
        RECT 1441.740 284.590 1442.000 284.910 ;
        RECT 1479.920 284.590 1480.180 284.910 ;
        RECT 1441.800 18.010 1441.940 284.590 ;
        RECT 1435.760 17.690 1436.020 18.010 ;
        RECT 1441.740 17.690 1442.000 18.010 ;
        RECT 1435.820 2.400 1435.960 17.690 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1455.510 283.120 1455.830 283.180 ;
        RECT 1494.610 283.120 1494.930 283.180 ;
        RECT 1455.510 282.980 1494.930 283.120 ;
        RECT 1455.510 282.920 1455.830 282.980 ;
        RECT 1494.610 282.920 1494.930 282.980 ;
      LAYER via ;
        RECT 1455.540 282.920 1455.800 283.180 ;
        RECT 1494.640 282.920 1494.900 283.180 ;
      LAYER met2 ;
        RECT 1494.640 300.000 1494.920 304.000 ;
        RECT 1494.700 283.210 1494.840 300.000 ;
        RECT 1455.540 282.890 1455.800 283.210 ;
        RECT 1494.640 282.890 1494.900 283.210 ;
        RECT 1455.600 17.410 1455.740 282.890 ;
        RECT 1453.760 17.270 1455.740 17.410 ;
        RECT 1453.760 2.400 1453.900 17.270 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1476.210 286.860 1476.530 286.920 ;
        RECT 1509.330 286.860 1509.650 286.920 ;
        RECT 1476.210 286.720 1509.650 286.860 ;
        RECT 1476.210 286.660 1476.530 286.720 ;
        RECT 1509.330 286.660 1509.650 286.720 ;
        RECT 1471.610 17.580 1471.930 17.640 ;
        RECT 1476.210 17.580 1476.530 17.640 ;
        RECT 1471.610 17.440 1476.530 17.580 ;
        RECT 1471.610 17.380 1471.930 17.440 ;
        RECT 1476.210 17.380 1476.530 17.440 ;
      LAYER via ;
        RECT 1476.240 286.660 1476.500 286.920 ;
        RECT 1509.360 286.660 1509.620 286.920 ;
        RECT 1471.640 17.380 1471.900 17.640 ;
        RECT 1476.240 17.380 1476.500 17.640 ;
      LAYER met2 ;
        RECT 1509.360 300.000 1509.640 304.000 ;
        RECT 1509.420 286.950 1509.560 300.000 ;
        RECT 1476.240 286.630 1476.500 286.950 ;
        RECT 1509.360 286.630 1509.620 286.950 ;
        RECT 1476.300 17.670 1476.440 286.630 ;
        RECT 1471.640 17.350 1471.900 17.670 ;
        RECT 1476.240 17.350 1476.500 17.670 ;
        RECT 1471.700 2.400 1471.840 17.350 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1490.010 286.520 1490.330 286.580 ;
        RECT 1524.050 286.520 1524.370 286.580 ;
        RECT 1490.010 286.380 1524.370 286.520 ;
        RECT 1490.010 286.320 1490.330 286.380 ;
        RECT 1524.050 286.320 1524.370 286.380 ;
      LAYER via ;
        RECT 1490.040 286.320 1490.300 286.580 ;
        RECT 1524.080 286.320 1524.340 286.580 ;
      LAYER met2 ;
        RECT 1524.080 300.000 1524.360 304.000 ;
        RECT 1524.140 286.610 1524.280 300.000 ;
        RECT 1490.040 286.290 1490.300 286.610 ;
        RECT 1524.080 286.290 1524.340 286.610 ;
        RECT 1490.100 17.410 1490.240 286.290 ;
        RECT 1489.640 17.270 1490.240 17.410 ;
        RECT 1489.640 2.400 1489.780 17.270 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1510.710 283.800 1511.030 283.860 ;
        RECT 1538.770 283.800 1539.090 283.860 ;
        RECT 1510.710 283.660 1539.090 283.800 ;
        RECT 1510.710 283.600 1511.030 283.660 ;
        RECT 1538.770 283.600 1539.090 283.660 ;
        RECT 1507.030 17.580 1507.350 17.640 ;
        RECT 1510.710 17.580 1511.030 17.640 ;
        RECT 1507.030 17.440 1511.030 17.580 ;
        RECT 1507.030 17.380 1507.350 17.440 ;
        RECT 1510.710 17.380 1511.030 17.440 ;
      LAYER via ;
        RECT 1510.740 283.600 1511.000 283.860 ;
        RECT 1538.800 283.600 1539.060 283.860 ;
        RECT 1507.060 17.380 1507.320 17.640 ;
        RECT 1510.740 17.380 1511.000 17.640 ;
      LAYER met2 ;
        RECT 1538.800 300.000 1539.080 304.000 ;
        RECT 1538.860 283.890 1539.000 300.000 ;
        RECT 1510.740 283.570 1511.000 283.890 ;
        RECT 1538.800 283.570 1539.060 283.890 ;
        RECT 1510.800 17.670 1510.940 283.570 ;
        RECT 1507.060 17.350 1507.320 17.670 ;
        RECT 1510.740 17.350 1511.000 17.670 ;
        RECT 1507.120 2.400 1507.260 17.350 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 727.880 20.840 731.700 20.980 ;
        RECT 704.330 20.640 704.650 20.700 ;
        RECT 727.880 20.640 728.020 20.840 ;
        RECT 704.330 20.500 728.020 20.640 ;
        RECT 731.560 20.640 731.700 20.840 ;
        RECT 876.830 20.640 877.150 20.700 ;
        RECT 731.560 20.500 877.150 20.640 ;
        RECT 704.330 20.440 704.650 20.500 ;
        RECT 876.830 20.440 877.150 20.500 ;
      LAYER via ;
        RECT 704.360 20.440 704.620 20.700 ;
        RECT 876.860 20.440 877.120 20.700 ;
      LAYER met2 ;
        RECT 877.780 300.290 878.060 304.000 ;
        RECT 876.920 300.150 878.060 300.290 ;
        RECT 876.920 20.730 877.060 300.150 ;
        RECT 877.780 300.000 878.060 300.150 ;
        RECT 704.360 20.410 704.620 20.730 ;
        RECT 876.860 20.410 877.120 20.730 ;
        RECT 704.420 2.400 704.560 20.410 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1530.950 286.520 1531.270 286.580 ;
        RECT 1553.490 286.520 1553.810 286.580 ;
        RECT 1530.950 286.380 1553.810 286.520 ;
        RECT 1530.950 286.320 1531.270 286.380 ;
        RECT 1553.490 286.320 1553.810 286.380 ;
        RECT 1524.970 17.920 1525.290 17.980 ;
        RECT 1530.950 17.920 1531.270 17.980 ;
        RECT 1524.970 17.780 1531.270 17.920 ;
        RECT 1524.970 17.720 1525.290 17.780 ;
        RECT 1530.950 17.720 1531.270 17.780 ;
      LAYER via ;
        RECT 1530.980 286.320 1531.240 286.580 ;
        RECT 1553.520 286.320 1553.780 286.580 ;
        RECT 1525.000 17.720 1525.260 17.980 ;
        RECT 1530.980 17.720 1531.240 17.980 ;
      LAYER met2 ;
        RECT 1553.520 300.000 1553.800 304.000 ;
        RECT 1553.580 286.610 1553.720 300.000 ;
        RECT 1530.980 286.290 1531.240 286.610 ;
        RECT 1553.520 286.290 1553.780 286.610 ;
        RECT 1531.040 18.010 1531.180 286.290 ;
        RECT 1525.000 17.690 1525.260 18.010 ;
        RECT 1530.980 17.690 1531.240 18.010 ;
        RECT 1525.060 2.400 1525.200 17.690 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1545.210 287.880 1545.530 287.940 ;
        RECT 1568.210 287.880 1568.530 287.940 ;
        RECT 1545.210 287.740 1568.530 287.880 ;
        RECT 1545.210 287.680 1545.530 287.740 ;
        RECT 1568.210 287.680 1568.530 287.740 ;
        RECT 1542.910 17.580 1543.230 17.640 ;
        RECT 1545.210 17.580 1545.530 17.640 ;
        RECT 1542.910 17.440 1545.530 17.580 ;
        RECT 1542.910 17.380 1543.230 17.440 ;
        RECT 1545.210 17.380 1545.530 17.440 ;
      LAYER via ;
        RECT 1545.240 287.680 1545.500 287.940 ;
        RECT 1568.240 287.680 1568.500 287.940 ;
        RECT 1542.940 17.380 1543.200 17.640 ;
        RECT 1545.240 17.380 1545.500 17.640 ;
      LAYER met2 ;
        RECT 1568.240 300.000 1568.520 304.000 ;
        RECT 1568.300 287.970 1568.440 300.000 ;
        RECT 1545.240 287.650 1545.500 287.970 ;
        RECT 1568.240 287.650 1568.500 287.970 ;
        RECT 1545.300 17.670 1545.440 287.650 ;
        RECT 1542.940 17.350 1543.200 17.670 ;
        RECT 1545.240 17.350 1545.500 17.670 ;
        RECT 1543.000 2.400 1543.140 17.350 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1565.910 283.800 1566.230 283.860 ;
        RECT 1582.930 283.800 1583.250 283.860 ;
        RECT 1565.910 283.660 1583.250 283.800 ;
        RECT 1565.910 283.600 1566.230 283.660 ;
        RECT 1582.930 283.600 1583.250 283.660 ;
        RECT 1560.850 17.580 1561.170 17.640 ;
        RECT 1565.910 17.580 1566.230 17.640 ;
        RECT 1560.850 17.440 1566.230 17.580 ;
        RECT 1560.850 17.380 1561.170 17.440 ;
        RECT 1565.910 17.380 1566.230 17.440 ;
      LAYER via ;
        RECT 1565.940 283.600 1566.200 283.860 ;
        RECT 1582.960 283.600 1583.220 283.860 ;
        RECT 1560.880 17.380 1561.140 17.640 ;
        RECT 1565.940 17.380 1566.200 17.640 ;
      LAYER met2 ;
        RECT 1582.960 300.000 1583.240 304.000 ;
        RECT 1583.020 283.890 1583.160 300.000 ;
        RECT 1565.940 283.570 1566.200 283.890 ;
        RECT 1582.960 283.570 1583.220 283.890 ;
        RECT 1566.000 17.670 1566.140 283.570 ;
        RECT 1560.880 17.350 1561.140 17.670 ;
        RECT 1565.940 17.350 1566.200 17.670 ;
        RECT 1560.940 2.400 1561.080 17.350 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1579.710 286.180 1580.030 286.240 ;
        RECT 1597.650 286.180 1597.970 286.240 ;
        RECT 1579.710 286.040 1597.970 286.180 ;
        RECT 1579.710 285.980 1580.030 286.040 ;
        RECT 1597.650 285.980 1597.970 286.040 ;
      LAYER via ;
        RECT 1579.740 285.980 1580.000 286.240 ;
        RECT 1597.680 285.980 1597.940 286.240 ;
      LAYER met2 ;
        RECT 1597.680 300.000 1597.960 304.000 ;
        RECT 1597.740 286.270 1597.880 300.000 ;
        RECT 1579.740 285.950 1580.000 286.270 ;
        RECT 1597.680 285.950 1597.940 286.270 ;
        RECT 1579.800 17.410 1579.940 285.950 ;
        RECT 1578.880 17.270 1579.940 17.410 ;
        RECT 1578.880 2.400 1579.020 17.270 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1600.410 287.540 1600.730 287.600 ;
        RECT 1612.370 287.540 1612.690 287.600 ;
        RECT 1600.410 287.400 1612.690 287.540 ;
        RECT 1600.410 287.340 1600.730 287.400 ;
        RECT 1612.370 287.340 1612.690 287.400 ;
        RECT 1596.270 17.240 1596.590 17.300 ;
        RECT 1600.410 17.240 1600.730 17.300 ;
        RECT 1596.270 17.100 1600.730 17.240 ;
        RECT 1596.270 17.040 1596.590 17.100 ;
        RECT 1600.410 17.040 1600.730 17.100 ;
      LAYER via ;
        RECT 1600.440 287.340 1600.700 287.600 ;
        RECT 1612.400 287.340 1612.660 287.600 ;
        RECT 1596.300 17.040 1596.560 17.300 ;
        RECT 1600.440 17.040 1600.700 17.300 ;
      LAYER met2 ;
        RECT 1612.400 300.000 1612.680 304.000 ;
        RECT 1612.460 287.630 1612.600 300.000 ;
        RECT 1600.440 287.310 1600.700 287.630 ;
        RECT 1612.400 287.310 1612.660 287.630 ;
        RECT 1600.500 17.330 1600.640 287.310 ;
        RECT 1596.300 17.010 1596.560 17.330 ;
        RECT 1600.440 17.010 1600.700 17.330 ;
        RECT 1596.360 2.400 1596.500 17.010 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1614.210 288.220 1614.530 288.280 ;
        RECT 1627.090 288.220 1627.410 288.280 ;
        RECT 1614.210 288.080 1627.410 288.220 ;
        RECT 1614.210 288.020 1614.530 288.080 ;
        RECT 1627.090 288.020 1627.410 288.080 ;
      LAYER via ;
        RECT 1614.240 288.020 1614.500 288.280 ;
        RECT 1627.120 288.020 1627.380 288.280 ;
      LAYER met2 ;
        RECT 1627.120 300.000 1627.400 304.000 ;
        RECT 1627.180 288.310 1627.320 300.000 ;
        RECT 1614.240 287.990 1614.500 288.310 ;
        RECT 1627.120 287.990 1627.380 288.310 ;
        RECT 1614.300 2.400 1614.440 287.990 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1634.910 288.900 1635.230 288.960 ;
        RECT 1641.810 288.900 1642.130 288.960 ;
        RECT 1634.910 288.760 1642.130 288.900 ;
        RECT 1634.910 288.700 1635.230 288.760 ;
        RECT 1641.810 288.700 1642.130 288.760 ;
        RECT 1632.150 17.580 1632.470 17.640 ;
        RECT 1634.910 17.580 1635.230 17.640 ;
        RECT 1632.150 17.440 1635.230 17.580 ;
        RECT 1632.150 17.380 1632.470 17.440 ;
        RECT 1634.910 17.380 1635.230 17.440 ;
      LAYER via ;
        RECT 1634.940 288.700 1635.200 288.960 ;
        RECT 1641.840 288.700 1642.100 288.960 ;
        RECT 1632.180 17.380 1632.440 17.640 ;
        RECT 1634.940 17.380 1635.200 17.640 ;
      LAYER met2 ;
        RECT 1641.840 300.000 1642.120 304.000 ;
        RECT 1641.900 288.990 1642.040 300.000 ;
        RECT 1634.940 288.670 1635.200 288.990 ;
        RECT 1641.840 288.670 1642.100 288.990 ;
        RECT 1635.000 17.670 1635.140 288.670 ;
        RECT 1632.180 17.350 1632.440 17.670 ;
        RECT 1634.940 17.350 1635.200 17.670 ;
        RECT 1632.240 2.400 1632.380 17.350 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1650.090 16.560 1650.410 16.620 ;
        RECT 1655.610 16.560 1655.930 16.620 ;
        RECT 1650.090 16.420 1655.930 16.560 ;
        RECT 1650.090 16.360 1650.410 16.420 ;
        RECT 1655.610 16.360 1655.930 16.420 ;
      LAYER via ;
        RECT 1650.120 16.360 1650.380 16.620 ;
        RECT 1655.640 16.360 1655.900 16.620 ;
      LAYER met2 ;
        RECT 1656.560 300.290 1656.840 304.000 ;
        RECT 1656.160 300.150 1656.840 300.290 ;
        RECT 1656.160 288.050 1656.300 300.150 ;
        RECT 1656.560 300.000 1656.840 300.150 ;
        RECT 1655.700 287.910 1656.300 288.050 ;
        RECT 1655.700 16.650 1655.840 287.910 ;
        RECT 1650.120 16.330 1650.380 16.650 ;
        RECT 1655.640 16.330 1655.900 16.650 ;
        RECT 1650.180 2.400 1650.320 16.330 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1668.105 2.805 1668.275 14.195 ;
      LAYER mcon ;
        RECT 1668.105 14.025 1668.275 14.195 ;
      LAYER met1 ;
        RECT 1668.045 14.180 1668.335 14.225 ;
        RECT 1669.410 14.180 1669.730 14.240 ;
        RECT 1668.045 14.040 1669.730 14.180 ;
        RECT 1668.045 13.995 1668.335 14.040 ;
        RECT 1669.410 13.980 1669.730 14.040 ;
        RECT 1668.030 2.960 1668.350 3.020 ;
        RECT 1667.835 2.820 1668.350 2.960 ;
        RECT 1668.030 2.760 1668.350 2.820 ;
      LAYER via ;
        RECT 1669.440 13.980 1669.700 14.240 ;
        RECT 1668.060 2.760 1668.320 3.020 ;
      LAYER met2 ;
        RECT 1671.280 300.290 1671.560 304.000 ;
        RECT 1669.960 300.150 1671.560 300.290 ;
        RECT 1669.960 283.290 1670.100 300.150 ;
        RECT 1671.280 300.000 1671.560 300.150 ;
        RECT 1669.500 283.150 1670.100 283.290 ;
        RECT 1669.500 14.270 1669.640 283.150 ;
        RECT 1669.440 13.950 1669.700 14.270 ;
        RECT 1668.060 2.730 1668.320 3.050 ;
        RECT 1668.120 2.400 1668.260 2.730 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1683.745 234.685 1683.915 282.455 ;
        RECT 1683.745 138.125 1683.915 186.235 ;
        RECT 1683.745 47.685 1683.915 89.675 ;
      LAYER mcon ;
        RECT 1683.745 282.285 1683.915 282.455 ;
        RECT 1683.745 186.065 1683.915 186.235 ;
        RECT 1683.745 89.505 1683.915 89.675 ;
      LAYER met1 ;
        RECT 1683.670 283.120 1683.990 283.180 ;
        RECT 1685.970 283.120 1686.290 283.180 ;
        RECT 1683.670 282.980 1686.290 283.120 ;
        RECT 1683.670 282.920 1683.990 282.980 ;
        RECT 1685.970 282.920 1686.290 282.980 ;
        RECT 1683.670 282.440 1683.990 282.500 ;
        RECT 1683.670 282.300 1684.185 282.440 ;
        RECT 1683.670 282.240 1683.990 282.300 ;
        RECT 1683.670 234.840 1683.990 234.900 ;
        RECT 1683.670 234.700 1684.185 234.840 ;
        RECT 1683.670 234.640 1683.990 234.700 ;
        RECT 1683.670 186.220 1683.990 186.280 ;
        RECT 1683.670 186.080 1684.185 186.220 ;
        RECT 1683.670 186.020 1683.990 186.080 ;
        RECT 1683.670 138.280 1683.990 138.340 ;
        RECT 1683.670 138.140 1684.185 138.280 ;
        RECT 1683.670 138.080 1683.990 138.140 ;
        RECT 1683.670 89.660 1683.990 89.720 ;
        RECT 1683.670 89.520 1684.185 89.660 ;
        RECT 1683.670 89.460 1683.990 89.520 ;
        RECT 1683.685 47.840 1683.975 47.885 ;
        RECT 1685.510 47.840 1685.830 47.900 ;
        RECT 1683.685 47.700 1685.830 47.840 ;
        RECT 1683.685 47.655 1683.975 47.700 ;
        RECT 1685.510 47.640 1685.830 47.700 ;
      LAYER via ;
        RECT 1683.700 282.920 1683.960 283.180 ;
        RECT 1686.000 282.920 1686.260 283.180 ;
        RECT 1683.700 282.240 1683.960 282.500 ;
        RECT 1683.700 234.640 1683.960 234.900 ;
        RECT 1683.700 186.020 1683.960 186.280 ;
        RECT 1683.700 138.080 1683.960 138.340 ;
        RECT 1683.700 89.460 1683.960 89.720 ;
        RECT 1685.540 47.640 1685.800 47.900 ;
      LAYER met2 ;
        RECT 1686.000 300.000 1686.280 304.000 ;
        RECT 1686.060 283.210 1686.200 300.000 ;
        RECT 1683.700 282.890 1683.960 283.210 ;
        RECT 1686.000 282.890 1686.260 283.210 ;
        RECT 1683.760 282.530 1683.900 282.890 ;
        RECT 1683.700 282.210 1683.960 282.530 ;
        RECT 1683.700 234.610 1683.960 234.930 ;
        RECT 1683.760 186.310 1683.900 234.610 ;
        RECT 1683.700 185.990 1683.960 186.310 ;
        RECT 1683.700 138.050 1683.960 138.370 ;
        RECT 1683.760 90.850 1683.900 138.050 ;
        RECT 1683.760 90.710 1684.360 90.850 ;
        RECT 1684.220 90.170 1684.360 90.710 ;
        RECT 1683.760 90.030 1684.360 90.170 ;
        RECT 1683.760 89.750 1683.900 90.030 ;
        RECT 1683.700 89.430 1683.960 89.750 ;
        RECT 1685.540 47.610 1685.800 47.930 ;
        RECT 1685.600 2.400 1685.740 47.610 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 722.270 20.300 722.590 20.360 ;
        RECT 890.170 20.300 890.490 20.360 ;
        RECT 722.270 20.160 890.490 20.300 ;
        RECT 722.270 20.100 722.590 20.160 ;
        RECT 890.170 20.100 890.490 20.160 ;
      LAYER via ;
        RECT 722.300 20.100 722.560 20.360 ;
        RECT 890.200 20.100 890.460 20.360 ;
      LAYER met2 ;
        RECT 892.500 300.290 892.780 304.000 ;
        RECT 890.260 300.150 892.780 300.290 ;
        RECT 890.260 20.390 890.400 300.150 ;
        RECT 892.500 300.000 892.780 300.150 ;
        RECT 722.300 20.070 722.560 20.390 ;
        RECT 890.200 20.070 890.460 20.390 ;
        RECT 722.360 2.400 722.500 20.070 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1697.470 20.640 1697.790 20.700 ;
        RECT 1703.450 20.640 1703.770 20.700 ;
        RECT 1697.470 20.500 1703.770 20.640 ;
        RECT 1697.470 20.440 1697.790 20.500 ;
        RECT 1703.450 20.440 1703.770 20.500 ;
      LAYER via ;
        RECT 1697.500 20.440 1697.760 20.700 ;
        RECT 1703.480 20.440 1703.740 20.700 ;
      LAYER met2 ;
        RECT 1700.720 300.290 1701.000 304.000 ;
        RECT 1697.560 300.150 1701.000 300.290 ;
        RECT 1697.560 20.730 1697.700 300.150 ;
        RECT 1700.720 300.000 1701.000 300.150 ;
        RECT 1697.500 20.410 1697.760 20.730 ;
        RECT 1703.480 20.410 1703.740 20.730 ;
        RECT 1703.540 2.400 1703.680 20.410 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1714.950 283.460 1715.270 283.520 ;
        RECT 1718.630 283.460 1718.950 283.520 ;
        RECT 1714.950 283.320 1718.950 283.460 ;
        RECT 1714.950 283.260 1715.270 283.320 ;
        RECT 1718.630 283.260 1718.950 283.320 ;
      LAYER via ;
        RECT 1714.980 283.260 1715.240 283.520 ;
        RECT 1718.660 283.260 1718.920 283.520 ;
      LAYER met2 ;
        RECT 1714.980 300.000 1715.260 304.000 ;
        RECT 1715.040 283.550 1715.180 300.000 ;
        RECT 1714.980 283.230 1715.240 283.550 ;
        RECT 1718.660 283.230 1718.920 283.550 ;
        RECT 1718.720 17.410 1718.860 283.230 ;
        RECT 1718.720 17.270 1721.620 17.410 ;
        RECT 1721.480 2.400 1721.620 17.270 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1731.050 17.240 1731.370 17.300 ;
        RECT 1739.330 17.240 1739.650 17.300 ;
        RECT 1731.050 17.100 1739.650 17.240 ;
        RECT 1731.050 17.040 1731.370 17.100 ;
        RECT 1739.330 17.040 1739.650 17.100 ;
      LAYER via ;
        RECT 1731.080 17.040 1731.340 17.300 ;
        RECT 1739.360 17.040 1739.620 17.300 ;
      LAYER met2 ;
        RECT 1729.700 300.290 1729.980 304.000 ;
        RECT 1729.700 300.150 1731.280 300.290 ;
        RECT 1729.700 300.000 1729.980 300.150 ;
        RECT 1731.140 17.330 1731.280 300.150 ;
        RECT 1731.080 17.010 1731.340 17.330 ;
        RECT 1739.360 17.010 1739.620 17.330 ;
        RECT 1739.420 2.400 1739.560 17.010 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1744.850 17.920 1745.170 17.980 ;
        RECT 1756.810 17.920 1757.130 17.980 ;
        RECT 1744.850 17.780 1757.130 17.920 ;
        RECT 1744.850 17.720 1745.170 17.780 ;
        RECT 1756.810 17.720 1757.130 17.780 ;
      LAYER via ;
        RECT 1744.880 17.720 1745.140 17.980 ;
        RECT 1756.840 17.720 1757.100 17.980 ;
      LAYER met2 ;
        RECT 1744.420 300.290 1744.700 304.000 ;
        RECT 1744.420 300.150 1745.080 300.290 ;
        RECT 1744.420 300.000 1744.700 300.150 ;
        RECT 1744.940 18.010 1745.080 300.150 ;
        RECT 1744.880 17.690 1745.140 18.010 ;
        RECT 1756.840 17.690 1757.100 18.010 ;
        RECT 1756.900 2.400 1757.040 17.690 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1758.650 17.920 1758.970 17.980 ;
        RECT 1774.750 17.920 1775.070 17.980 ;
        RECT 1758.650 17.780 1775.070 17.920 ;
        RECT 1758.650 17.720 1758.970 17.780 ;
        RECT 1774.750 17.720 1775.070 17.780 ;
      LAYER via ;
        RECT 1758.680 17.720 1758.940 17.980 ;
        RECT 1774.780 17.720 1775.040 17.980 ;
      LAYER met2 ;
        RECT 1759.140 300.290 1759.420 304.000 ;
        RECT 1758.740 300.150 1759.420 300.290 ;
        RECT 1758.740 18.010 1758.880 300.150 ;
        RECT 1759.140 300.000 1759.420 300.150 ;
        RECT 1758.680 17.690 1758.940 18.010 ;
        RECT 1774.780 17.690 1775.040 18.010 ;
        RECT 1774.840 2.400 1774.980 17.690 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1773.830 286.180 1774.150 286.240 ;
        RECT 1779.350 286.180 1779.670 286.240 ;
        RECT 1773.830 286.040 1779.670 286.180 ;
        RECT 1773.830 285.980 1774.150 286.040 ;
        RECT 1779.350 285.980 1779.670 286.040 ;
        RECT 1779.350 15.880 1779.670 15.940 ;
        RECT 1792.690 15.880 1793.010 15.940 ;
        RECT 1779.350 15.740 1793.010 15.880 ;
        RECT 1779.350 15.680 1779.670 15.740 ;
        RECT 1792.690 15.680 1793.010 15.740 ;
      LAYER via ;
        RECT 1773.860 285.980 1774.120 286.240 ;
        RECT 1779.380 285.980 1779.640 286.240 ;
        RECT 1779.380 15.680 1779.640 15.940 ;
        RECT 1792.720 15.680 1792.980 15.940 ;
      LAYER met2 ;
        RECT 1773.860 300.000 1774.140 304.000 ;
        RECT 1773.920 286.270 1774.060 300.000 ;
        RECT 1773.860 285.950 1774.120 286.270 ;
        RECT 1779.380 285.950 1779.640 286.270 ;
        RECT 1779.440 15.970 1779.580 285.950 ;
        RECT 1779.380 15.650 1779.640 15.970 ;
        RECT 1792.720 15.650 1792.980 15.970 ;
        RECT 1792.780 2.400 1792.920 15.650 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1788.550 288.220 1788.870 288.280 ;
        RECT 1793.150 288.220 1793.470 288.280 ;
        RECT 1788.550 288.080 1793.470 288.220 ;
        RECT 1788.550 288.020 1788.870 288.080 ;
        RECT 1793.150 288.020 1793.470 288.080 ;
        RECT 1793.150 16.560 1793.470 16.620 ;
        RECT 1810.630 16.560 1810.950 16.620 ;
        RECT 1793.150 16.420 1810.950 16.560 ;
        RECT 1793.150 16.360 1793.470 16.420 ;
        RECT 1810.630 16.360 1810.950 16.420 ;
      LAYER via ;
        RECT 1788.580 288.020 1788.840 288.280 ;
        RECT 1793.180 288.020 1793.440 288.280 ;
        RECT 1793.180 16.360 1793.440 16.620 ;
        RECT 1810.660 16.360 1810.920 16.620 ;
      LAYER met2 ;
        RECT 1788.580 300.000 1788.860 304.000 ;
        RECT 1788.640 288.310 1788.780 300.000 ;
        RECT 1788.580 287.990 1788.840 288.310 ;
        RECT 1793.180 287.990 1793.440 288.310 ;
        RECT 1793.240 16.650 1793.380 287.990 ;
        RECT 1793.180 16.330 1793.440 16.650 ;
        RECT 1810.660 16.330 1810.920 16.650 ;
        RECT 1810.720 2.400 1810.860 16.330 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1803.270 288.220 1803.590 288.280 ;
        RECT 1811.090 288.220 1811.410 288.280 ;
        RECT 1803.270 288.080 1811.410 288.220 ;
        RECT 1803.270 288.020 1803.590 288.080 ;
        RECT 1811.090 288.020 1811.410 288.080 ;
        RECT 1811.090 20.640 1811.410 20.700 ;
        RECT 1828.570 20.640 1828.890 20.700 ;
        RECT 1811.090 20.500 1828.890 20.640 ;
        RECT 1811.090 20.440 1811.410 20.500 ;
        RECT 1828.570 20.440 1828.890 20.500 ;
      LAYER via ;
        RECT 1803.300 288.020 1803.560 288.280 ;
        RECT 1811.120 288.020 1811.380 288.280 ;
        RECT 1811.120 20.440 1811.380 20.700 ;
        RECT 1828.600 20.440 1828.860 20.700 ;
      LAYER met2 ;
        RECT 1803.300 300.000 1803.580 304.000 ;
        RECT 1803.360 288.310 1803.500 300.000 ;
        RECT 1803.300 287.990 1803.560 288.310 ;
        RECT 1811.120 287.990 1811.380 288.310 ;
        RECT 1811.180 20.730 1811.320 287.990 ;
        RECT 1811.120 20.410 1811.380 20.730 ;
        RECT 1828.600 20.410 1828.860 20.730 ;
        RECT 1828.660 2.400 1828.800 20.410 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1821.210 18.600 1821.530 18.660 ;
        RECT 1846.050 18.600 1846.370 18.660 ;
        RECT 1821.210 18.460 1846.370 18.600 ;
        RECT 1821.210 18.400 1821.530 18.460 ;
        RECT 1846.050 18.400 1846.370 18.460 ;
      LAYER via ;
        RECT 1821.240 18.400 1821.500 18.660 ;
        RECT 1846.080 18.400 1846.340 18.660 ;
      LAYER met2 ;
        RECT 1818.020 300.290 1818.300 304.000 ;
        RECT 1818.020 300.150 1821.440 300.290 ;
        RECT 1818.020 300.000 1818.300 300.150 ;
        RECT 1821.300 18.690 1821.440 300.150 ;
        RECT 1821.240 18.370 1821.500 18.690 ;
        RECT 1846.080 18.370 1846.340 18.690 ;
        RECT 1846.140 2.400 1846.280 18.370 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1835.010 17.580 1835.330 17.640 ;
        RECT 1863.990 17.580 1864.310 17.640 ;
        RECT 1835.010 17.440 1864.310 17.580 ;
        RECT 1835.010 17.380 1835.330 17.440 ;
        RECT 1863.990 17.380 1864.310 17.440 ;
      LAYER via ;
        RECT 1835.040 17.380 1835.300 17.640 ;
        RECT 1864.020 17.380 1864.280 17.640 ;
      LAYER met2 ;
        RECT 1832.740 300.290 1833.020 304.000 ;
        RECT 1832.740 300.150 1835.240 300.290 ;
        RECT 1832.740 300.000 1833.020 300.150 ;
        RECT 1835.100 17.670 1835.240 300.150 ;
        RECT 1835.040 17.350 1835.300 17.670 ;
        RECT 1864.020 17.350 1864.280 17.670 ;
        RECT 1864.080 2.400 1864.220 17.350 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 740.210 25.740 740.530 25.800 ;
        RECT 903.970 25.740 904.290 25.800 ;
        RECT 740.210 25.600 904.290 25.740 ;
        RECT 740.210 25.540 740.530 25.600 ;
        RECT 903.970 25.540 904.290 25.600 ;
      LAYER via ;
        RECT 740.240 25.540 740.500 25.800 ;
        RECT 904.000 25.540 904.260 25.800 ;
      LAYER met2 ;
        RECT 907.220 300.290 907.500 304.000 ;
        RECT 904.060 300.150 907.500 300.290 ;
        RECT 904.060 25.830 904.200 300.150 ;
        RECT 907.220 300.000 907.500 300.150 ;
        RECT 740.240 25.510 740.500 25.830 ;
        RECT 904.000 25.510 904.260 25.830 ;
        RECT 740.300 2.400 740.440 25.510 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1848.810 19.280 1849.130 19.340 ;
        RECT 1881.930 19.280 1882.250 19.340 ;
        RECT 1848.810 19.140 1882.250 19.280 ;
        RECT 1848.810 19.080 1849.130 19.140 ;
        RECT 1881.930 19.080 1882.250 19.140 ;
      LAYER via ;
        RECT 1848.840 19.080 1849.100 19.340 ;
        RECT 1881.960 19.080 1882.220 19.340 ;
      LAYER met2 ;
        RECT 1847.460 300.290 1847.740 304.000 ;
        RECT 1847.460 300.150 1849.040 300.290 ;
        RECT 1847.460 300.000 1847.740 300.150 ;
        RECT 1848.900 19.370 1849.040 300.150 ;
        RECT 1848.840 19.050 1849.100 19.370 ;
        RECT 1881.960 19.050 1882.220 19.370 ;
        RECT 1882.020 2.400 1882.160 19.050 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1862.610 17.240 1862.930 17.300 ;
        RECT 1899.870 17.240 1900.190 17.300 ;
        RECT 1862.610 17.100 1900.190 17.240 ;
        RECT 1862.610 17.040 1862.930 17.100 ;
        RECT 1899.870 17.040 1900.190 17.100 ;
      LAYER via ;
        RECT 1862.640 17.040 1862.900 17.300 ;
        RECT 1899.900 17.040 1900.160 17.300 ;
      LAYER met2 ;
        RECT 1862.180 300.290 1862.460 304.000 ;
        RECT 1862.180 300.150 1862.840 300.290 ;
        RECT 1862.180 300.000 1862.460 300.150 ;
        RECT 1862.700 17.330 1862.840 300.150 ;
        RECT 1862.640 17.010 1862.900 17.330 ;
        RECT 1899.900 17.010 1900.160 17.330 ;
        RECT 1899.960 2.400 1900.100 17.010 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1876.870 288.220 1877.190 288.280 ;
        RECT 1882.850 288.220 1883.170 288.280 ;
        RECT 1876.870 288.080 1883.170 288.220 ;
        RECT 1876.870 288.020 1877.190 288.080 ;
        RECT 1882.850 288.020 1883.170 288.080 ;
        RECT 1882.850 16.220 1883.170 16.280 ;
        RECT 1917.810 16.220 1918.130 16.280 ;
        RECT 1882.850 16.080 1918.130 16.220 ;
        RECT 1882.850 16.020 1883.170 16.080 ;
        RECT 1917.810 16.020 1918.130 16.080 ;
      LAYER via ;
        RECT 1876.900 288.020 1877.160 288.280 ;
        RECT 1882.880 288.020 1883.140 288.280 ;
        RECT 1882.880 16.020 1883.140 16.280 ;
        RECT 1917.840 16.020 1918.100 16.280 ;
      LAYER met2 ;
        RECT 1876.900 300.000 1877.180 304.000 ;
        RECT 1876.960 288.310 1877.100 300.000 ;
        RECT 1876.900 287.990 1877.160 288.310 ;
        RECT 1882.880 287.990 1883.140 288.310 ;
        RECT 1882.940 16.310 1883.080 287.990 ;
        RECT 1882.880 15.990 1883.140 16.310 ;
        RECT 1917.840 15.990 1918.100 16.310 ;
        RECT 1917.900 2.400 1918.040 15.990 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1891.590 287.880 1891.910 287.940 ;
        RECT 1897.110 287.880 1897.430 287.940 ;
        RECT 1891.590 287.740 1897.430 287.880 ;
        RECT 1891.590 287.680 1891.910 287.740 ;
        RECT 1897.110 287.680 1897.430 287.740 ;
        RECT 1897.110 20.640 1897.430 20.700 ;
        RECT 1935.290 20.640 1935.610 20.700 ;
        RECT 1897.110 20.500 1935.610 20.640 ;
        RECT 1897.110 20.440 1897.430 20.500 ;
        RECT 1935.290 20.440 1935.610 20.500 ;
      LAYER via ;
        RECT 1891.620 287.680 1891.880 287.940 ;
        RECT 1897.140 287.680 1897.400 287.940 ;
        RECT 1897.140 20.440 1897.400 20.700 ;
        RECT 1935.320 20.440 1935.580 20.700 ;
      LAYER met2 ;
        RECT 1891.620 300.000 1891.900 304.000 ;
        RECT 1891.680 287.970 1891.820 300.000 ;
        RECT 1891.620 287.650 1891.880 287.970 ;
        RECT 1897.140 287.650 1897.400 287.970 ;
        RECT 1897.200 20.730 1897.340 287.650 ;
        RECT 1897.140 20.410 1897.400 20.730 ;
        RECT 1935.320 20.410 1935.580 20.730 ;
        RECT 1935.380 2.400 1935.520 20.410 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1906.310 288.220 1906.630 288.280 ;
        RECT 1910.450 288.220 1910.770 288.280 ;
        RECT 1906.310 288.080 1910.770 288.220 ;
        RECT 1906.310 288.020 1906.630 288.080 ;
        RECT 1910.450 288.020 1910.770 288.080 ;
        RECT 1910.450 17.920 1910.770 17.980 ;
        RECT 1953.230 17.920 1953.550 17.980 ;
        RECT 1910.450 17.780 1953.550 17.920 ;
        RECT 1910.450 17.720 1910.770 17.780 ;
        RECT 1953.230 17.720 1953.550 17.780 ;
      LAYER via ;
        RECT 1906.340 288.020 1906.600 288.280 ;
        RECT 1910.480 288.020 1910.740 288.280 ;
        RECT 1910.480 17.720 1910.740 17.980 ;
        RECT 1953.260 17.720 1953.520 17.980 ;
      LAYER met2 ;
        RECT 1906.340 300.000 1906.620 304.000 ;
        RECT 1906.400 288.310 1906.540 300.000 ;
        RECT 1906.340 287.990 1906.600 288.310 ;
        RECT 1910.480 287.990 1910.740 288.310 ;
        RECT 1910.540 18.010 1910.680 287.990 ;
        RECT 1910.480 17.690 1910.740 18.010 ;
        RECT 1953.260 17.690 1953.520 18.010 ;
        RECT 1953.320 2.400 1953.460 17.690 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1921.030 286.860 1921.350 286.920 ;
        RECT 1924.710 286.860 1925.030 286.920 ;
        RECT 1921.030 286.720 1925.030 286.860 ;
        RECT 1921.030 286.660 1921.350 286.720 ;
        RECT 1924.710 286.660 1925.030 286.720 ;
        RECT 1924.710 20.300 1925.030 20.360 ;
        RECT 1971.170 20.300 1971.490 20.360 ;
        RECT 1924.710 20.160 1971.490 20.300 ;
        RECT 1924.710 20.100 1925.030 20.160 ;
        RECT 1971.170 20.100 1971.490 20.160 ;
      LAYER via ;
        RECT 1921.060 286.660 1921.320 286.920 ;
        RECT 1924.740 286.660 1925.000 286.920 ;
        RECT 1924.740 20.100 1925.000 20.360 ;
        RECT 1971.200 20.100 1971.460 20.360 ;
      LAYER met2 ;
        RECT 1921.060 300.000 1921.340 304.000 ;
        RECT 1921.120 286.950 1921.260 300.000 ;
        RECT 1921.060 286.630 1921.320 286.950 ;
        RECT 1924.740 286.630 1925.000 286.950 ;
        RECT 1924.800 20.390 1924.940 286.630 ;
        RECT 1924.740 20.070 1925.000 20.390 ;
        RECT 1971.200 20.070 1971.460 20.390 ;
        RECT 1971.260 2.400 1971.400 20.070 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1938.510 18.260 1938.830 18.320 ;
        RECT 1989.110 18.260 1989.430 18.320 ;
        RECT 1938.510 18.120 1989.430 18.260 ;
        RECT 1938.510 18.060 1938.830 18.120 ;
        RECT 1989.110 18.060 1989.430 18.120 ;
      LAYER via ;
        RECT 1938.540 18.060 1938.800 18.320 ;
        RECT 1989.140 18.060 1989.400 18.320 ;
      LAYER met2 ;
        RECT 1935.780 300.290 1936.060 304.000 ;
        RECT 1935.780 300.150 1938.740 300.290 ;
        RECT 1935.780 300.000 1936.060 300.150 ;
        RECT 1938.600 18.350 1938.740 300.150 ;
        RECT 1938.540 18.030 1938.800 18.350 ;
        RECT 1989.140 18.030 1989.400 18.350 ;
        RECT 1989.200 2.400 1989.340 18.030 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1952.310 18.940 1952.630 19.000 ;
        RECT 2006.590 18.940 2006.910 19.000 ;
        RECT 1952.310 18.800 2006.910 18.940 ;
        RECT 1952.310 18.740 1952.630 18.800 ;
        RECT 2006.590 18.740 2006.910 18.800 ;
      LAYER via ;
        RECT 1952.340 18.740 1952.600 19.000 ;
        RECT 2006.620 18.740 2006.880 19.000 ;
      LAYER met2 ;
        RECT 1950.500 300.290 1950.780 304.000 ;
        RECT 1950.500 300.150 1952.540 300.290 ;
        RECT 1950.500 300.000 1950.780 300.150 ;
        RECT 1952.400 19.030 1952.540 300.150 ;
        RECT 1952.340 18.710 1952.600 19.030 ;
        RECT 2006.620 18.710 2006.880 19.030 ;
        RECT 2006.680 2.400 2006.820 18.710 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1965.650 19.620 1965.970 19.680 ;
        RECT 2024.530 19.620 2024.850 19.680 ;
        RECT 1965.650 19.480 2024.850 19.620 ;
        RECT 1965.650 19.420 1965.970 19.480 ;
        RECT 2024.530 19.420 2024.850 19.480 ;
      LAYER via ;
        RECT 1965.680 19.420 1965.940 19.680 ;
        RECT 2024.560 19.420 2024.820 19.680 ;
      LAYER met2 ;
        RECT 1964.760 300.290 1965.040 304.000 ;
        RECT 1964.760 300.150 1965.880 300.290 ;
        RECT 1964.760 300.000 1965.040 300.150 ;
        RECT 1965.740 19.710 1965.880 300.150 ;
        RECT 1965.680 19.390 1965.940 19.710 ;
        RECT 2024.560 19.390 2024.820 19.710 ;
        RECT 2024.620 2.400 2024.760 19.390 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1979.910 17.920 1980.230 17.980 ;
        RECT 2042.470 17.920 2042.790 17.980 ;
        RECT 1979.910 17.780 2042.790 17.920 ;
        RECT 1979.910 17.720 1980.230 17.780 ;
        RECT 2042.470 17.720 2042.790 17.780 ;
      LAYER via ;
        RECT 1979.940 17.720 1980.200 17.980 ;
        RECT 2042.500 17.720 2042.760 17.980 ;
      LAYER met2 ;
        RECT 1979.480 300.290 1979.760 304.000 ;
        RECT 1979.480 300.150 1980.140 300.290 ;
        RECT 1979.480 300.000 1979.760 300.150 ;
        RECT 1980.000 18.010 1980.140 300.150 ;
        RECT 1979.940 17.690 1980.200 18.010 ;
        RECT 2042.500 17.690 2042.760 18.010 ;
        RECT 2042.560 2.400 2042.700 17.690 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 757.690 18.260 758.010 18.320 ;
        RECT 917.770 18.260 918.090 18.320 ;
        RECT 757.690 18.120 918.090 18.260 ;
        RECT 757.690 18.060 758.010 18.120 ;
        RECT 917.770 18.060 918.090 18.120 ;
      LAYER via ;
        RECT 757.720 18.060 757.980 18.320 ;
        RECT 917.800 18.060 918.060 18.320 ;
      LAYER met2 ;
        RECT 921.940 300.290 922.220 304.000 ;
        RECT 917.860 300.150 922.220 300.290 ;
        RECT 917.860 18.350 918.000 300.150 ;
        RECT 921.940 300.000 922.220 300.150 ;
        RECT 757.720 18.030 757.980 18.350 ;
        RECT 917.800 18.030 918.060 18.350 ;
        RECT 757.780 2.400 757.920 18.030 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1994.170 288.220 1994.490 288.280 ;
        RECT 2000.150 288.220 2000.470 288.280 ;
        RECT 1994.170 288.080 2000.470 288.220 ;
        RECT 1994.170 288.020 1994.490 288.080 ;
        RECT 2000.150 288.020 2000.470 288.080 ;
        RECT 2000.150 19.960 2000.470 20.020 ;
        RECT 2060.410 19.960 2060.730 20.020 ;
        RECT 2000.150 19.820 2060.730 19.960 ;
        RECT 2000.150 19.760 2000.470 19.820 ;
        RECT 2060.410 19.760 2060.730 19.820 ;
      LAYER via ;
        RECT 1994.200 288.020 1994.460 288.280 ;
        RECT 2000.180 288.020 2000.440 288.280 ;
        RECT 2000.180 19.760 2000.440 20.020 ;
        RECT 2060.440 19.760 2060.700 20.020 ;
      LAYER met2 ;
        RECT 1994.200 300.000 1994.480 304.000 ;
        RECT 1994.260 288.310 1994.400 300.000 ;
        RECT 1994.200 287.990 1994.460 288.310 ;
        RECT 2000.180 287.990 2000.440 288.310 ;
        RECT 2000.240 20.050 2000.380 287.990 ;
        RECT 2000.180 19.730 2000.440 20.050 ;
        RECT 2060.440 19.730 2060.700 20.050 ;
        RECT 2060.500 2.400 2060.640 19.730 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2008.890 288.220 2009.210 288.280 ;
        RECT 2013.950 288.220 2014.270 288.280 ;
        RECT 2008.890 288.080 2014.270 288.220 ;
        RECT 2008.890 288.020 2009.210 288.080 ;
        RECT 2013.950 288.020 2014.270 288.080 ;
        RECT 2013.950 18.260 2014.270 18.320 ;
        RECT 2078.350 18.260 2078.670 18.320 ;
        RECT 2013.950 18.120 2078.670 18.260 ;
        RECT 2013.950 18.060 2014.270 18.120 ;
        RECT 2078.350 18.060 2078.670 18.120 ;
      LAYER via ;
        RECT 2008.920 288.020 2009.180 288.280 ;
        RECT 2013.980 288.020 2014.240 288.280 ;
        RECT 2013.980 18.060 2014.240 18.320 ;
        RECT 2078.380 18.060 2078.640 18.320 ;
      LAYER met2 ;
        RECT 2008.920 300.000 2009.200 304.000 ;
        RECT 2008.980 288.310 2009.120 300.000 ;
        RECT 2008.920 287.990 2009.180 288.310 ;
        RECT 2013.980 287.990 2014.240 288.310 ;
        RECT 2014.040 18.350 2014.180 287.990 ;
        RECT 2013.980 18.030 2014.240 18.350 ;
        RECT 2078.380 18.030 2078.640 18.350 ;
        RECT 2078.440 2.400 2078.580 18.030 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2023.610 288.220 2023.930 288.280 ;
        RECT 2028.210 288.220 2028.530 288.280 ;
        RECT 2023.610 288.080 2028.530 288.220 ;
        RECT 2023.610 288.020 2023.930 288.080 ;
        RECT 2028.210 288.020 2028.530 288.080 ;
        RECT 2028.210 16.900 2028.530 16.960 ;
        RECT 2095.830 16.900 2096.150 16.960 ;
        RECT 2028.210 16.760 2096.150 16.900 ;
        RECT 2028.210 16.700 2028.530 16.760 ;
        RECT 2095.830 16.700 2096.150 16.760 ;
      LAYER via ;
        RECT 2023.640 288.020 2023.900 288.280 ;
        RECT 2028.240 288.020 2028.500 288.280 ;
        RECT 2028.240 16.700 2028.500 16.960 ;
        RECT 2095.860 16.700 2096.120 16.960 ;
      LAYER met2 ;
        RECT 2023.640 300.000 2023.920 304.000 ;
        RECT 2023.700 288.310 2023.840 300.000 ;
        RECT 2023.640 287.990 2023.900 288.310 ;
        RECT 2028.240 287.990 2028.500 288.310 ;
        RECT 2028.300 16.990 2028.440 287.990 ;
        RECT 2028.240 16.670 2028.500 16.990 ;
        RECT 2095.860 16.670 2096.120 16.990 ;
        RECT 2095.920 2.400 2096.060 16.670 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2042.010 17.240 2042.330 17.300 ;
        RECT 2113.770 17.240 2114.090 17.300 ;
        RECT 2042.010 17.100 2114.090 17.240 ;
        RECT 2042.010 17.040 2042.330 17.100 ;
        RECT 2113.770 17.040 2114.090 17.100 ;
      LAYER via ;
        RECT 2042.040 17.040 2042.300 17.300 ;
        RECT 2113.800 17.040 2114.060 17.300 ;
      LAYER met2 ;
        RECT 2038.360 300.290 2038.640 304.000 ;
        RECT 2038.360 300.150 2042.240 300.290 ;
        RECT 2038.360 300.000 2038.640 300.150 ;
        RECT 2042.100 17.330 2042.240 300.150 ;
        RECT 2042.040 17.010 2042.300 17.330 ;
        RECT 2113.800 17.010 2114.060 17.330 ;
        RECT 2113.860 2.400 2114.000 17.010 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2055.810 15.880 2056.130 15.940 ;
        RECT 2131.710 15.880 2132.030 15.940 ;
        RECT 2055.810 15.740 2132.030 15.880 ;
        RECT 2055.810 15.680 2056.130 15.740 ;
        RECT 2131.710 15.680 2132.030 15.740 ;
      LAYER via ;
        RECT 2055.840 15.680 2056.100 15.940 ;
        RECT 2131.740 15.680 2132.000 15.940 ;
      LAYER met2 ;
        RECT 2053.080 300.290 2053.360 304.000 ;
        RECT 2053.080 300.150 2056.040 300.290 ;
        RECT 2053.080 300.000 2053.360 300.150 ;
        RECT 2055.900 15.970 2056.040 300.150 ;
        RECT 2055.840 15.650 2056.100 15.970 ;
        RECT 2131.740 15.650 2132.000 15.970 ;
        RECT 2131.800 2.400 2131.940 15.650 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2069.610 18.600 2069.930 18.660 ;
        RECT 2149.650 18.600 2149.970 18.660 ;
        RECT 2069.610 18.460 2149.970 18.600 ;
        RECT 2069.610 18.400 2069.930 18.460 ;
        RECT 2149.650 18.400 2149.970 18.460 ;
      LAYER via ;
        RECT 2069.640 18.400 2069.900 18.660 ;
        RECT 2149.680 18.400 2149.940 18.660 ;
      LAYER met2 ;
        RECT 2067.800 300.290 2068.080 304.000 ;
        RECT 2067.800 300.150 2069.840 300.290 ;
        RECT 2067.800 300.000 2068.080 300.150 ;
        RECT 2069.700 18.690 2069.840 300.150 ;
        RECT 2069.640 18.370 2069.900 18.690 ;
        RECT 2149.680 18.370 2149.940 18.690 ;
        RECT 2149.740 2.400 2149.880 18.370 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2082.950 18.260 2083.270 18.320 ;
        RECT 2167.590 18.260 2167.910 18.320 ;
        RECT 2082.950 18.120 2167.910 18.260 ;
        RECT 2082.950 18.060 2083.270 18.120 ;
        RECT 2167.590 18.060 2167.910 18.120 ;
      LAYER via ;
        RECT 2082.980 18.060 2083.240 18.320 ;
        RECT 2167.620 18.060 2167.880 18.320 ;
      LAYER met2 ;
        RECT 2082.520 300.290 2082.800 304.000 ;
        RECT 2082.520 300.150 2083.180 300.290 ;
        RECT 2082.520 300.000 2082.800 300.150 ;
        RECT 2083.040 18.350 2083.180 300.150 ;
        RECT 2082.980 18.030 2083.240 18.350 ;
        RECT 2167.620 18.030 2167.880 18.350 ;
        RECT 2167.680 2.400 2167.820 18.030 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2096.750 17.580 2097.070 17.640 ;
        RECT 2185.070 17.580 2185.390 17.640 ;
        RECT 2096.750 17.440 2185.390 17.580 ;
        RECT 2096.750 17.380 2097.070 17.440 ;
        RECT 2185.070 17.380 2185.390 17.440 ;
      LAYER via ;
        RECT 2096.780 17.380 2097.040 17.640 ;
        RECT 2185.100 17.380 2185.360 17.640 ;
      LAYER met2 ;
        RECT 2097.240 300.290 2097.520 304.000 ;
        RECT 2096.840 300.150 2097.520 300.290 ;
        RECT 2096.840 17.670 2096.980 300.150 ;
        RECT 2097.240 300.000 2097.520 300.150 ;
        RECT 2096.780 17.350 2097.040 17.670 ;
        RECT 2185.100 17.350 2185.360 17.670 ;
        RECT 2185.160 2.400 2185.300 17.350 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2111.930 288.220 2112.250 288.280 ;
        RECT 2117.450 288.220 2117.770 288.280 ;
        RECT 2111.930 288.080 2117.770 288.220 ;
        RECT 2111.930 288.020 2112.250 288.080 ;
        RECT 2117.450 288.020 2117.770 288.080 ;
        RECT 2117.450 19.620 2117.770 19.680 ;
        RECT 2203.010 19.620 2203.330 19.680 ;
        RECT 2117.450 19.480 2203.330 19.620 ;
        RECT 2117.450 19.420 2117.770 19.480 ;
        RECT 2203.010 19.420 2203.330 19.480 ;
      LAYER via ;
        RECT 2111.960 288.020 2112.220 288.280 ;
        RECT 2117.480 288.020 2117.740 288.280 ;
        RECT 2117.480 19.420 2117.740 19.680 ;
        RECT 2203.040 19.420 2203.300 19.680 ;
      LAYER met2 ;
        RECT 2111.960 300.000 2112.240 304.000 ;
        RECT 2112.020 288.310 2112.160 300.000 ;
        RECT 2111.960 287.990 2112.220 288.310 ;
        RECT 2117.480 287.990 2117.740 288.310 ;
        RECT 2117.540 19.710 2117.680 287.990 ;
        RECT 2117.480 19.390 2117.740 19.710 ;
        RECT 2203.040 19.390 2203.300 19.710 ;
        RECT 2203.100 2.400 2203.240 19.390 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2126.650 288.220 2126.970 288.280 ;
        RECT 2131.250 288.220 2131.570 288.280 ;
        RECT 2126.650 288.080 2131.570 288.220 ;
        RECT 2126.650 288.020 2126.970 288.080 ;
        RECT 2131.250 288.020 2131.570 288.080 ;
        RECT 2131.250 15.540 2131.570 15.600 ;
        RECT 2220.950 15.540 2221.270 15.600 ;
        RECT 2131.250 15.400 2221.270 15.540 ;
        RECT 2131.250 15.340 2131.570 15.400 ;
        RECT 2220.950 15.340 2221.270 15.400 ;
      LAYER via ;
        RECT 2126.680 288.020 2126.940 288.280 ;
        RECT 2131.280 288.020 2131.540 288.280 ;
        RECT 2131.280 15.340 2131.540 15.600 ;
        RECT 2220.980 15.340 2221.240 15.600 ;
      LAYER met2 ;
        RECT 2126.680 300.000 2126.960 304.000 ;
        RECT 2126.740 288.310 2126.880 300.000 ;
        RECT 2126.680 287.990 2126.940 288.310 ;
        RECT 2131.280 287.990 2131.540 288.310 ;
        RECT 2131.340 15.630 2131.480 287.990 ;
        RECT 2131.280 15.310 2131.540 15.630 ;
        RECT 2220.980 15.310 2221.240 15.630 ;
        RECT 2221.040 2.400 2221.180 15.310 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 775.630 26.080 775.950 26.140 ;
        RECT 932.030 26.080 932.350 26.140 ;
        RECT 775.630 25.940 932.350 26.080 ;
        RECT 775.630 25.880 775.950 25.940 ;
        RECT 932.030 25.880 932.350 25.940 ;
      LAYER via ;
        RECT 775.660 25.880 775.920 26.140 ;
        RECT 932.060 25.880 932.320 26.140 ;
      LAYER met2 ;
        RECT 936.660 300.290 936.940 304.000 ;
        RECT 932.120 300.150 936.940 300.290 ;
        RECT 932.120 26.170 932.260 300.150 ;
        RECT 936.660 300.000 936.940 300.150 ;
        RECT 775.660 25.850 775.920 26.170 ;
        RECT 932.060 25.850 932.320 26.170 ;
        RECT 775.720 2.400 775.860 25.850 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2141.370 288.220 2141.690 288.280 ;
        RECT 2145.510 288.220 2145.830 288.280 ;
        RECT 2141.370 288.080 2145.830 288.220 ;
        RECT 2141.370 288.020 2141.690 288.080 ;
        RECT 2145.510 288.020 2145.830 288.080 ;
        RECT 2145.510 19.960 2145.830 20.020 ;
        RECT 2238.890 19.960 2239.210 20.020 ;
        RECT 2145.510 19.820 2239.210 19.960 ;
        RECT 2145.510 19.760 2145.830 19.820 ;
        RECT 2238.890 19.760 2239.210 19.820 ;
      LAYER via ;
        RECT 2141.400 288.020 2141.660 288.280 ;
        RECT 2145.540 288.020 2145.800 288.280 ;
        RECT 2145.540 19.760 2145.800 20.020 ;
        RECT 2238.920 19.760 2239.180 20.020 ;
      LAYER met2 ;
        RECT 2141.400 300.000 2141.680 304.000 ;
        RECT 2141.460 288.310 2141.600 300.000 ;
        RECT 2141.400 287.990 2141.660 288.310 ;
        RECT 2145.540 287.990 2145.800 288.310 ;
        RECT 2145.600 20.050 2145.740 287.990 ;
        RECT 2145.540 19.730 2145.800 20.050 ;
        RECT 2238.920 19.730 2239.180 20.050 ;
        RECT 2238.980 2.400 2239.120 19.730 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2159.310 20.640 2159.630 20.700 ;
        RECT 2256.370 20.640 2256.690 20.700 ;
        RECT 2159.310 20.500 2256.690 20.640 ;
        RECT 2159.310 20.440 2159.630 20.500 ;
        RECT 2256.370 20.440 2256.690 20.500 ;
      LAYER via ;
        RECT 2159.340 20.440 2159.600 20.700 ;
        RECT 2256.400 20.440 2256.660 20.700 ;
      LAYER met2 ;
        RECT 2156.120 300.290 2156.400 304.000 ;
        RECT 2156.120 300.150 2159.540 300.290 ;
        RECT 2156.120 300.000 2156.400 300.150 ;
        RECT 2159.400 20.730 2159.540 300.150 ;
        RECT 2159.340 20.410 2159.600 20.730 ;
        RECT 2256.400 20.410 2256.660 20.730 ;
        RECT 2256.460 2.400 2256.600 20.410 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2173.110 19.280 2173.430 19.340 ;
        RECT 2274.310 19.280 2274.630 19.340 ;
        RECT 2173.110 19.140 2274.630 19.280 ;
        RECT 2173.110 19.080 2173.430 19.140 ;
        RECT 2274.310 19.080 2274.630 19.140 ;
      LAYER via ;
        RECT 2173.140 19.080 2173.400 19.340 ;
        RECT 2274.340 19.080 2274.600 19.340 ;
      LAYER met2 ;
        RECT 2170.840 300.290 2171.120 304.000 ;
        RECT 2170.840 300.150 2173.340 300.290 ;
        RECT 2170.840 300.000 2171.120 300.150 ;
        RECT 2173.200 19.370 2173.340 300.150 ;
        RECT 2173.140 19.050 2173.400 19.370 ;
        RECT 2274.340 19.050 2274.600 19.370 ;
        RECT 2274.400 2.400 2274.540 19.050 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2185.530 286.180 2185.850 286.240 ;
        RECT 2291.330 286.180 2291.650 286.240 ;
        RECT 2185.530 286.040 2291.650 286.180 ;
        RECT 2185.530 285.980 2185.850 286.040 ;
        RECT 2291.330 285.980 2291.650 286.040 ;
      LAYER via ;
        RECT 2185.560 285.980 2185.820 286.240 ;
        RECT 2291.360 285.980 2291.620 286.240 ;
      LAYER met2 ;
        RECT 2185.560 300.000 2185.840 304.000 ;
        RECT 2185.620 286.270 2185.760 300.000 ;
        RECT 2185.560 285.950 2185.820 286.270 ;
        RECT 2291.360 285.950 2291.620 286.270 ;
        RECT 2291.420 3.130 2291.560 285.950 ;
        RECT 2291.420 2.990 2292.480 3.130 ;
        RECT 2292.340 2.400 2292.480 2.990 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2280.365 17.425 2280.535 19.635 ;
      LAYER mcon ;
        RECT 2280.365 19.465 2280.535 19.635 ;
      LAYER met1 ;
        RECT 2280.305 19.620 2280.595 19.665 ;
        RECT 2310.190 19.620 2310.510 19.680 ;
        RECT 2280.305 19.480 2310.510 19.620 ;
        RECT 2280.305 19.435 2280.595 19.480 ;
        RECT 2310.190 19.420 2310.510 19.480 ;
        RECT 2200.250 17.580 2200.570 17.640 ;
        RECT 2280.305 17.580 2280.595 17.625 ;
        RECT 2200.250 17.440 2280.595 17.580 ;
        RECT 2200.250 17.380 2200.570 17.440 ;
        RECT 2280.305 17.395 2280.595 17.440 ;
      LAYER via ;
        RECT 2310.220 19.420 2310.480 19.680 ;
        RECT 2200.280 17.380 2200.540 17.640 ;
      LAYER met2 ;
        RECT 2200.280 300.000 2200.560 304.000 ;
        RECT 2200.340 17.670 2200.480 300.000 ;
        RECT 2310.220 19.390 2310.480 19.710 ;
        RECT 2200.280 17.350 2200.540 17.670 ;
        RECT 2310.280 2.400 2310.420 19.390 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2214.050 17.240 2214.370 17.300 ;
        RECT 2328.130 17.240 2328.450 17.300 ;
        RECT 2214.050 17.100 2328.450 17.240 ;
        RECT 2214.050 17.040 2214.370 17.100 ;
        RECT 2328.130 17.040 2328.450 17.100 ;
      LAYER via ;
        RECT 2214.080 17.040 2214.340 17.300 ;
        RECT 2328.160 17.040 2328.420 17.300 ;
      LAYER met2 ;
        RECT 2214.540 300.290 2214.820 304.000 ;
        RECT 2214.140 300.150 2214.820 300.290 ;
        RECT 2214.140 17.330 2214.280 300.150 ;
        RECT 2214.540 300.000 2214.820 300.150 ;
        RECT 2214.080 17.010 2214.340 17.330 ;
        RECT 2328.160 17.010 2328.420 17.330 ;
        RECT 2328.220 2.400 2328.360 17.010 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2229.230 285.500 2229.550 285.560 ;
        RECT 2234.750 285.500 2235.070 285.560 ;
        RECT 2229.230 285.360 2235.070 285.500 ;
        RECT 2229.230 285.300 2229.550 285.360 ;
        RECT 2234.750 285.300 2235.070 285.360 ;
        RECT 2234.750 15.540 2235.070 15.600 ;
        RECT 2241.650 15.540 2241.970 15.600 ;
        RECT 2234.750 15.400 2241.970 15.540 ;
        RECT 2234.750 15.340 2235.070 15.400 ;
        RECT 2241.650 15.340 2241.970 15.400 ;
        RECT 2255.910 15.200 2256.230 15.260 ;
        RECT 2345.610 15.200 2345.930 15.260 ;
        RECT 2255.910 15.060 2345.930 15.200 ;
        RECT 2255.910 15.000 2256.230 15.060 ;
        RECT 2345.610 15.000 2345.930 15.060 ;
      LAYER via ;
        RECT 2229.260 285.300 2229.520 285.560 ;
        RECT 2234.780 285.300 2235.040 285.560 ;
        RECT 2234.780 15.340 2235.040 15.600 ;
        RECT 2241.680 15.340 2241.940 15.600 ;
        RECT 2255.940 15.000 2256.200 15.260 ;
        RECT 2345.640 15.000 2345.900 15.260 ;
      LAYER met2 ;
        RECT 2229.260 300.000 2229.540 304.000 ;
        RECT 2229.320 285.590 2229.460 300.000 ;
        RECT 2229.260 285.270 2229.520 285.590 ;
        RECT 2234.780 285.270 2235.040 285.590 ;
        RECT 2234.840 15.630 2234.980 285.270 ;
        RECT 2234.780 15.310 2235.040 15.630 ;
        RECT 2241.680 15.485 2241.940 15.630 ;
        RECT 2241.670 15.115 2241.950 15.485 ;
        RECT 2255.930 15.115 2256.210 15.485 ;
        RECT 2255.940 14.970 2256.200 15.115 ;
        RECT 2345.640 14.970 2345.900 15.290 ;
        RECT 2345.700 2.400 2345.840 14.970 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
      LAYER via2 ;
        RECT 2241.670 15.160 2241.950 15.440 ;
        RECT 2255.930 15.160 2256.210 15.440 ;
      LAYER met3 ;
        RECT 2241.645 15.450 2241.975 15.465 ;
        RECT 2255.905 15.450 2256.235 15.465 ;
        RECT 2241.645 15.150 2256.235 15.450 ;
        RECT 2241.645 15.135 2241.975 15.150 ;
        RECT 2255.905 15.135 2256.235 15.150 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2243.950 288.220 2244.270 288.280 ;
        RECT 2248.550 288.220 2248.870 288.280 ;
        RECT 2243.950 288.080 2248.870 288.220 ;
        RECT 2243.950 288.020 2244.270 288.080 ;
        RECT 2248.550 288.020 2248.870 288.080 ;
        RECT 2248.550 20.300 2248.870 20.360 ;
        RECT 2363.550 20.300 2363.870 20.360 ;
        RECT 2248.550 20.160 2363.870 20.300 ;
        RECT 2248.550 20.100 2248.870 20.160 ;
        RECT 2363.550 20.100 2363.870 20.160 ;
      LAYER via ;
        RECT 2243.980 288.020 2244.240 288.280 ;
        RECT 2248.580 288.020 2248.840 288.280 ;
        RECT 2248.580 20.100 2248.840 20.360 ;
        RECT 2363.580 20.100 2363.840 20.360 ;
      LAYER met2 ;
        RECT 2243.980 300.000 2244.260 304.000 ;
        RECT 2244.040 288.310 2244.180 300.000 ;
        RECT 2243.980 287.990 2244.240 288.310 ;
        RECT 2248.580 287.990 2248.840 288.310 ;
        RECT 2248.640 20.390 2248.780 287.990 ;
        RECT 2248.580 20.070 2248.840 20.390 ;
        RECT 2363.580 20.070 2363.840 20.390 ;
        RECT 2363.640 2.400 2363.780 20.070 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2258.670 288.220 2258.990 288.280 ;
        RECT 2262.810 288.220 2263.130 288.280 ;
        RECT 2258.670 288.080 2263.130 288.220 ;
        RECT 2258.670 288.020 2258.990 288.080 ;
        RECT 2262.810 288.020 2263.130 288.080 ;
        RECT 2262.810 20.640 2263.130 20.700 ;
        RECT 2381.490 20.640 2381.810 20.700 ;
        RECT 2262.810 20.500 2381.810 20.640 ;
        RECT 2262.810 20.440 2263.130 20.500 ;
        RECT 2381.490 20.440 2381.810 20.500 ;
      LAYER via ;
        RECT 2258.700 288.020 2258.960 288.280 ;
        RECT 2262.840 288.020 2263.100 288.280 ;
        RECT 2262.840 20.440 2263.100 20.700 ;
        RECT 2381.520 20.440 2381.780 20.700 ;
      LAYER met2 ;
        RECT 2258.700 300.000 2258.980 304.000 ;
        RECT 2258.760 288.310 2258.900 300.000 ;
        RECT 2258.700 287.990 2258.960 288.310 ;
        RECT 2262.840 287.990 2263.100 288.310 ;
        RECT 2262.900 20.730 2263.040 287.990 ;
        RECT 2262.840 20.410 2263.100 20.730 ;
        RECT 2381.520 20.410 2381.780 20.730 ;
        RECT 2381.580 2.400 2381.720 20.410 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2279.445 14.535 2279.615 16.575 ;
        RECT 2279.445 14.365 2280.995 14.535 ;
      LAYER mcon ;
        RECT 2279.445 16.405 2279.615 16.575 ;
        RECT 2280.825 14.365 2280.995 14.535 ;
      LAYER met1 ;
        RECT 2276.610 16.560 2276.930 16.620 ;
        RECT 2279.385 16.560 2279.675 16.605 ;
        RECT 2276.610 16.420 2279.675 16.560 ;
        RECT 2276.610 16.360 2276.930 16.420 ;
        RECT 2279.385 16.375 2279.675 16.420 ;
        RECT 2280.765 14.520 2281.055 14.565 ;
        RECT 2399.430 14.520 2399.750 14.580 ;
        RECT 2280.765 14.380 2399.750 14.520 ;
        RECT 2280.765 14.335 2281.055 14.380 ;
        RECT 2399.430 14.320 2399.750 14.380 ;
      LAYER via ;
        RECT 2276.640 16.360 2276.900 16.620 ;
        RECT 2399.460 14.320 2399.720 14.580 ;
      LAYER met2 ;
        RECT 2273.420 300.290 2273.700 304.000 ;
        RECT 2273.420 300.150 2276.840 300.290 ;
        RECT 2273.420 300.000 2273.700 300.150 ;
        RECT 2276.700 16.650 2276.840 300.150 ;
        RECT 2276.640 16.330 2276.900 16.650 ;
        RECT 2399.460 14.290 2399.720 14.610 ;
        RECT 2399.520 2.400 2399.660 14.290 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 799.550 285.160 799.870 285.220 ;
        RECT 951.350 285.160 951.670 285.220 ;
        RECT 799.550 285.020 951.670 285.160 ;
        RECT 799.550 284.960 799.870 285.020 ;
        RECT 951.350 284.960 951.670 285.020 ;
        RECT 793.570 17.920 793.890 17.980 ;
        RECT 799.550 17.920 799.870 17.980 ;
        RECT 793.570 17.780 799.870 17.920 ;
        RECT 793.570 17.720 793.890 17.780 ;
        RECT 799.550 17.720 799.870 17.780 ;
      LAYER via ;
        RECT 799.580 284.960 799.840 285.220 ;
        RECT 951.380 284.960 951.640 285.220 ;
        RECT 793.600 17.720 793.860 17.980 ;
        RECT 799.580 17.720 799.840 17.980 ;
      LAYER met2 ;
        RECT 951.380 300.000 951.660 304.000 ;
        RECT 951.440 285.250 951.580 300.000 ;
        RECT 799.580 284.930 799.840 285.250 ;
        RECT 951.380 284.930 951.640 285.250 ;
        RECT 799.640 18.010 799.780 284.930 ;
        RECT 793.600 17.690 793.860 18.010 ;
        RECT 799.580 17.690 799.840 18.010 ;
        RECT 793.660 2.400 793.800 17.690 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 639.010 24.380 639.330 24.440 ;
        RECT 821.170 24.380 821.490 24.440 ;
        RECT 639.010 24.240 821.490 24.380 ;
        RECT 639.010 24.180 639.330 24.240 ;
        RECT 821.170 24.180 821.490 24.240 ;
      LAYER via ;
        RECT 639.040 24.180 639.300 24.440 ;
        RECT 821.200 24.180 821.460 24.440 ;
      LAYER met2 ;
        RECT 823.960 300.290 824.240 304.000 ;
        RECT 821.260 300.150 824.240 300.290 ;
        RECT 821.260 24.470 821.400 300.150 ;
        RECT 823.960 300.000 824.240 300.150 ;
        RECT 639.040 24.150 639.300 24.470 ;
        RECT 821.200 24.150 821.460 24.470 ;
        RECT 639.100 2.400 639.240 24.150 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2293.170 288.220 2293.490 288.280 ;
        RECT 2297.310 288.220 2297.630 288.280 ;
        RECT 2293.170 288.080 2297.630 288.220 ;
        RECT 2293.170 288.020 2293.490 288.080 ;
        RECT 2297.310 288.020 2297.630 288.080 ;
        RECT 2297.310 18.600 2297.630 18.660 ;
        RECT 2422.890 18.600 2423.210 18.660 ;
        RECT 2297.310 18.460 2423.210 18.600 ;
        RECT 2297.310 18.400 2297.630 18.460 ;
        RECT 2422.890 18.400 2423.210 18.460 ;
      LAYER via ;
        RECT 2293.200 288.020 2293.460 288.280 ;
        RECT 2297.340 288.020 2297.600 288.280 ;
        RECT 2297.340 18.400 2297.600 18.660 ;
        RECT 2422.920 18.400 2423.180 18.660 ;
      LAYER met2 ;
        RECT 2293.200 300.000 2293.480 304.000 ;
        RECT 2293.260 288.310 2293.400 300.000 ;
        RECT 2293.200 287.990 2293.460 288.310 ;
        RECT 2297.340 287.990 2297.600 288.310 ;
        RECT 2297.400 18.690 2297.540 287.990 ;
        RECT 2297.340 18.370 2297.600 18.690 ;
        RECT 2422.920 18.370 2423.180 18.690 ;
        RECT 2422.980 2.400 2423.120 18.370 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2311.110 19.280 2311.430 19.340 ;
        RECT 2440.830 19.280 2441.150 19.340 ;
        RECT 2311.110 19.140 2441.150 19.280 ;
        RECT 2311.110 19.080 2311.430 19.140 ;
        RECT 2440.830 19.080 2441.150 19.140 ;
      LAYER via ;
        RECT 2311.140 19.080 2311.400 19.340 ;
        RECT 2440.860 19.080 2441.120 19.340 ;
      LAYER met2 ;
        RECT 2307.920 300.290 2308.200 304.000 ;
        RECT 2307.920 300.150 2311.340 300.290 ;
        RECT 2307.920 300.000 2308.200 300.150 ;
        RECT 2311.200 19.370 2311.340 300.150 ;
        RECT 2311.140 19.050 2311.400 19.370 ;
        RECT 2440.860 19.050 2441.120 19.370 ;
        RECT 2440.920 2.400 2441.060 19.050 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2324.910 19.620 2325.230 19.680 ;
        RECT 2458.770 19.620 2459.090 19.680 ;
        RECT 2324.910 19.480 2459.090 19.620 ;
        RECT 2324.910 19.420 2325.230 19.480 ;
        RECT 2458.770 19.420 2459.090 19.480 ;
      LAYER via ;
        RECT 2324.940 19.420 2325.200 19.680 ;
        RECT 2458.800 19.420 2459.060 19.680 ;
      LAYER met2 ;
        RECT 2322.640 300.290 2322.920 304.000 ;
        RECT 2322.640 300.150 2325.140 300.290 ;
        RECT 2322.640 300.000 2322.920 300.150 ;
        RECT 2325.000 19.710 2325.140 300.150 ;
        RECT 2324.940 19.390 2325.200 19.710 ;
        RECT 2458.800 19.390 2459.060 19.710 ;
        RECT 2458.860 2.400 2459.000 19.390 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2476.710 15.200 2477.030 15.260 ;
        RECT 2346.160 15.060 2477.030 15.200 ;
        RECT 2338.710 14.860 2339.030 14.920 ;
        RECT 2346.160 14.860 2346.300 15.060 ;
        RECT 2476.710 15.000 2477.030 15.060 ;
        RECT 2338.710 14.720 2346.300 14.860 ;
        RECT 2338.710 14.660 2339.030 14.720 ;
      LAYER via ;
        RECT 2338.740 14.660 2339.000 14.920 ;
        RECT 2476.740 15.000 2477.000 15.260 ;
      LAYER met2 ;
        RECT 2337.360 300.290 2337.640 304.000 ;
        RECT 2337.360 300.150 2338.940 300.290 ;
        RECT 2337.360 300.000 2337.640 300.150 ;
        RECT 2338.800 14.950 2338.940 300.150 ;
        RECT 2476.740 14.970 2477.000 15.290 ;
        RECT 2338.740 14.630 2339.000 14.950 ;
        RECT 2476.800 2.400 2476.940 14.970 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2352.510 17.920 2352.830 17.980 ;
        RECT 2494.650 17.920 2494.970 17.980 ;
        RECT 2352.510 17.780 2494.970 17.920 ;
        RECT 2352.510 17.720 2352.830 17.780 ;
        RECT 2494.650 17.720 2494.970 17.780 ;
      LAYER via ;
        RECT 2352.540 17.720 2352.800 17.980 ;
        RECT 2494.680 17.720 2494.940 17.980 ;
      LAYER met2 ;
        RECT 2352.080 300.290 2352.360 304.000 ;
        RECT 2352.080 300.150 2352.740 300.290 ;
        RECT 2352.080 300.000 2352.360 300.150 ;
        RECT 2352.600 18.010 2352.740 300.150 ;
        RECT 2352.540 17.690 2352.800 18.010 ;
        RECT 2494.680 17.690 2494.940 18.010 ;
        RECT 2494.740 2.400 2494.880 17.690 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2366.770 287.880 2367.090 287.940 ;
        RECT 2372.750 287.880 2373.070 287.940 ;
        RECT 2366.770 287.740 2373.070 287.880 ;
        RECT 2366.770 287.680 2367.090 287.740 ;
        RECT 2372.750 287.680 2373.070 287.740 ;
        RECT 2372.750 20.300 2373.070 20.360 ;
        RECT 2512.130 20.300 2512.450 20.360 ;
        RECT 2372.750 20.160 2512.450 20.300 ;
        RECT 2372.750 20.100 2373.070 20.160 ;
        RECT 2512.130 20.100 2512.450 20.160 ;
      LAYER via ;
        RECT 2366.800 287.680 2367.060 287.940 ;
        RECT 2372.780 287.680 2373.040 287.940 ;
        RECT 2372.780 20.100 2373.040 20.360 ;
        RECT 2512.160 20.100 2512.420 20.360 ;
      LAYER met2 ;
        RECT 2366.800 300.000 2367.080 304.000 ;
        RECT 2366.860 287.970 2367.000 300.000 ;
        RECT 2366.800 287.650 2367.060 287.970 ;
        RECT 2372.780 287.650 2373.040 287.970 ;
        RECT 2372.840 20.390 2372.980 287.650 ;
        RECT 2372.780 20.070 2373.040 20.390 ;
        RECT 2512.160 20.070 2512.420 20.390 ;
        RECT 2512.220 2.400 2512.360 20.070 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2381.030 284.820 2381.350 284.880 ;
        RECT 2387.010 284.820 2387.330 284.880 ;
        RECT 2381.030 284.680 2387.330 284.820 ;
        RECT 2381.030 284.620 2381.350 284.680 ;
        RECT 2387.010 284.620 2387.330 284.680 ;
        RECT 2387.010 16.220 2387.330 16.280 ;
        RECT 2530.070 16.220 2530.390 16.280 ;
        RECT 2387.010 16.080 2530.390 16.220 ;
        RECT 2387.010 16.020 2387.330 16.080 ;
        RECT 2530.070 16.020 2530.390 16.080 ;
      LAYER via ;
        RECT 2381.060 284.620 2381.320 284.880 ;
        RECT 2387.040 284.620 2387.300 284.880 ;
        RECT 2387.040 16.020 2387.300 16.280 ;
        RECT 2530.100 16.020 2530.360 16.280 ;
      LAYER met2 ;
        RECT 2381.060 300.000 2381.340 304.000 ;
        RECT 2381.120 284.910 2381.260 300.000 ;
        RECT 2381.060 284.590 2381.320 284.910 ;
        RECT 2387.040 284.590 2387.300 284.910 ;
        RECT 2387.100 16.310 2387.240 284.590 ;
        RECT 2387.040 15.990 2387.300 16.310 ;
        RECT 2530.100 15.990 2530.360 16.310 ;
        RECT 2530.160 2.400 2530.300 15.990 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2395.750 286.180 2396.070 286.240 ;
        RECT 2400.810 286.180 2401.130 286.240 ;
        RECT 2395.750 286.040 2401.130 286.180 ;
        RECT 2395.750 285.980 2396.070 286.040 ;
        RECT 2400.810 285.980 2401.130 286.040 ;
        RECT 2400.810 16.560 2401.130 16.620 ;
        RECT 2548.010 16.560 2548.330 16.620 ;
        RECT 2400.810 16.420 2548.330 16.560 ;
        RECT 2400.810 16.360 2401.130 16.420 ;
        RECT 2548.010 16.360 2548.330 16.420 ;
      LAYER via ;
        RECT 2395.780 285.980 2396.040 286.240 ;
        RECT 2400.840 285.980 2401.100 286.240 ;
        RECT 2400.840 16.360 2401.100 16.620 ;
        RECT 2548.040 16.360 2548.300 16.620 ;
      LAYER met2 ;
        RECT 2395.780 300.000 2396.060 304.000 ;
        RECT 2395.840 286.270 2395.980 300.000 ;
        RECT 2395.780 285.950 2396.040 286.270 ;
        RECT 2400.840 285.950 2401.100 286.270 ;
        RECT 2400.900 16.650 2401.040 285.950 ;
        RECT 2400.840 16.330 2401.100 16.650 ;
        RECT 2548.040 16.330 2548.300 16.650 ;
        RECT 2548.100 2.400 2548.240 16.330 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2410.470 288.900 2410.790 288.960 ;
        RECT 2414.610 288.900 2414.930 288.960 ;
        RECT 2410.470 288.760 2414.930 288.900 ;
        RECT 2410.470 288.700 2410.790 288.760 ;
        RECT 2414.610 288.700 2414.930 288.760 ;
        RECT 2414.610 16.900 2414.930 16.960 ;
        RECT 2565.950 16.900 2566.270 16.960 ;
        RECT 2414.610 16.760 2566.270 16.900 ;
        RECT 2414.610 16.700 2414.930 16.760 ;
        RECT 2565.950 16.700 2566.270 16.760 ;
      LAYER via ;
        RECT 2410.500 288.700 2410.760 288.960 ;
        RECT 2414.640 288.700 2414.900 288.960 ;
        RECT 2414.640 16.700 2414.900 16.960 ;
        RECT 2565.980 16.700 2566.240 16.960 ;
      LAYER met2 ;
        RECT 2410.500 300.000 2410.780 304.000 ;
        RECT 2410.560 288.990 2410.700 300.000 ;
        RECT 2410.500 288.670 2410.760 288.990 ;
        RECT 2414.640 288.670 2414.900 288.990 ;
        RECT 2414.700 16.990 2414.840 288.670 ;
        RECT 2414.640 16.670 2414.900 16.990 ;
        RECT 2565.980 16.670 2566.240 16.990 ;
        RECT 2566.040 2.400 2566.180 16.670 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2428.410 18.940 2428.730 19.000 ;
        RECT 2583.890 18.940 2584.210 19.000 ;
        RECT 2428.410 18.800 2584.210 18.940 ;
        RECT 2428.410 18.740 2428.730 18.800 ;
        RECT 2583.890 18.740 2584.210 18.800 ;
      LAYER via ;
        RECT 2428.440 18.740 2428.700 19.000 ;
        RECT 2583.920 18.740 2584.180 19.000 ;
      LAYER met2 ;
        RECT 2425.220 300.290 2425.500 304.000 ;
        RECT 2425.220 300.150 2428.640 300.290 ;
        RECT 2425.220 300.000 2425.500 300.150 ;
        RECT 2428.500 19.030 2428.640 300.150 ;
        RECT 2428.440 18.710 2428.700 19.030 ;
        RECT 2583.920 18.710 2584.180 19.030 ;
        RECT 2583.980 2.400 2584.120 18.710 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 847.005 284.325 847.175 286.535 ;
      LAYER mcon ;
        RECT 847.005 286.365 847.175 286.535 ;
      LAYER met1 ;
        RECT 846.945 286.520 847.235 286.565 ;
        RECT 970.670 286.520 970.990 286.580 ;
        RECT 846.945 286.380 970.990 286.520 ;
        RECT 846.945 286.335 847.235 286.380 ;
        RECT 970.670 286.320 970.990 286.380 ;
        RECT 820.710 284.480 821.030 284.540 ;
        RECT 846.945 284.480 847.235 284.525 ;
        RECT 820.710 284.340 847.235 284.480 ;
        RECT 820.710 284.280 821.030 284.340 ;
        RECT 846.945 284.295 847.235 284.340 ;
        RECT 817.490 17.580 817.810 17.640 ;
        RECT 820.710 17.580 821.030 17.640 ;
        RECT 817.490 17.440 821.030 17.580 ;
        RECT 817.490 17.380 817.810 17.440 ;
        RECT 820.710 17.380 821.030 17.440 ;
      LAYER via ;
        RECT 970.700 286.320 970.960 286.580 ;
        RECT 820.740 284.280 821.000 284.540 ;
        RECT 817.520 17.380 817.780 17.640 ;
        RECT 820.740 17.380 821.000 17.640 ;
      LAYER met2 ;
        RECT 970.700 300.000 970.980 304.000 ;
        RECT 970.760 286.610 970.900 300.000 ;
        RECT 970.700 286.290 970.960 286.610 ;
        RECT 820.740 284.250 821.000 284.570 ;
        RECT 820.800 17.670 820.940 284.250 ;
        RECT 817.520 17.350 817.780 17.670 ;
        RECT 820.740 17.350 821.000 17.670 ;
        RECT 817.580 2.400 817.720 17.350 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2442.210 18.600 2442.530 18.660 ;
        RECT 2601.370 18.600 2601.690 18.660 ;
        RECT 2442.210 18.460 2601.690 18.600 ;
        RECT 2442.210 18.400 2442.530 18.460 ;
        RECT 2601.370 18.400 2601.690 18.460 ;
      LAYER via ;
        RECT 2442.240 18.400 2442.500 18.660 ;
        RECT 2601.400 18.400 2601.660 18.660 ;
      LAYER met2 ;
        RECT 2439.940 300.290 2440.220 304.000 ;
        RECT 2439.940 300.150 2442.440 300.290 ;
        RECT 2439.940 300.000 2440.220 300.150 ;
        RECT 2442.300 18.690 2442.440 300.150 ;
        RECT 2442.240 18.370 2442.500 18.690 ;
        RECT 2601.400 18.370 2601.660 18.690 ;
        RECT 2601.460 2.400 2601.600 18.370 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2456.010 18.260 2456.330 18.320 ;
        RECT 2619.310 18.260 2619.630 18.320 ;
        RECT 2456.010 18.120 2619.630 18.260 ;
        RECT 2456.010 18.060 2456.330 18.120 ;
        RECT 2619.310 18.060 2619.630 18.120 ;
      LAYER via ;
        RECT 2456.040 18.060 2456.300 18.320 ;
        RECT 2619.340 18.060 2619.600 18.320 ;
      LAYER met2 ;
        RECT 2454.660 300.290 2454.940 304.000 ;
        RECT 2454.660 300.150 2456.240 300.290 ;
        RECT 2454.660 300.000 2454.940 300.150 ;
        RECT 2456.100 18.350 2456.240 300.150 ;
        RECT 2456.040 18.030 2456.300 18.350 ;
        RECT 2619.340 18.030 2619.600 18.350 ;
        RECT 2619.400 2.400 2619.540 18.030 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2469.810 17.580 2470.130 17.640 ;
        RECT 2637.250 17.580 2637.570 17.640 ;
        RECT 2469.810 17.440 2637.570 17.580 ;
        RECT 2469.810 17.380 2470.130 17.440 ;
        RECT 2637.250 17.380 2637.570 17.440 ;
      LAYER via ;
        RECT 2469.840 17.380 2470.100 17.640 ;
        RECT 2637.280 17.380 2637.540 17.640 ;
      LAYER met2 ;
        RECT 2469.380 300.290 2469.660 304.000 ;
        RECT 2469.380 300.150 2470.040 300.290 ;
        RECT 2469.380 300.000 2469.660 300.150 ;
        RECT 2469.900 17.670 2470.040 300.150 ;
        RECT 2469.840 17.350 2470.100 17.670 ;
        RECT 2637.280 17.350 2637.540 17.670 ;
        RECT 2637.340 2.400 2637.480 17.350 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2484.070 288.220 2484.390 288.280 ;
        RECT 2490.510 288.220 2490.830 288.280 ;
        RECT 2484.070 288.080 2490.830 288.220 ;
        RECT 2484.070 288.020 2484.390 288.080 ;
        RECT 2490.510 288.020 2490.830 288.080 ;
        RECT 2490.510 14.860 2490.830 14.920 ;
        RECT 2655.190 14.860 2655.510 14.920 ;
        RECT 2490.510 14.720 2655.510 14.860 ;
        RECT 2490.510 14.660 2490.830 14.720 ;
        RECT 2655.190 14.660 2655.510 14.720 ;
      LAYER via ;
        RECT 2484.100 288.020 2484.360 288.280 ;
        RECT 2490.540 288.020 2490.800 288.280 ;
        RECT 2490.540 14.660 2490.800 14.920 ;
        RECT 2655.220 14.660 2655.480 14.920 ;
      LAYER met2 ;
        RECT 2484.100 300.000 2484.380 304.000 ;
        RECT 2484.160 288.310 2484.300 300.000 ;
        RECT 2484.100 287.990 2484.360 288.310 ;
        RECT 2490.540 287.990 2490.800 288.310 ;
        RECT 2490.600 14.950 2490.740 287.990 ;
        RECT 2490.540 14.630 2490.800 14.950 ;
        RECT 2655.220 14.630 2655.480 14.950 ;
        RECT 2655.280 2.400 2655.420 14.630 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2498.790 288.220 2499.110 288.280 ;
        RECT 2504.310 288.220 2504.630 288.280 ;
        RECT 2498.790 288.080 2504.630 288.220 ;
        RECT 2498.790 288.020 2499.110 288.080 ;
        RECT 2504.310 288.020 2504.630 288.080 ;
        RECT 2504.310 17.920 2504.630 17.980 ;
        RECT 2504.310 17.780 2645.760 17.920 ;
        RECT 2504.310 17.720 2504.630 17.780 ;
        RECT 2645.620 17.580 2645.760 17.780 ;
        RECT 2672.670 17.580 2672.990 17.640 ;
        RECT 2645.620 17.440 2672.990 17.580 ;
        RECT 2672.670 17.380 2672.990 17.440 ;
      LAYER via ;
        RECT 2498.820 288.020 2499.080 288.280 ;
        RECT 2504.340 288.020 2504.600 288.280 ;
        RECT 2504.340 17.720 2504.600 17.980 ;
        RECT 2672.700 17.380 2672.960 17.640 ;
      LAYER met2 ;
        RECT 2498.820 300.000 2499.100 304.000 ;
        RECT 2498.880 288.310 2499.020 300.000 ;
        RECT 2498.820 287.990 2499.080 288.310 ;
        RECT 2504.340 287.990 2504.600 288.310 ;
        RECT 2504.400 18.010 2504.540 287.990 ;
        RECT 2504.340 17.690 2504.600 18.010 ;
        RECT 2672.700 17.350 2672.960 17.670 ;
        RECT 2672.760 2.400 2672.900 17.350 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2664.465 17.765 2664.635 19.975 ;
      LAYER mcon ;
        RECT 2664.465 19.805 2664.635 19.975 ;
      LAYER met1 ;
        RECT 2513.510 288.220 2513.830 288.280 ;
        RECT 2518.110 288.220 2518.430 288.280 ;
        RECT 2513.510 288.080 2518.430 288.220 ;
        RECT 2513.510 288.020 2513.830 288.080 ;
        RECT 2518.110 288.020 2518.430 288.080 ;
        RECT 2518.110 20.300 2518.430 20.360 ;
        RECT 2518.110 20.160 2655.880 20.300 ;
        RECT 2518.110 20.100 2518.430 20.160 ;
        RECT 2655.740 19.960 2655.880 20.160 ;
        RECT 2664.405 19.960 2664.695 20.005 ;
        RECT 2655.740 19.820 2664.695 19.960 ;
        RECT 2664.405 19.775 2664.695 19.820 ;
        RECT 2664.405 17.920 2664.695 17.965 ;
        RECT 2664.405 17.780 2673.360 17.920 ;
        RECT 2664.405 17.735 2664.695 17.780 ;
        RECT 2673.220 17.580 2673.360 17.780 ;
        RECT 2673.220 17.440 2679.340 17.580 ;
        RECT 2679.200 17.240 2679.340 17.440 ;
        RECT 2690.150 17.240 2690.470 17.300 ;
        RECT 2679.200 17.100 2690.470 17.240 ;
        RECT 2690.150 17.040 2690.470 17.100 ;
      LAYER via ;
        RECT 2513.540 288.020 2513.800 288.280 ;
        RECT 2518.140 288.020 2518.400 288.280 ;
        RECT 2518.140 20.100 2518.400 20.360 ;
        RECT 2690.180 17.040 2690.440 17.300 ;
      LAYER met2 ;
        RECT 2513.540 300.000 2513.820 304.000 ;
        RECT 2513.600 288.310 2513.740 300.000 ;
        RECT 2513.540 287.990 2513.800 288.310 ;
        RECT 2518.140 287.990 2518.400 288.310 ;
        RECT 2518.200 20.390 2518.340 287.990 ;
        RECT 2518.140 20.070 2518.400 20.390 ;
        RECT 2690.180 17.010 2690.440 17.330 ;
        RECT 2690.240 16.730 2690.380 17.010 ;
        RECT 2690.240 16.590 2690.840 16.730 ;
        RECT 2690.700 2.400 2690.840 16.590 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2528.230 288.220 2528.550 288.280 ;
        RECT 2531.910 288.220 2532.230 288.280 ;
        RECT 2528.230 288.080 2532.230 288.220 ;
        RECT 2528.230 288.020 2528.550 288.080 ;
        RECT 2531.910 288.020 2532.230 288.080 ;
        RECT 2531.910 15.880 2532.230 15.940 ;
        RECT 2708.550 15.880 2708.870 15.940 ;
        RECT 2531.910 15.740 2708.870 15.880 ;
        RECT 2531.910 15.680 2532.230 15.740 ;
        RECT 2708.550 15.680 2708.870 15.740 ;
      LAYER via ;
        RECT 2528.260 288.020 2528.520 288.280 ;
        RECT 2531.940 288.020 2532.200 288.280 ;
        RECT 2531.940 15.680 2532.200 15.940 ;
        RECT 2708.580 15.680 2708.840 15.940 ;
      LAYER met2 ;
        RECT 2528.260 300.000 2528.540 304.000 ;
        RECT 2528.320 288.310 2528.460 300.000 ;
        RECT 2528.260 287.990 2528.520 288.310 ;
        RECT 2531.940 287.990 2532.200 288.310 ;
        RECT 2532.000 15.970 2532.140 287.990 ;
        RECT 2531.940 15.650 2532.200 15.970 ;
        RECT 2708.580 15.650 2708.840 15.970 ;
        RECT 2708.640 2.400 2708.780 15.650 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2545.710 15.540 2546.030 15.600 ;
        RECT 2726.490 15.540 2726.810 15.600 ;
        RECT 2545.710 15.400 2726.810 15.540 ;
        RECT 2545.710 15.340 2546.030 15.400 ;
        RECT 2726.490 15.340 2726.810 15.400 ;
      LAYER via ;
        RECT 2545.740 15.340 2546.000 15.600 ;
        RECT 2726.520 15.340 2726.780 15.600 ;
      LAYER met2 ;
        RECT 2542.980 300.290 2543.260 304.000 ;
        RECT 2542.980 300.150 2545.940 300.290 ;
        RECT 2542.980 300.000 2543.260 300.150 ;
        RECT 2545.800 15.630 2545.940 300.150 ;
        RECT 2545.740 15.310 2546.000 15.630 ;
        RECT 2726.520 15.310 2726.780 15.630 ;
        RECT 2726.580 2.400 2726.720 15.310 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2559.510 15.200 2559.830 15.260 ;
        RECT 2744.430 15.200 2744.750 15.260 ;
        RECT 2559.510 15.060 2744.750 15.200 ;
        RECT 2559.510 15.000 2559.830 15.060 ;
        RECT 2744.430 15.000 2744.750 15.060 ;
      LAYER via ;
        RECT 2559.540 15.000 2559.800 15.260 ;
        RECT 2744.460 15.000 2744.720 15.260 ;
      LAYER met2 ;
        RECT 2557.700 300.290 2557.980 304.000 ;
        RECT 2557.700 300.150 2559.740 300.290 ;
        RECT 2557.700 300.000 2557.980 300.150 ;
        RECT 2559.600 15.290 2559.740 300.150 ;
        RECT 2559.540 14.970 2559.800 15.290 ;
        RECT 2744.460 14.970 2744.720 15.290 ;
        RECT 2744.520 2.400 2744.660 14.970 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2573.310 20.640 2573.630 20.700 ;
        RECT 2761.910 20.640 2762.230 20.700 ;
        RECT 2573.310 20.500 2762.230 20.640 ;
        RECT 2573.310 20.440 2573.630 20.500 ;
        RECT 2761.910 20.440 2762.230 20.500 ;
      LAYER via ;
        RECT 2573.340 20.440 2573.600 20.700 ;
        RECT 2761.940 20.440 2762.200 20.700 ;
      LAYER met2 ;
        RECT 2572.420 300.290 2572.700 304.000 ;
        RECT 2572.420 300.150 2573.540 300.290 ;
        RECT 2572.420 300.000 2572.700 300.150 ;
        RECT 2573.400 20.730 2573.540 300.150 ;
        RECT 2573.340 20.410 2573.600 20.730 ;
        RECT 2761.940 20.410 2762.200 20.730 ;
        RECT 2762.000 2.400 2762.140 20.410 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 841.410 284.140 841.730 284.200 ;
        RECT 985.390 284.140 985.710 284.200 ;
        RECT 841.410 284.000 985.710 284.140 ;
        RECT 841.410 283.940 841.730 284.000 ;
        RECT 985.390 283.940 985.710 284.000 ;
        RECT 835.430 15.880 835.750 15.940 ;
        RECT 841.410 15.880 841.730 15.940 ;
        RECT 835.430 15.740 841.730 15.880 ;
        RECT 835.430 15.680 835.750 15.740 ;
        RECT 841.410 15.680 841.730 15.740 ;
      LAYER via ;
        RECT 841.440 283.940 841.700 284.200 ;
        RECT 985.420 283.940 985.680 284.200 ;
        RECT 835.460 15.680 835.720 15.940 ;
        RECT 841.440 15.680 841.700 15.940 ;
      LAYER met2 ;
        RECT 985.420 300.000 985.700 304.000 ;
        RECT 985.480 284.230 985.620 300.000 ;
        RECT 841.440 283.910 841.700 284.230 ;
        RECT 985.420 283.910 985.680 284.230 ;
        RECT 841.500 15.970 841.640 283.910 ;
        RECT 835.460 15.650 835.720 15.970 ;
        RECT 841.440 15.650 841.700 15.970 ;
        RECT 835.520 2.400 835.660 15.650 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2749.105 15.045 2749.275 16.915 ;
      LAYER mcon ;
        RECT 2749.105 16.745 2749.275 16.915 ;
      LAYER met1 ;
        RECT 2587.110 16.900 2587.430 16.960 ;
        RECT 2749.045 16.900 2749.335 16.945 ;
        RECT 2587.110 16.760 2749.335 16.900 ;
        RECT 2587.110 16.700 2587.430 16.760 ;
        RECT 2749.045 16.715 2749.335 16.760 ;
        RECT 2749.045 15.200 2749.335 15.245 ;
        RECT 2779.850 15.200 2780.170 15.260 ;
        RECT 2749.045 15.060 2780.170 15.200 ;
        RECT 2749.045 15.015 2749.335 15.060 ;
        RECT 2779.850 15.000 2780.170 15.060 ;
      LAYER via ;
        RECT 2587.140 16.700 2587.400 16.960 ;
        RECT 2779.880 15.000 2780.140 15.260 ;
      LAYER met2 ;
        RECT 2587.140 300.000 2587.420 304.000 ;
        RECT 2587.200 16.990 2587.340 300.000 ;
        RECT 2587.140 16.670 2587.400 16.990 ;
        RECT 2779.880 14.970 2780.140 15.290 ;
        RECT 2779.940 2.400 2780.080 14.970 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2601.830 289.240 2602.150 289.300 ;
        RECT 2607.810 289.240 2608.130 289.300 ;
        RECT 2601.830 289.100 2608.130 289.240 ;
        RECT 2601.830 289.040 2602.150 289.100 ;
        RECT 2607.810 289.040 2608.130 289.100 ;
        RECT 2606.890 27.440 2607.210 27.500 ;
        RECT 2607.810 27.440 2608.130 27.500 ;
        RECT 2606.890 27.300 2608.130 27.440 ;
        RECT 2606.890 27.240 2607.210 27.300 ;
        RECT 2607.810 27.240 2608.130 27.300 ;
        RECT 2606.890 16.220 2607.210 16.280 ;
        RECT 2797.790 16.220 2798.110 16.280 ;
        RECT 2606.890 16.080 2798.110 16.220 ;
        RECT 2606.890 16.020 2607.210 16.080 ;
        RECT 2797.790 16.020 2798.110 16.080 ;
      LAYER via ;
        RECT 2601.860 289.040 2602.120 289.300 ;
        RECT 2607.840 289.040 2608.100 289.300 ;
        RECT 2606.920 27.240 2607.180 27.500 ;
        RECT 2607.840 27.240 2608.100 27.500 ;
        RECT 2606.920 16.020 2607.180 16.280 ;
        RECT 2797.820 16.020 2798.080 16.280 ;
      LAYER met2 ;
        RECT 2601.860 300.000 2602.140 304.000 ;
        RECT 2601.920 289.330 2602.060 300.000 ;
        RECT 2601.860 289.010 2602.120 289.330 ;
        RECT 2607.840 289.010 2608.100 289.330 ;
        RECT 2607.900 27.530 2608.040 289.010 ;
        RECT 2606.920 27.210 2607.180 27.530 ;
        RECT 2607.840 27.210 2608.100 27.530 ;
        RECT 2606.980 16.310 2607.120 27.210 ;
        RECT 2606.920 15.990 2607.180 16.310 ;
        RECT 2797.820 15.990 2798.080 16.310 ;
        RECT 2797.880 2.400 2798.020 15.990 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2664.925 19.125 2665.095 19.975 ;
      LAYER mcon ;
        RECT 2664.925 19.805 2665.095 19.975 ;
      LAYER met1 ;
        RECT 2616.550 283.460 2616.870 283.520 ;
        RECT 2621.610 283.460 2621.930 283.520 ;
        RECT 2616.550 283.320 2621.930 283.460 ;
        RECT 2616.550 283.260 2616.870 283.320 ;
        RECT 2621.610 283.260 2621.930 283.320 ;
        RECT 2664.865 19.960 2665.155 20.005 ;
        RECT 2815.730 19.960 2816.050 20.020 ;
        RECT 2664.865 19.820 2816.050 19.960 ;
        RECT 2664.865 19.775 2665.155 19.820 ;
        RECT 2815.730 19.760 2816.050 19.820 ;
        RECT 2621.610 19.280 2621.930 19.340 ;
        RECT 2664.865 19.280 2665.155 19.325 ;
        RECT 2621.610 19.140 2665.155 19.280 ;
        RECT 2621.610 19.080 2621.930 19.140 ;
        RECT 2664.865 19.095 2665.155 19.140 ;
      LAYER via ;
        RECT 2616.580 283.260 2616.840 283.520 ;
        RECT 2621.640 283.260 2621.900 283.520 ;
        RECT 2815.760 19.760 2816.020 20.020 ;
        RECT 2621.640 19.080 2621.900 19.340 ;
      LAYER met2 ;
        RECT 2616.580 300.000 2616.860 304.000 ;
        RECT 2616.640 283.550 2616.780 300.000 ;
        RECT 2616.580 283.230 2616.840 283.550 ;
        RECT 2621.640 283.230 2621.900 283.550 ;
        RECT 2621.700 19.370 2621.840 283.230 ;
        RECT 2815.760 19.730 2816.020 20.050 ;
        RECT 2621.640 19.050 2621.900 19.370 ;
        RECT 2815.820 2.400 2815.960 19.730 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2630.810 285.500 2631.130 285.560 ;
        RECT 2666.690 285.500 2667.010 285.560 ;
        RECT 2630.810 285.360 2667.010 285.500 ;
        RECT 2630.810 285.300 2631.130 285.360 ;
        RECT 2666.690 285.300 2667.010 285.360 ;
        RECT 2666.690 14.860 2667.010 14.920 ;
        RECT 2666.690 14.720 2715.220 14.860 ;
        RECT 2666.690 14.660 2667.010 14.720 ;
        RECT 2715.080 14.520 2715.220 14.720 ;
        RECT 2833.670 14.520 2833.990 14.580 ;
        RECT 2715.080 14.380 2833.990 14.520 ;
        RECT 2833.670 14.320 2833.990 14.380 ;
      LAYER via ;
        RECT 2630.840 285.300 2631.100 285.560 ;
        RECT 2666.720 285.300 2666.980 285.560 ;
        RECT 2666.720 14.660 2666.980 14.920 ;
        RECT 2833.700 14.320 2833.960 14.580 ;
      LAYER met2 ;
        RECT 2630.840 300.000 2631.120 304.000 ;
        RECT 2630.900 285.590 2631.040 300.000 ;
        RECT 2630.840 285.270 2631.100 285.590 ;
        RECT 2666.720 285.270 2666.980 285.590 ;
        RECT 2666.780 14.950 2666.920 285.270 ;
        RECT 2666.720 14.630 2666.980 14.950 ;
        RECT 2833.700 14.290 2833.960 14.610 ;
        RECT 2833.760 2.400 2833.900 14.290 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2645.530 285.840 2645.850 285.900 ;
        RECT 2687.390 285.840 2687.710 285.900 ;
        RECT 2645.530 285.700 2687.710 285.840 ;
        RECT 2645.530 285.640 2645.850 285.700 ;
        RECT 2687.390 285.640 2687.710 285.700 ;
        RECT 2687.390 14.520 2687.710 14.580 ;
        RECT 2687.390 14.380 2713.840 14.520 ;
        RECT 2687.390 14.320 2687.710 14.380 ;
        RECT 2713.700 14.180 2713.840 14.380 ;
        RECT 2851.150 14.180 2851.470 14.240 ;
        RECT 2713.700 14.040 2851.470 14.180 ;
        RECT 2851.150 13.980 2851.470 14.040 ;
      LAYER via ;
        RECT 2645.560 285.640 2645.820 285.900 ;
        RECT 2687.420 285.640 2687.680 285.900 ;
        RECT 2687.420 14.320 2687.680 14.580 ;
        RECT 2851.180 13.980 2851.440 14.240 ;
      LAYER met2 ;
        RECT 2645.560 300.000 2645.840 304.000 ;
        RECT 2645.620 285.930 2645.760 300.000 ;
        RECT 2645.560 285.610 2645.820 285.930 ;
        RECT 2687.420 285.610 2687.680 285.930 ;
        RECT 2687.480 14.610 2687.620 285.610 ;
        RECT 2687.420 14.290 2687.680 14.610 ;
        RECT 2851.180 13.950 2851.440 14.270 ;
        RECT 2851.240 2.400 2851.380 13.950 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2663.010 18.260 2663.330 18.320 ;
        RECT 2869.090 18.260 2869.410 18.320 ;
        RECT 2663.010 18.120 2869.410 18.260 ;
        RECT 2663.010 18.060 2663.330 18.120 ;
        RECT 2869.090 18.060 2869.410 18.120 ;
      LAYER via ;
        RECT 2663.040 18.060 2663.300 18.320 ;
        RECT 2869.120 18.060 2869.380 18.320 ;
      LAYER met2 ;
        RECT 2660.280 300.290 2660.560 304.000 ;
        RECT 2660.280 300.150 2663.240 300.290 ;
        RECT 2660.280 300.000 2660.560 300.150 ;
        RECT 2663.100 18.350 2663.240 300.150 ;
        RECT 2663.040 18.030 2663.300 18.350 ;
        RECT 2869.120 18.030 2869.380 18.350 ;
        RECT 2869.180 2.400 2869.320 18.030 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2674.970 284.820 2675.290 284.880 ;
        RECT 2694.750 284.820 2695.070 284.880 ;
        RECT 2674.970 284.680 2695.070 284.820 ;
        RECT 2674.970 284.620 2675.290 284.680 ;
        RECT 2694.750 284.620 2695.070 284.680 ;
        RECT 2694.750 20.300 2695.070 20.360 ;
        RECT 2887.030 20.300 2887.350 20.360 ;
        RECT 2694.750 20.160 2887.350 20.300 ;
        RECT 2694.750 20.100 2695.070 20.160 ;
        RECT 2887.030 20.100 2887.350 20.160 ;
      LAYER via ;
        RECT 2675.000 284.620 2675.260 284.880 ;
        RECT 2694.780 284.620 2695.040 284.880 ;
        RECT 2694.780 20.100 2695.040 20.360 ;
        RECT 2887.060 20.100 2887.320 20.360 ;
      LAYER met2 ;
        RECT 2675.000 300.000 2675.280 304.000 ;
        RECT 2675.060 284.910 2675.200 300.000 ;
        RECT 2675.000 284.590 2675.260 284.910 ;
        RECT 2694.780 284.590 2695.040 284.910 ;
        RECT 2694.840 20.390 2694.980 284.590 ;
        RECT 2694.780 20.070 2695.040 20.390 ;
        RECT 2887.060 20.070 2887.320 20.390 ;
        RECT 2887.120 2.400 2887.260 20.070 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2689.690 283.120 2690.010 283.180 ;
        RECT 2701.190 283.120 2701.510 283.180 ;
        RECT 2689.690 282.980 2701.510 283.120 ;
        RECT 2689.690 282.920 2690.010 282.980 ;
        RECT 2701.190 282.920 2701.510 282.980 ;
      LAYER via ;
        RECT 2689.720 282.920 2689.980 283.180 ;
        RECT 2701.220 282.920 2701.480 283.180 ;
      LAYER met2 ;
        RECT 2689.720 300.000 2690.000 304.000 ;
        RECT 2689.780 283.210 2689.920 300.000 ;
        RECT 2689.720 282.890 2689.980 283.210 ;
        RECT 2701.220 282.890 2701.480 283.210 ;
        RECT 2701.280 16.845 2701.420 282.890 ;
        RECT 2701.210 16.475 2701.490 16.845 ;
        RECT 2904.990 16.475 2905.270 16.845 ;
        RECT 2905.060 2.400 2905.200 16.475 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 2701.210 16.520 2701.490 16.800 ;
        RECT 2904.990 16.520 2905.270 16.800 ;
      LAYER met3 ;
        RECT 2701.185 16.810 2701.515 16.825 ;
        RECT 2904.965 16.810 2905.295 16.825 ;
        RECT 2701.185 16.510 2905.295 16.810 ;
        RECT 2701.185 16.495 2701.515 16.510 ;
        RECT 2904.965 16.495 2905.295 16.510 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 855.210 283.800 855.530 283.860 ;
        RECT 998.270 283.800 998.590 283.860 ;
        RECT 855.210 283.660 998.590 283.800 ;
        RECT 855.210 283.600 855.530 283.660 ;
        RECT 998.270 283.600 998.590 283.660 ;
        RECT 852.910 15.200 853.230 15.260 ;
        RECT 855.210 15.200 855.530 15.260 ;
        RECT 852.910 15.060 855.530 15.200 ;
        RECT 852.910 15.000 853.230 15.060 ;
        RECT 855.210 15.000 855.530 15.060 ;
      LAYER via ;
        RECT 855.240 283.600 855.500 283.860 ;
        RECT 998.300 283.600 998.560 283.860 ;
        RECT 852.940 15.000 853.200 15.260 ;
        RECT 855.240 15.000 855.500 15.260 ;
      LAYER met2 ;
        RECT 1000.140 300.290 1000.420 304.000 ;
        RECT 998.360 300.150 1000.420 300.290 ;
        RECT 998.360 283.890 998.500 300.150 ;
        RECT 1000.140 300.000 1000.420 300.150 ;
        RECT 855.240 283.570 855.500 283.890 ;
        RECT 998.300 283.570 998.560 283.890 ;
        RECT 855.300 15.290 855.440 283.570 ;
        RECT 852.940 14.970 853.200 15.290 ;
        RECT 855.240 14.970 855.500 15.290 ;
        RECT 853.000 2.400 853.140 14.970 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 927.965 286.705 928.135 287.555 ;
      LAYER mcon ;
        RECT 927.965 287.385 928.135 287.555 ;
      LAYER met1 ;
        RECT 927.905 287.540 928.195 287.585 ;
        RECT 887.960 287.400 928.195 287.540 ;
        RECT 875.910 287.200 876.230 287.260 ;
        RECT 887.960 287.200 888.100 287.400 ;
        RECT 927.905 287.355 928.195 287.400 ;
        RECT 875.910 287.060 888.100 287.200 ;
        RECT 875.910 287.000 876.230 287.060 ;
        RECT 927.905 286.860 928.195 286.905 ;
        RECT 1014.830 286.860 1015.150 286.920 ;
        RECT 927.905 286.720 1015.150 286.860 ;
        RECT 927.905 286.675 928.195 286.720 ;
        RECT 1014.830 286.660 1015.150 286.720 ;
        RECT 870.850 16.900 871.170 16.960 ;
        RECT 875.910 16.900 876.230 16.960 ;
        RECT 870.850 16.760 876.230 16.900 ;
        RECT 870.850 16.700 871.170 16.760 ;
        RECT 875.910 16.700 876.230 16.760 ;
      LAYER via ;
        RECT 875.940 287.000 876.200 287.260 ;
        RECT 1014.860 286.660 1015.120 286.920 ;
        RECT 870.880 16.700 871.140 16.960 ;
        RECT 875.940 16.700 876.200 16.960 ;
      LAYER met2 ;
        RECT 1014.860 300.000 1015.140 304.000 ;
        RECT 875.940 286.970 876.200 287.290 ;
        RECT 876.000 16.990 876.140 286.970 ;
        RECT 1014.920 286.950 1015.060 300.000 ;
        RECT 1014.860 286.630 1015.120 286.950 ;
        RECT 870.880 16.670 871.140 16.990 ;
        RECT 875.940 16.670 876.200 16.990 ;
        RECT 870.940 2.400 871.080 16.670 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 889.710 287.200 890.030 287.260 ;
        RECT 1029.550 287.200 1029.870 287.260 ;
        RECT 889.710 287.060 1029.870 287.200 ;
        RECT 889.710 287.000 890.030 287.060 ;
        RECT 1029.550 287.000 1029.870 287.060 ;
      LAYER via ;
        RECT 889.740 287.000 890.000 287.260 ;
        RECT 1029.580 287.000 1029.840 287.260 ;
      LAYER met2 ;
        RECT 1029.580 300.000 1029.860 304.000 ;
        RECT 1029.640 287.290 1029.780 300.000 ;
        RECT 889.740 286.970 890.000 287.290 ;
        RECT 1029.580 286.970 1029.840 287.290 ;
        RECT 889.800 16.730 889.940 286.970 ;
        RECT 888.880 16.590 889.940 16.730 ;
        RECT 888.880 2.400 889.020 16.590 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 955.565 287.725 955.735 288.575 ;
      LAYER mcon ;
        RECT 955.565 288.405 955.735 288.575 ;
      LAYER met1 ;
        RECT 910.410 288.560 910.730 288.620 ;
        RECT 955.505 288.560 955.795 288.605 ;
        RECT 910.410 288.420 955.795 288.560 ;
        RECT 910.410 288.360 910.730 288.420 ;
        RECT 955.505 288.375 955.795 288.420 ;
        RECT 955.505 287.880 955.795 287.925 ;
        RECT 1044.270 287.880 1044.590 287.940 ;
        RECT 955.505 287.740 1044.590 287.880 ;
        RECT 955.505 287.695 955.795 287.740 ;
        RECT 1044.270 287.680 1044.590 287.740 ;
        RECT 906.730 16.900 907.050 16.960 ;
        RECT 910.410 16.900 910.730 16.960 ;
        RECT 906.730 16.760 910.730 16.900 ;
        RECT 906.730 16.700 907.050 16.760 ;
        RECT 910.410 16.700 910.730 16.760 ;
      LAYER via ;
        RECT 910.440 288.360 910.700 288.620 ;
        RECT 1044.300 287.680 1044.560 287.940 ;
        RECT 906.760 16.700 907.020 16.960 ;
        RECT 910.440 16.700 910.700 16.960 ;
      LAYER met2 ;
        RECT 1044.300 300.000 1044.580 304.000 ;
        RECT 910.440 288.330 910.700 288.650 ;
        RECT 910.500 16.990 910.640 288.330 ;
        RECT 1044.360 287.970 1044.500 300.000 ;
        RECT 1044.300 287.650 1044.560 287.970 ;
        RECT 906.760 16.670 907.020 16.990 ;
        RECT 910.440 16.670 910.700 16.990 ;
        RECT 906.820 2.400 906.960 16.670 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 955.105 285.005 955.275 287.895 ;
        RECT 979.485 285.005 979.655 287.555 ;
      LAYER mcon ;
        RECT 955.105 287.725 955.275 287.895 ;
        RECT 979.485 287.385 979.655 287.555 ;
      LAYER met1 ;
        RECT 924.210 287.880 924.530 287.940 ;
        RECT 955.045 287.880 955.335 287.925 ;
        RECT 924.210 287.740 955.335 287.880 ;
        RECT 924.210 287.680 924.530 287.740 ;
        RECT 955.045 287.695 955.335 287.740 ;
        RECT 979.425 287.540 979.715 287.585 ;
        RECT 1058.990 287.540 1059.310 287.600 ;
        RECT 979.425 287.400 1059.310 287.540 ;
        RECT 979.425 287.355 979.715 287.400 ;
        RECT 1058.990 287.340 1059.310 287.400 ;
        RECT 955.045 285.160 955.335 285.205 ;
        RECT 979.425 285.160 979.715 285.205 ;
        RECT 955.045 285.020 979.715 285.160 ;
        RECT 955.045 284.975 955.335 285.020 ;
        RECT 979.425 284.975 979.715 285.020 ;
      LAYER via ;
        RECT 924.240 287.680 924.500 287.940 ;
        RECT 1059.020 287.340 1059.280 287.600 ;
      LAYER met2 ;
        RECT 1059.020 300.000 1059.300 304.000 ;
        RECT 924.240 287.650 924.500 287.970 ;
        RECT 924.300 2.400 924.440 287.650 ;
        RECT 1059.080 287.630 1059.220 300.000 ;
        RECT 1059.020 287.310 1059.280 287.630 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 956.485 285.685 956.655 289.255 ;
      LAYER mcon ;
        RECT 956.485 289.085 956.655 289.255 ;
      LAYER met1 ;
        RECT 956.425 289.240 956.715 289.285 ;
        RECT 1073.710 289.240 1074.030 289.300 ;
        RECT 956.425 289.100 1074.030 289.240 ;
        RECT 956.425 289.055 956.715 289.100 ;
        RECT 1073.710 289.040 1074.030 289.100 ;
        RECT 944.910 285.840 945.230 285.900 ;
        RECT 956.425 285.840 956.715 285.885 ;
        RECT 944.910 285.700 956.715 285.840 ;
        RECT 944.910 285.640 945.230 285.700 ;
        RECT 956.425 285.655 956.715 285.700 ;
        RECT 942.150 15.200 942.470 15.260 ;
        RECT 944.910 15.200 945.230 15.260 ;
        RECT 942.150 15.060 945.230 15.200 ;
        RECT 942.150 15.000 942.470 15.060 ;
        RECT 944.910 15.000 945.230 15.060 ;
      LAYER via ;
        RECT 1073.740 289.040 1074.000 289.300 ;
        RECT 944.940 285.640 945.200 285.900 ;
        RECT 942.180 15.000 942.440 15.260 ;
        RECT 944.940 15.000 945.200 15.260 ;
      LAYER met2 ;
        RECT 1073.740 300.000 1074.020 304.000 ;
        RECT 1073.800 289.330 1073.940 300.000 ;
        RECT 1073.740 289.010 1074.000 289.330 ;
        RECT 944.940 285.610 945.200 285.930 ;
        RECT 945.000 15.290 945.140 285.610 ;
        RECT 942.180 14.970 942.440 15.290 ;
        RECT 944.940 14.970 945.200 15.290 ;
        RECT 942.240 2.400 942.380 14.970 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 965.610 285.500 965.930 285.560 ;
        RECT 1088.430 285.500 1088.750 285.560 ;
        RECT 965.610 285.360 1088.750 285.500 ;
        RECT 965.610 285.300 965.930 285.360 ;
        RECT 1088.430 285.300 1088.750 285.360 ;
        RECT 960.090 16.900 960.410 16.960 ;
        RECT 965.610 16.900 965.930 16.960 ;
        RECT 960.090 16.760 965.930 16.900 ;
        RECT 960.090 16.700 960.410 16.760 ;
        RECT 965.610 16.700 965.930 16.760 ;
      LAYER via ;
        RECT 965.640 285.300 965.900 285.560 ;
        RECT 1088.460 285.300 1088.720 285.560 ;
        RECT 960.120 16.700 960.380 16.960 ;
        RECT 965.640 16.700 965.900 16.960 ;
      LAYER met2 ;
        RECT 1088.460 300.000 1088.740 304.000 ;
        RECT 1088.520 285.590 1088.660 300.000 ;
        RECT 965.640 285.270 965.900 285.590 ;
        RECT 1088.460 285.270 1088.720 285.590 ;
        RECT 965.700 16.990 965.840 285.270 ;
        RECT 960.120 16.670 960.380 16.990 ;
        RECT 965.640 16.670 965.900 16.990 ;
        RECT 960.180 2.400 960.320 16.670 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 979.945 241.485 980.115 285.855 ;
        RECT 979.485 144.925 979.655 193.035 ;
        RECT 978.105 2.805 978.275 48.195 ;
      LAYER mcon ;
        RECT 979.945 285.685 980.115 285.855 ;
        RECT 979.485 192.865 979.655 193.035 ;
        RECT 978.105 48.025 978.275 48.195 ;
      LAYER met1 ;
        RECT 979.885 285.840 980.175 285.885 ;
        RECT 1103.150 285.840 1103.470 285.900 ;
        RECT 979.885 285.700 1103.470 285.840 ;
        RECT 979.885 285.655 980.175 285.700 ;
        RECT 1103.150 285.640 1103.470 285.700 ;
        RECT 979.410 241.640 979.730 241.700 ;
        RECT 979.885 241.640 980.175 241.685 ;
        RECT 979.410 241.500 980.175 241.640 ;
        RECT 979.410 241.440 979.730 241.500 ;
        RECT 979.885 241.455 980.175 241.500 ;
        RECT 979.410 193.020 979.730 193.080 ;
        RECT 979.215 192.880 979.730 193.020 ;
        RECT 979.410 192.820 979.730 192.880 ;
        RECT 979.410 145.080 979.730 145.140 ;
        RECT 979.215 144.940 979.730 145.080 ;
        RECT 979.410 144.880 979.730 144.940 ;
        RECT 979.410 97.280 979.730 97.540 ;
        RECT 979.500 96.860 979.640 97.280 ;
        RECT 979.410 96.600 979.730 96.860 ;
        RECT 978.045 48.180 978.335 48.225 ;
        RECT 979.410 48.180 979.730 48.240 ;
        RECT 978.045 48.040 979.730 48.180 ;
        RECT 978.045 47.995 978.335 48.040 ;
        RECT 979.410 47.980 979.730 48.040 ;
        RECT 978.030 2.960 978.350 3.020 ;
        RECT 977.835 2.820 978.350 2.960 ;
        RECT 978.030 2.760 978.350 2.820 ;
      LAYER via ;
        RECT 1103.180 285.640 1103.440 285.900 ;
        RECT 979.440 241.440 979.700 241.700 ;
        RECT 979.440 192.820 979.700 193.080 ;
        RECT 979.440 144.880 979.700 145.140 ;
        RECT 979.440 97.280 979.700 97.540 ;
        RECT 979.440 96.600 979.700 96.860 ;
        RECT 979.440 47.980 979.700 48.240 ;
        RECT 978.060 2.760 978.320 3.020 ;
      LAYER met2 ;
        RECT 1103.180 300.000 1103.460 304.000 ;
        RECT 1103.240 285.930 1103.380 300.000 ;
        RECT 1103.180 285.610 1103.440 285.930 ;
        RECT 979.440 241.410 979.700 241.730 ;
        RECT 979.500 193.110 979.640 241.410 ;
        RECT 979.440 192.790 979.700 193.110 ;
        RECT 979.440 144.850 979.700 145.170 ;
        RECT 979.500 97.570 979.640 144.850 ;
        RECT 979.440 97.250 979.700 97.570 ;
        RECT 979.440 96.570 979.700 96.890 ;
        RECT 979.500 96.405 979.640 96.570 ;
        RECT 979.430 96.035 979.710 96.405 ;
        RECT 980.810 96.035 981.090 96.405 ;
        RECT 980.880 48.805 981.020 96.035 ;
        RECT 979.430 48.435 979.710 48.805 ;
        RECT 980.810 48.435 981.090 48.805 ;
        RECT 979.500 48.270 979.640 48.435 ;
        RECT 979.440 47.950 979.700 48.270 ;
        RECT 978.060 2.730 978.320 3.050 ;
        RECT 978.120 2.400 978.260 2.730 ;
        RECT 977.910 -4.800 978.470 2.400 ;
      LAYER via2 ;
        RECT 979.430 96.080 979.710 96.360 ;
        RECT 980.810 96.080 981.090 96.360 ;
        RECT 979.430 48.480 979.710 48.760 ;
        RECT 980.810 48.480 981.090 48.760 ;
      LAYER met3 ;
        RECT 979.405 96.370 979.735 96.385 ;
        RECT 980.785 96.370 981.115 96.385 ;
        RECT 979.405 96.070 981.115 96.370 ;
        RECT 979.405 96.055 979.735 96.070 ;
        RECT 980.785 96.055 981.115 96.070 ;
        RECT 979.405 48.770 979.735 48.785 ;
        RECT 980.785 48.770 981.115 48.785 ;
        RECT 979.405 48.470 981.115 48.770 ;
        RECT 979.405 48.455 979.735 48.470 ;
        RECT 980.785 48.455 981.115 48.470 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 25.060 657.270 25.120 ;
        RECT 834.970 25.060 835.290 25.120 ;
        RECT 656.950 24.920 835.290 25.060 ;
        RECT 656.950 24.860 657.270 24.920 ;
        RECT 834.970 24.860 835.290 24.920 ;
      LAYER via ;
        RECT 656.980 24.860 657.240 25.120 ;
        RECT 835.000 24.860 835.260 25.120 ;
      LAYER met2 ;
        RECT 838.680 300.290 838.960 304.000 ;
        RECT 835.060 300.150 838.960 300.290 ;
        RECT 835.060 25.150 835.200 300.150 ;
        RECT 838.680 300.000 838.960 300.150 ;
        RECT 656.980 24.830 657.240 25.150 ;
        RECT 835.000 24.830 835.260 25.150 ;
        RECT 657.040 2.400 657.180 24.830 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1000.110 286.520 1000.430 286.580 ;
        RECT 1117.870 286.520 1118.190 286.580 ;
        RECT 1000.110 286.380 1118.190 286.520 ;
        RECT 1000.110 286.320 1000.430 286.380 ;
        RECT 1117.870 286.320 1118.190 286.380 ;
        RECT 995.970 20.640 996.290 20.700 ;
        RECT 1000.110 20.640 1000.430 20.700 ;
        RECT 995.970 20.500 1000.430 20.640 ;
        RECT 995.970 20.440 996.290 20.500 ;
        RECT 1000.110 20.440 1000.430 20.500 ;
      LAYER via ;
        RECT 1000.140 286.320 1000.400 286.580 ;
        RECT 1117.900 286.320 1118.160 286.580 ;
        RECT 996.000 20.440 996.260 20.700 ;
        RECT 1000.140 20.440 1000.400 20.700 ;
      LAYER met2 ;
        RECT 1117.900 300.000 1118.180 304.000 ;
        RECT 1117.960 286.610 1118.100 300.000 ;
        RECT 1000.140 286.290 1000.400 286.610 ;
        RECT 1117.900 286.290 1118.160 286.610 ;
        RECT 1000.200 20.730 1000.340 286.290 ;
        RECT 996.000 20.410 996.260 20.730 ;
        RECT 1000.140 20.410 1000.400 20.730 ;
        RECT 996.060 2.400 996.200 20.410 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1132.160 300.000 1132.440 304.000 ;
        RECT 1132.220 286.125 1132.360 300.000 ;
        RECT 1013.930 285.755 1014.210 286.125 ;
        RECT 1132.150 285.755 1132.430 286.125 ;
        RECT 1014.000 20.130 1014.140 285.755 ;
        RECT 1013.540 19.990 1014.140 20.130 ;
        RECT 1013.540 2.400 1013.680 19.990 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
      LAYER via2 ;
        RECT 1013.930 285.800 1014.210 286.080 ;
        RECT 1132.150 285.800 1132.430 286.080 ;
      LAYER met3 ;
        RECT 1013.905 286.090 1014.235 286.105 ;
        RECT 1132.125 286.090 1132.455 286.105 ;
        RECT 1013.905 285.790 1132.455 286.090 ;
        RECT 1013.905 285.775 1014.235 285.790 ;
        RECT 1132.125 285.775 1132.455 285.790 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1033.690 287.200 1034.010 287.260 ;
        RECT 1146.850 287.200 1147.170 287.260 ;
        RECT 1033.690 287.060 1147.170 287.200 ;
        RECT 1033.690 287.000 1034.010 287.060 ;
        RECT 1146.850 287.000 1147.170 287.060 ;
        RECT 1031.390 15.540 1031.710 15.600 ;
        RECT 1034.610 15.540 1034.930 15.600 ;
        RECT 1031.390 15.400 1034.930 15.540 ;
        RECT 1031.390 15.340 1031.710 15.400 ;
        RECT 1034.610 15.340 1034.930 15.400 ;
      LAYER via ;
        RECT 1033.720 287.000 1033.980 287.260 ;
        RECT 1146.880 287.000 1147.140 287.260 ;
        RECT 1031.420 15.340 1031.680 15.600 ;
        RECT 1034.640 15.340 1034.900 15.600 ;
      LAYER met2 ;
        RECT 1146.880 300.000 1147.160 304.000 ;
        RECT 1146.940 287.290 1147.080 300.000 ;
        RECT 1033.720 286.970 1033.980 287.290 ;
        RECT 1146.880 286.970 1147.140 287.290 ;
        RECT 1033.780 271.050 1033.920 286.970 ;
        RECT 1033.780 270.910 1034.840 271.050 ;
        RECT 1034.700 15.630 1034.840 270.910 ;
        RECT 1031.420 15.310 1031.680 15.630 ;
        RECT 1034.640 15.310 1034.900 15.630 ;
        RECT 1031.480 2.400 1031.620 15.310 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1079.305 282.965 1079.475 288.575 ;
      LAYER mcon ;
        RECT 1079.305 288.405 1079.475 288.575 ;
      LAYER met1 ;
        RECT 1079.245 288.560 1079.535 288.605 ;
        RECT 1161.570 288.560 1161.890 288.620 ;
        RECT 1079.245 288.420 1161.890 288.560 ;
        RECT 1079.245 288.375 1079.535 288.420 ;
        RECT 1161.570 288.360 1161.890 288.420 ;
        RECT 1054.850 283.120 1055.170 283.180 ;
        RECT 1079.245 283.120 1079.535 283.165 ;
        RECT 1054.850 282.980 1079.535 283.120 ;
        RECT 1054.850 282.920 1055.170 282.980 ;
        RECT 1079.245 282.935 1079.535 282.980 ;
        RECT 1049.330 14.860 1049.650 14.920 ;
        RECT 1054.850 14.860 1055.170 14.920 ;
        RECT 1049.330 14.720 1055.170 14.860 ;
        RECT 1049.330 14.660 1049.650 14.720 ;
        RECT 1054.850 14.660 1055.170 14.720 ;
      LAYER via ;
        RECT 1161.600 288.360 1161.860 288.620 ;
        RECT 1054.880 282.920 1055.140 283.180 ;
        RECT 1049.360 14.660 1049.620 14.920 ;
        RECT 1054.880 14.660 1055.140 14.920 ;
      LAYER met2 ;
        RECT 1161.600 300.000 1161.880 304.000 ;
        RECT 1161.660 288.650 1161.800 300.000 ;
        RECT 1161.600 288.330 1161.860 288.650 ;
        RECT 1054.880 282.890 1055.140 283.210 ;
        RECT 1054.940 14.950 1055.080 282.890 ;
        RECT 1049.360 14.630 1049.620 14.950 ;
        RECT 1054.880 14.630 1055.140 14.950 ;
        RECT 1049.420 2.400 1049.560 14.630 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1078.845 288.405 1079.015 289.595 ;
        RECT 1121.165 288.745 1121.335 289.595 ;
        RECT 1067.345 2.805 1067.515 14.195 ;
      LAYER mcon ;
        RECT 1078.845 289.425 1079.015 289.595 ;
        RECT 1121.165 289.425 1121.335 289.595 ;
        RECT 1067.345 14.025 1067.515 14.195 ;
      LAYER met1 ;
        RECT 1078.785 289.580 1079.075 289.625 ;
        RECT 1121.105 289.580 1121.395 289.625 ;
        RECT 1078.785 289.440 1121.395 289.580 ;
        RECT 1078.785 289.395 1079.075 289.440 ;
        RECT 1121.105 289.395 1121.395 289.440 ;
        RECT 1121.105 288.900 1121.395 288.945 ;
        RECT 1176.290 288.900 1176.610 288.960 ;
        RECT 1121.105 288.760 1176.610 288.900 ;
        RECT 1121.105 288.715 1121.395 288.760 ;
        RECT 1176.290 288.700 1176.610 288.760 ;
        RECT 1069.110 288.560 1069.430 288.620 ;
        RECT 1078.785 288.560 1079.075 288.605 ;
        RECT 1069.110 288.420 1079.075 288.560 ;
        RECT 1069.110 288.360 1069.430 288.420 ;
        RECT 1078.785 288.375 1079.075 288.420 ;
        RECT 1067.285 14.180 1067.575 14.225 ;
        RECT 1069.110 14.180 1069.430 14.240 ;
        RECT 1067.285 14.040 1069.430 14.180 ;
        RECT 1067.285 13.995 1067.575 14.040 ;
        RECT 1069.110 13.980 1069.430 14.040 ;
        RECT 1067.270 2.960 1067.590 3.020 ;
        RECT 1067.075 2.820 1067.590 2.960 ;
        RECT 1067.270 2.760 1067.590 2.820 ;
      LAYER via ;
        RECT 1176.320 288.700 1176.580 288.960 ;
        RECT 1069.140 288.360 1069.400 288.620 ;
        RECT 1069.140 13.980 1069.400 14.240 ;
        RECT 1067.300 2.760 1067.560 3.020 ;
      LAYER met2 ;
        RECT 1176.320 300.000 1176.600 304.000 ;
        RECT 1176.380 288.990 1176.520 300.000 ;
        RECT 1176.320 288.670 1176.580 288.990 ;
        RECT 1069.140 288.330 1069.400 288.650 ;
        RECT 1069.200 14.270 1069.340 288.330 ;
        RECT 1069.140 13.950 1069.400 14.270 ;
        RECT 1067.300 2.730 1067.560 3.050 ;
        RECT 1067.360 2.400 1067.500 2.730 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1089.810 285.160 1090.130 285.220 ;
        RECT 1191.010 285.160 1191.330 285.220 ;
        RECT 1089.810 285.020 1191.330 285.160 ;
        RECT 1089.810 284.960 1090.130 285.020 ;
        RECT 1191.010 284.960 1191.330 285.020 ;
        RECT 1085.210 17.580 1085.530 17.640 ;
        RECT 1089.810 17.580 1090.130 17.640 ;
        RECT 1085.210 17.440 1090.130 17.580 ;
        RECT 1085.210 17.380 1085.530 17.440 ;
        RECT 1089.810 17.380 1090.130 17.440 ;
      LAYER via ;
        RECT 1089.840 284.960 1090.100 285.220 ;
        RECT 1191.040 284.960 1191.300 285.220 ;
        RECT 1085.240 17.380 1085.500 17.640 ;
        RECT 1089.840 17.380 1090.100 17.640 ;
      LAYER met2 ;
        RECT 1191.040 300.000 1191.320 304.000 ;
        RECT 1191.100 285.250 1191.240 300.000 ;
        RECT 1089.840 284.930 1090.100 285.250 ;
        RECT 1191.040 284.930 1191.300 285.250 ;
        RECT 1089.900 17.670 1090.040 284.930 ;
        RECT 1085.240 17.350 1085.500 17.670 ;
        RECT 1089.840 17.350 1090.100 17.670 ;
        RECT 1085.300 2.400 1085.440 17.350 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1103.610 285.840 1103.930 285.900 ;
        RECT 1205.730 285.840 1206.050 285.900 ;
        RECT 1103.610 285.700 1206.050 285.840 ;
        RECT 1103.610 285.640 1103.930 285.700 ;
        RECT 1205.730 285.640 1206.050 285.700 ;
      LAYER via ;
        RECT 1103.640 285.640 1103.900 285.900 ;
        RECT 1205.760 285.640 1206.020 285.900 ;
      LAYER met2 ;
        RECT 1205.760 300.000 1206.040 304.000 ;
        RECT 1205.820 285.930 1205.960 300.000 ;
        RECT 1103.640 285.610 1103.900 285.930 ;
        RECT 1205.760 285.610 1206.020 285.930 ;
        RECT 1103.700 17.410 1103.840 285.610 ;
        RECT 1102.780 17.270 1103.840 17.410 ;
        RECT 1102.780 2.400 1102.920 17.270 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1124.310 284.480 1124.630 284.540 ;
        RECT 1220.450 284.480 1220.770 284.540 ;
        RECT 1124.310 284.340 1220.770 284.480 ;
        RECT 1124.310 284.280 1124.630 284.340 ;
        RECT 1220.450 284.280 1220.770 284.340 ;
        RECT 1120.630 15.200 1120.950 15.260 ;
        RECT 1124.310 15.200 1124.630 15.260 ;
        RECT 1120.630 15.060 1124.630 15.200 ;
        RECT 1120.630 15.000 1120.950 15.060 ;
        RECT 1124.310 15.000 1124.630 15.060 ;
      LAYER via ;
        RECT 1124.340 284.280 1124.600 284.540 ;
        RECT 1220.480 284.280 1220.740 284.540 ;
        RECT 1120.660 15.000 1120.920 15.260 ;
        RECT 1124.340 15.000 1124.600 15.260 ;
      LAYER met2 ;
        RECT 1220.480 300.000 1220.760 304.000 ;
        RECT 1220.540 284.570 1220.680 300.000 ;
        RECT 1124.340 284.250 1124.600 284.570 ;
        RECT 1220.480 284.250 1220.740 284.570 ;
        RECT 1124.400 15.290 1124.540 284.250 ;
        RECT 1120.660 14.970 1120.920 15.290 ;
        RECT 1124.340 14.970 1124.600 15.290 ;
        RECT 1120.720 2.400 1120.860 14.970 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1145.010 288.220 1145.330 288.280 ;
        RECT 1235.170 288.220 1235.490 288.280 ;
        RECT 1145.010 288.080 1235.490 288.220 ;
        RECT 1145.010 288.020 1145.330 288.080 ;
        RECT 1235.170 288.020 1235.490 288.080 ;
        RECT 1138.570 17.240 1138.890 17.300 ;
        RECT 1145.010 17.240 1145.330 17.300 ;
        RECT 1138.570 17.100 1145.330 17.240 ;
        RECT 1138.570 17.040 1138.890 17.100 ;
        RECT 1145.010 17.040 1145.330 17.100 ;
      LAYER via ;
        RECT 1145.040 288.020 1145.300 288.280 ;
        RECT 1235.200 288.020 1235.460 288.280 ;
        RECT 1138.600 17.040 1138.860 17.300 ;
        RECT 1145.040 17.040 1145.300 17.300 ;
      LAYER met2 ;
        RECT 1235.200 300.000 1235.480 304.000 ;
        RECT 1235.260 288.310 1235.400 300.000 ;
        RECT 1145.040 287.990 1145.300 288.310 ;
        RECT 1235.200 287.990 1235.460 288.310 ;
        RECT 1145.100 17.330 1145.240 287.990 ;
        RECT 1138.600 17.010 1138.860 17.330 ;
        RECT 1145.040 17.010 1145.300 17.330 ;
        RECT 1138.660 2.400 1138.800 17.010 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1158.810 286.860 1159.130 286.920 ;
        RECT 1249.890 286.860 1250.210 286.920 ;
        RECT 1158.810 286.720 1250.210 286.860 ;
        RECT 1158.810 286.660 1159.130 286.720 ;
        RECT 1249.890 286.660 1250.210 286.720 ;
        RECT 1156.510 17.580 1156.830 17.640 ;
        RECT 1158.810 17.580 1159.130 17.640 ;
        RECT 1156.510 17.440 1159.130 17.580 ;
        RECT 1156.510 17.380 1156.830 17.440 ;
        RECT 1158.810 17.380 1159.130 17.440 ;
      LAYER via ;
        RECT 1158.840 286.660 1159.100 286.920 ;
        RECT 1249.920 286.660 1250.180 286.920 ;
        RECT 1156.540 17.380 1156.800 17.640 ;
        RECT 1158.840 17.380 1159.100 17.640 ;
      LAYER met2 ;
        RECT 1249.920 300.000 1250.200 304.000 ;
        RECT 1249.980 286.950 1250.120 300.000 ;
        RECT 1158.840 286.630 1159.100 286.950 ;
        RECT 1249.920 286.630 1250.180 286.950 ;
        RECT 1158.900 17.670 1159.040 286.630 ;
        RECT 1156.540 17.350 1156.800 17.670 ;
        RECT 1158.840 17.350 1159.100 17.670 ;
        RECT 1156.600 2.400 1156.740 17.350 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 674.430 25.400 674.750 25.460 ;
        RECT 848.770 25.400 849.090 25.460 ;
        RECT 674.430 25.260 849.090 25.400 ;
        RECT 674.430 25.200 674.750 25.260 ;
        RECT 848.770 25.200 849.090 25.260 ;
      LAYER via ;
        RECT 674.460 25.200 674.720 25.460 ;
        RECT 848.800 25.200 849.060 25.460 ;
      LAYER met2 ;
        RECT 853.400 300.290 853.680 304.000 ;
        RECT 848.860 300.150 853.680 300.290 ;
        RECT 848.860 25.490 849.000 300.150 ;
        RECT 853.400 300.000 853.680 300.150 ;
        RECT 674.460 25.170 674.720 25.490 ;
        RECT 848.800 25.170 849.060 25.490 ;
        RECT 674.520 2.400 674.660 25.170 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1179.510 283.800 1179.830 283.860 ;
        RECT 1264.610 283.800 1264.930 283.860 ;
        RECT 1179.510 283.660 1264.930 283.800 ;
        RECT 1179.510 283.600 1179.830 283.660 ;
        RECT 1264.610 283.600 1264.930 283.660 ;
        RECT 1173.990 16.560 1174.310 16.620 ;
        RECT 1179.510 16.560 1179.830 16.620 ;
        RECT 1173.990 16.420 1179.830 16.560 ;
        RECT 1173.990 16.360 1174.310 16.420 ;
        RECT 1179.510 16.360 1179.830 16.420 ;
      LAYER via ;
        RECT 1179.540 283.600 1179.800 283.860 ;
        RECT 1264.640 283.600 1264.900 283.860 ;
        RECT 1174.020 16.360 1174.280 16.620 ;
        RECT 1179.540 16.360 1179.800 16.620 ;
      LAYER met2 ;
        RECT 1264.640 300.000 1264.920 304.000 ;
        RECT 1264.700 283.890 1264.840 300.000 ;
        RECT 1179.540 283.570 1179.800 283.890 ;
        RECT 1264.640 283.570 1264.900 283.890 ;
        RECT 1179.600 16.650 1179.740 283.570 ;
        RECT 1174.020 16.330 1174.280 16.650 ;
        RECT 1179.540 16.330 1179.800 16.650 ;
        RECT 1174.080 2.400 1174.220 16.330 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1193.310 285.160 1193.630 285.220 ;
        RECT 1279.330 285.160 1279.650 285.220 ;
        RECT 1193.310 285.020 1279.650 285.160 ;
        RECT 1193.310 284.960 1193.630 285.020 ;
        RECT 1279.330 284.960 1279.650 285.020 ;
      LAYER via ;
        RECT 1193.340 284.960 1193.600 285.220 ;
        RECT 1279.360 284.960 1279.620 285.220 ;
      LAYER met2 ;
        RECT 1279.360 300.000 1279.640 304.000 ;
        RECT 1279.420 285.250 1279.560 300.000 ;
        RECT 1193.340 284.930 1193.600 285.250 ;
        RECT 1279.360 284.930 1279.620 285.250 ;
        RECT 1193.400 17.410 1193.540 284.930 ;
        RECT 1192.020 17.270 1193.540 17.410 ;
        RECT 1192.020 2.400 1192.160 17.270 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1214.010 285.500 1214.330 285.560 ;
        RECT 1294.050 285.500 1294.370 285.560 ;
        RECT 1214.010 285.360 1294.370 285.500 ;
        RECT 1214.010 285.300 1214.330 285.360 ;
        RECT 1294.050 285.300 1294.370 285.360 ;
        RECT 1209.870 17.240 1210.190 17.300 ;
        RECT 1214.010 17.240 1214.330 17.300 ;
        RECT 1209.870 17.100 1214.330 17.240 ;
        RECT 1209.870 17.040 1210.190 17.100 ;
        RECT 1214.010 17.040 1214.330 17.100 ;
      LAYER via ;
        RECT 1214.040 285.300 1214.300 285.560 ;
        RECT 1294.080 285.300 1294.340 285.560 ;
        RECT 1209.900 17.040 1210.160 17.300 ;
        RECT 1214.040 17.040 1214.300 17.300 ;
      LAYER met2 ;
        RECT 1294.080 300.000 1294.360 304.000 ;
        RECT 1294.140 285.590 1294.280 300.000 ;
        RECT 1214.040 285.270 1214.300 285.590 ;
        RECT 1294.080 285.270 1294.340 285.590 ;
        RECT 1214.100 17.330 1214.240 285.270 ;
        RECT 1209.900 17.010 1210.160 17.330 ;
        RECT 1214.040 17.010 1214.300 17.330 ;
        RECT 1209.960 2.400 1210.100 17.010 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 289.580 1228.130 289.640 ;
        RECT 1308.770 289.580 1309.090 289.640 ;
        RECT 1227.810 289.440 1309.090 289.580 ;
        RECT 1227.810 289.380 1228.130 289.440 ;
        RECT 1308.770 289.380 1309.090 289.440 ;
      LAYER via ;
        RECT 1227.840 289.380 1228.100 289.640 ;
        RECT 1308.800 289.380 1309.060 289.640 ;
      LAYER met2 ;
        RECT 1308.800 300.000 1309.080 304.000 ;
        RECT 1308.860 289.670 1309.000 300.000 ;
        RECT 1227.840 289.350 1228.100 289.670 ;
        RECT 1308.800 289.350 1309.060 289.670 ;
        RECT 1227.900 2.400 1228.040 289.350 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1248.510 284.820 1248.830 284.880 ;
        RECT 1323.490 284.820 1323.810 284.880 ;
        RECT 1248.510 284.680 1323.810 284.820 ;
        RECT 1248.510 284.620 1248.830 284.680 ;
        RECT 1323.490 284.620 1323.810 284.680 ;
        RECT 1245.750 17.580 1246.070 17.640 ;
        RECT 1248.510 17.580 1248.830 17.640 ;
        RECT 1245.750 17.440 1248.830 17.580 ;
        RECT 1245.750 17.380 1246.070 17.440 ;
        RECT 1248.510 17.380 1248.830 17.440 ;
      LAYER via ;
        RECT 1248.540 284.620 1248.800 284.880 ;
        RECT 1323.520 284.620 1323.780 284.880 ;
        RECT 1245.780 17.380 1246.040 17.640 ;
        RECT 1248.540 17.380 1248.800 17.640 ;
      LAYER met2 ;
        RECT 1323.520 300.000 1323.800 304.000 ;
        RECT 1323.580 284.910 1323.720 300.000 ;
        RECT 1248.540 284.590 1248.800 284.910 ;
        RECT 1323.520 284.590 1323.780 284.910 ;
        RECT 1248.600 17.670 1248.740 284.590 ;
        RECT 1245.780 17.350 1246.040 17.670 ;
        RECT 1248.540 17.350 1248.800 17.670 ;
        RECT 1245.840 2.400 1245.980 17.350 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1269.210 284.140 1269.530 284.200 ;
        RECT 1336.830 284.140 1337.150 284.200 ;
        RECT 1269.210 284.000 1337.150 284.140 ;
        RECT 1269.210 283.940 1269.530 284.000 ;
        RECT 1336.830 283.940 1337.150 284.000 ;
        RECT 1263.230 17.920 1263.550 17.980 ;
        RECT 1269.210 17.920 1269.530 17.980 ;
        RECT 1263.230 17.780 1269.530 17.920 ;
        RECT 1263.230 17.720 1263.550 17.780 ;
        RECT 1269.210 17.720 1269.530 17.780 ;
      LAYER via ;
        RECT 1269.240 283.940 1269.500 284.200 ;
        RECT 1336.860 283.940 1337.120 284.200 ;
        RECT 1263.260 17.720 1263.520 17.980 ;
        RECT 1269.240 17.720 1269.500 17.980 ;
      LAYER met2 ;
        RECT 1338.240 300.290 1338.520 304.000 ;
        RECT 1336.920 300.150 1338.520 300.290 ;
        RECT 1336.920 284.230 1337.060 300.150 ;
        RECT 1338.240 300.000 1338.520 300.150 ;
        RECT 1269.240 283.910 1269.500 284.230 ;
        RECT 1336.860 283.910 1337.120 284.230 ;
        RECT 1269.300 18.010 1269.440 283.910 ;
        RECT 1263.260 17.690 1263.520 18.010 ;
        RECT 1269.240 17.690 1269.500 18.010 ;
        RECT 1263.320 2.400 1263.460 17.690 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.010 287.880 1283.330 287.940 ;
        RECT 1352.930 287.880 1353.250 287.940 ;
        RECT 1283.010 287.740 1353.250 287.880 ;
        RECT 1283.010 287.680 1283.330 287.740 ;
        RECT 1352.930 287.680 1353.250 287.740 ;
      LAYER via ;
        RECT 1283.040 287.680 1283.300 287.940 ;
        RECT 1352.960 287.680 1353.220 287.940 ;
      LAYER met2 ;
        RECT 1352.960 300.000 1353.240 304.000 ;
        RECT 1353.020 287.970 1353.160 300.000 ;
        RECT 1283.040 287.650 1283.300 287.970 ;
        RECT 1352.960 287.650 1353.220 287.970 ;
        RECT 1283.100 17.410 1283.240 287.650 ;
        RECT 1281.260 17.270 1283.240 17.410 ;
        RECT 1281.260 2.400 1281.400 17.270 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1303.710 287.540 1304.030 287.600 ;
        RECT 1367.650 287.540 1367.970 287.600 ;
        RECT 1303.710 287.400 1367.970 287.540 ;
        RECT 1303.710 287.340 1304.030 287.400 ;
        RECT 1367.650 287.340 1367.970 287.400 ;
        RECT 1299.110 17.580 1299.430 17.640 ;
        RECT 1303.710 17.580 1304.030 17.640 ;
        RECT 1299.110 17.440 1304.030 17.580 ;
        RECT 1299.110 17.380 1299.430 17.440 ;
        RECT 1303.710 17.380 1304.030 17.440 ;
      LAYER via ;
        RECT 1303.740 287.340 1304.000 287.600 ;
        RECT 1367.680 287.340 1367.940 287.600 ;
        RECT 1299.140 17.380 1299.400 17.640 ;
        RECT 1303.740 17.380 1304.000 17.640 ;
      LAYER met2 ;
        RECT 1367.680 300.000 1367.960 304.000 ;
        RECT 1367.740 287.630 1367.880 300.000 ;
        RECT 1303.740 287.310 1304.000 287.630 ;
        RECT 1367.680 287.310 1367.940 287.630 ;
        RECT 1303.800 17.670 1303.940 287.310 ;
        RECT 1299.140 17.350 1299.400 17.670 ;
        RECT 1303.740 17.350 1304.000 17.670 ;
        RECT 1299.200 2.400 1299.340 17.350 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.050 286.180 1317.370 286.240 ;
        RECT 1381.910 286.180 1382.230 286.240 ;
        RECT 1317.050 286.040 1382.230 286.180 ;
        RECT 1317.050 285.980 1317.370 286.040 ;
        RECT 1381.910 285.980 1382.230 286.040 ;
      LAYER via ;
        RECT 1317.080 285.980 1317.340 286.240 ;
        RECT 1381.940 285.980 1382.200 286.240 ;
      LAYER met2 ;
        RECT 1381.940 300.000 1382.220 304.000 ;
        RECT 1382.000 286.270 1382.140 300.000 ;
        RECT 1317.080 285.950 1317.340 286.270 ;
        RECT 1381.940 285.950 1382.200 286.270 ;
        RECT 1317.140 2.400 1317.280 285.950 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 288.220 1338.530 288.280 ;
        RECT 1396.630 288.220 1396.950 288.280 ;
        RECT 1338.210 288.080 1396.950 288.220 ;
        RECT 1338.210 288.020 1338.530 288.080 ;
        RECT 1396.630 288.020 1396.950 288.080 ;
        RECT 1334.990 17.240 1335.310 17.300 ;
        RECT 1338.210 17.240 1338.530 17.300 ;
        RECT 1334.990 17.100 1338.530 17.240 ;
        RECT 1334.990 17.040 1335.310 17.100 ;
        RECT 1338.210 17.040 1338.530 17.100 ;
      LAYER via ;
        RECT 1338.240 288.020 1338.500 288.280 ;
        RECT 1396.660 288.020 1396.920 288.280 ;
        RECT 1335.020 17.040 1335.280 17.300 ;
        RECT 1338.240 17.040 1338.500 17.300 ;
      LAYER met2 ;
        RECT 1396.660 300.000 1396.940 304.000 ;
        RECT 1396.720 288.310 1396.860 300.000 ;
        RECT 1338.240 287.990 1338.500 288.310 ;
        RECT 1396.660 287.990 1396.920 288.310 ;
        RECT 1338.300 17.330 1338.440 287.990 ;
        RECT 1335.020 17.010 1335.280 17.330 ;
        RECT 1338.240 17.010 1338.500 17.330 ;
        RECT 1335.080 2.400 1335.220 17.010 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 695.590 288.560 695.910 288.620 ;
        RECT 695.590 288.420 736.760 288.560 ;
        RECT 695.590 288.360 695.910 288.420 ;
        RECT 736.620 288.220 736.760 288.420 ;
        RECT 868.090 288.220 868.410 288.280 ;
        RECT 736.620 288.080 868.410 288.220 ;
        RECT 868.090 288.020 868.410 288.080 ;
        RECT 692.370 20.640 692.690 20.700 ;
        RECT 696.510 20.640 696.830 20.700 ;
        RECT 692.370 20.500 696.830 20.640 ;
        RECT 692.370 20.440 692.690 20.500 ;
        RECT 696.510 20.440 696.830 20.500 ;
      LAYER via ;
        RECT 695.620 288.360 695.880 288.620 ;
        RECT 868.120 288.020 868.380 288.280 ;
        RECT 692.400 20.440 692.660 20.700 ;
        RECT 696.540 20.440 696.800 20.700 ;
      LAYER met2 ;
        RECT 868.120 300.000 868.400 304.000 ;
        RECT 695.620 288.330 695.880 288.650 ;
        RECT 695.680 271.730 695.820 288.330 ;
        RECT 868.180 288.310 868.320 300.000 ;
        RECT 868.120 287.990 868.380 288.310 ;
        RECT 695.680 271.590 696.740 271.730 ;
        RECT 696.600 20.730 696.740 271.590 ;
        RECT 692.400 20.410 692.660 20.730 ;
        RECT 696.540 20.410 696.800 20.730 ;
        RECT 692.460 2.400 692.600 20.410 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1358.450 288.560 1358.770 288.620 ;
        RECT 1411.350 288.560 1411.670 288.620 ;
        RECT 1358.450 288.420 1411.670 288.560 ;
        RECT 1358.450 288.360 1358.770 288.420 ;
        RECT 1411.350 288.360 1411.670 288.420 ;
        RECT 1352.470 17.920 1352.790 17.980 ;
        RECT 1358.450 17.920 1358.770 17.980 ;
        RECT 1352.470 17.780 1358.770 17.920 ;
        RECT 1352.470 17.720 1352.790 17.780 ;
        RECT 1358.450 17.720 1358.770 17.780 ;
      LAYER via ;
        RECT 1358.480 288.360 1358.740 288.620 ;
        RECT 1411.380 288.360 1411.640 288.620 ;
        RECT 1352.500 17.720 1352.760 17.980 ;
        RECT 1358.480 17.720 1358.740 17.980 ;
      LAYER met2 ;
        RECT 1411.380 300.000 1411.660 304.000 ;
        RECT 1411.440 288.650 1411.580 300.000 ;
        RECT 1358.480 288.330 1358.740 288.650 ;
        RECT 1411.380 288.330 1411.640 288.650 ;
        RECT 1358.540 18.010 1358.680 288.330 ;
        RECT 1352.500 17.690 1352.760 18.010 ;
        RECT 1358.480 17.690 1358.740 18.010 ;
        RECT 1352.560 2.400 1352.700 17.690 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1372.710 289.240 1373.030 289.300 ;
        RECT 1426.070 289.240 1426.390 289.300 ;
        RECT 1372.710 289.100 1426.390 289.240 ;
        RECT 1372.710 289.040 1373.030 289.100 ;
        RECT 1426.070 289.040 1426.390 289.100 ;
        RECT 1370.410 17.580 1370.730 17.640 ;
        RECT 1372.710 17.580 1373.030 17.640 ;
        RECT 1370.410 17.440 1373.030 17.580 ;
        RECT 1370.410 17.380 1370.730 17.440 ;
        RECT 1372.710 17.380 1373.030 17.440 ;
      LAYER via ;
        RECT 1372.740 289.040 1373.000 289.300 ;
        RECT 1426.100 289.040 1426.360 289.300 ;
        RECT 1370.440 17.380 1370.700 17.640 ;
        RECT 1372.740 17.380 1373.000 17.640 ;
      LAYER met2 ;
        RECT 1426.100 300.000 1426.380 304.000 ;
        RECT 1426.160 289.330 1426.300 300.000 ;
        RECT 1372.740 289.010 1373.000 289.330 ;
        RECT 1426.100 289.010 1426.360 289.330 ;
        RECT 1372.800 17.670 1372.940 289.010 ;
        RECT 1370.440 17.350 1370.700 17.670 ;
        RECT 1372.740 17.350 1373.000 17.670 ;
        RECT 1370.500 2.400 1370.640 17.350 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1393.410 286.520 1393.730 286.580 ;
        RECT 1440.790 286.520 1441.110 286.580 ;
        RECT 1393.410 286.380 1441.110 286.520 ;
        RECT 1393.410 286.320 1393.730 286.380 ;
        RECT 1440.790 286.320 1441.110 286.380 ;
        RECT 1388.350 17.580 1388.670 17.640 ;
        RECT 1393.410 17.580 1393.730 17.640 ;
        RECT 1388.350 17.440 1393.730 17.580 ;
        RECT 1388.350 17.380 1388.670 17.440 ;
        RECT 1393.410 17.380 1393.730 17.440 ;
      LAYER via ;
        RECT 1393.440 286.320 1393.700 286.580 ;
        RECT 1440.820 286.320 1441.080 286.580 ;
        RECT 1388.380 17.380 1388.640 17.640 ;
        RECT 1393.440 17.380 1393.700 17.640 ;
      LAYER met2 ;
        RECT 1440.820 300.000 1441.100 304.000 ;
        RECT 1440.880 286.610 1441.020 300.000 ;
        RECT 1393.440 286.290 1393.700 286.610 ;
        RECT 1440.820 286.290 1441.080 286.610 ;
        RECT 1393.500 17.670 1393.640 286.290 ;
        RECT 1388.380 17.350 1388.640 17.670 ;
        RECT 1393.440 17.350 1393.700 17.670 ;
        RECT 1388.440 2.400 1388.580 17.350 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1407.210 288.220 1407.530 288.280 ;
        RECT 1455.510 288.220 1455.830 288.280 ;
        RECT 1407.210 288.080 1455.830 288.220 ;
        RECT 1407.210 288.020 1407.530 288.080 ;
        RECT 1455.510 288.020 1455.830 288.080 ;
      LAYER via ;
        RECT 1407.240 288.020 1407.500 288.280 ;
        RECT 1455.540 288.020 1455.800 288.280 ;
      LAYER met2 ;
        RECT 1455.540 300.000 1455.820 304.000 ;
        RECT 1455.600 288.310 1455.740 300.000 ;
        RECT 1407.240 287.990 1407.500 288.310 ;
        RECT 1455.540 287.990 1455.800 288.310 ;
        RECT 1407.300 17.580 1407.440 287.990 ;
        RECT 1406.380 17.440 1407.440 17.580 ;
        RECT 1406.380 2.400 1406.520 17.440 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1427.910 286.860 1428.230 286.920 ;
        RECT 1470.230 286.860 1470.550 286.920 ;
        RECT 1427.910 286.720 1470.550 286.860 ;
        RECT 1427.910 286.660 1428.230 286.720 ;
        RECT 1470.230 286.660 1470.550 286.720 ;
        RECT 1423.770 17.580 1424.090 17.640 ;
        RECT 1427.910 17.580 1428.230 17.640 ;
        RECT 1423.770 17.440 1428.230 17.580 ;
        RECT 1423.770 17.380 1424.090 17.440 ;
        RECT 1427.910 17.380 1428.230 17.440 ;
      LAYER via ;
        RECT 1427.940 286.660 1428.200 286.920 ;
        RECT 1470.260 286.660 1470.520 286.920 ;
        RECT 1423.800 17.380 1424.060 17.640 ;
        RECT 1427.940 17.380 1428.200 17.640 ;
      LAYER met2 ;
        RECT 1470.260 300.000 1470.540 304.000 ;
        RECT 1470.320 286.950 1470.460 300.000 ;
        RECT 1427.940 286.630 1428.200 286.950 ;
        RECT 1470.260 286.630 1470.520 286.950 ;
        RECT 1428.000 17.670 1428.140 286.630 ;
        RECT 1423.800 17.350 1424.060 17.670 ;
        RECT 1427.940 17.350 1428.200 17.670 ;
        RECT 1423.860 2.400 1424.000 17.350 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1441.250 286.520 1441.570 286.580 ;
        RECT 1484.950 286.520 1485.270 286.580 ;
        RECT 1441.250 286.380 1485.270 286.520 ;
        RECT 1441.250 286.320 1441.570 286.380 ;
        RECT 1484.950 286.320 1485.270 286.380 ;
      LAYER via ;
        RECT 1441.280 286.320 1441.540 286.580 ;
        RECT 1484.980 286.320 1485.240 286.580 ;
      LAYER met2 ;
        RECT 1484.980 300.000 1485.260 304.000 ;
        RECT 1485.040 286.610 1485.180 300.000 ;
        RECT 1441.280 286.290 1441.540 286.610 ;
        RECT 1484.980 286.290 1485.240 286.610 ;
        RECT 1441.340 17.410 1441.480 286.290 ;
        RECT 1441.340 17.270 1441.940 17.410 ;
        RECT 1441.800 2.400 1441.940 17.270 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1462.410 287.200 1462.730 287.260 ;
        RECT 1499.670 287.200 1499.990 287.260 ;
        RECT 1462.410 287.060 1499.990 287.200 ;
        RECT 1462.410 287.000 1462.730 287.060 ;
        RECT 1499.670 287.000 1499.990 287.060 ;
        RECT 1459.650 17.580 1459.970 17.640 ;
        RECT 1462.410 17.580 1462.730 17.640 ;
        RECT 1459.650 17.440 1462.730 17.580 ;
        RECT 1459.650 17.380 1459.970 17.440 ;
        RECT 1462.410 17.380 1462.730 17.440 ;
      LAYER via ;
        RECT 1462.440 287.000 1462.700 287.260 ;
        RECT 1499.700 287.000 1499.960 287.260 ;
        RECT 1459.680 17.380 1459.940 17.640 ;
        RECT 1462.440 17.380 1462.700 17.640 ;
      LAYER met2 ;
        RECT 1499.700 300.000 1499.980 304.000 ;
        RECT 1499.760 287.290 1499.900 300.000 ;
        RECT 1462.440 286.970 1462.700 287.290 ;
        RECT 1499.700 286.970 1499.960 287.290 ;
        RECT 1462.500 17.670 1462.640 286.970 ;
        RECT 1459.680 17.350 1459.940 17.670 ;
        RECT 1462.440 17.350 1462.700 17.670 ;
        RECT 1459.740 2.400 1459.880 17.350 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1483.110 288.560 1483.430 288.620 ;
        RECT 1514.390 288.560 1514.710 288.620 ;
        RECT 1483.110 288.420 1514.710 288.560 ;
        RECT 1483.110 288.360 1483.430 288.420 ;
        RECT 1514.390 288.360 1514.710 288.420 ;
        RECT 1477.590 17.580 1477.910 17.640 ;
        RECT 1483.110 17.580 1483.430 17.640 ;
        RECT 1477.590 17.440 1483.430 17.580 ;
        RECT 1477.590 17.380 1477.910 17.440 ;
        RECT 1483.110 17.380 1483.430 17.440 ;
      LAYER via ;
        RECT 1483.140 288.360 1483.400 288.620 ;
        RECT 1514.420 288.360 1514.680 288.620 ;
        RECT 1477.620 17.380 1477.880 17.640 ;
        RECT 1483.140 17.380 1483.400 17.640 ;
      LAYER met2 ;
        RECT 1514.420 300.000 1514.700 304.000 ;
        RECT 1514.480 288.650 1514.620 300.000 ;
        RECT 1483.140 288.330 1483.400 288.650 ;
        RECT 1514.420 288.330 1514.680 288.650 ;
        RECT 1483.200 17.670 1483.340 288.330 ;
        RECT 1477.620 17.350 1477.880 17.670 ;
        RECT 1483.140 17.350 1483.400 17.670 ;
        RECT 1477.680 2.400 1477.820 17.350 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1496.910 287.540 1497.230 287.600 ;
        RECT 1529.110 287.540 1529.430 287.600 ;
        RECT 1496.910 287.400 1529.430 287.540 ;
        RECT 1496.910 287.340 1497.230 287.400 ;
        RECT 1529.110 287.340 1529.430 287.400 ;
      LAYER via ;
        RECT 1496.940 287.340 1497.200 287.600 ;
        RECT 1529.140 287.340 1529.400 287.600 ;
      LAYER met2 ;
        RECT 1529.140 300.000 1529.420 304.000 ;
        RECT 1529.200 287.630 1529.340 300.000 ;
        RECT 1496.940 287.310 1497.200 287.630 ;
        RECT 1529.140 287.310 1529.400 287.630 ;
        RECT 1497.000 17.410 1497.140 287.310 ;
        RECT 1495.620 17.270 1497.140 17.410 ;
        RECT 1495.620 2.400 1495.760 17.270 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1517.610 283.460 1517.930 283.520 ;
        RECT 1543.830 283.460 1544.150 283.520 ;
        RECT 1517.610 283.320 1544.150 283.460 ;
        RECT 1517.610 283.260 1517.930 283.320 ;
        RECT 1543.830 283.260 1544.150 283.320 ;
        RECT 1513.010 17.580 1513.330 17.640 ;
        RECT 1517.610 17.580 1517.930 17.640 ;
        RECT 1513.010 17.440 1517.930 17.580 ;
        RECT 1513.010 17.380 1513.330 17.440 ;
        RECT 1517.610 17.380 1517.930 17.440 ;
      LAYER via ;
        RECT 1517.640 283.260 1517.900 283.520 ;
        RECT 1543.860 283.260 1544.120 283.520 ;
        RECT 1513.040 17.380 1513.300 17.640 ;
        RECT 1517.640 17.380 1517.900 17.640 ;
      LAYER met2 ;
        RECT 1543.860 300.000 1544.140 304.000 ;
        RECT 1543.920 283.550 1544.060 300.000 ;
        RECT 1517.640 283.230 1517.900 283.550 ;
        RECT 1543.860 283.230 1544.120 283.550 ;
        RECT 1517.700 17.670 1517.840 283.230 ;
        RECT 1513.040 17.350 1513.300 17.670 ;
        RECT 1517.640 17.350 1517.900 17.670 ;
        RECT 1513.100 2.400 1513.240 17.350 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 758.685 285.685 758.855 287.895 ;
      LAYER mcon ;
        RECT 758.685 287.725 758.855 287.895 ;
      LAYER met1 ;
        RECT 758.625 287.880 758.915 287.925 ;
        RECT 882.350 287.880 882.670 287.940 ;
        RECT 758.625 287.740 882.670 287.880 ;
        RECT 758.625 287.695 758.915 287.740 ;
        RECT 882.350 287.680 882.670 287.740 ;
        RECT 710.310 285.840 710.630 285.900 ;
        RECT 758.625 285.840 758.915 285.885 ;
        RECT 710.310 285.700 758.915 285.840 ;
        RECT 710.310 285.640 710.630 285.700 ;
        RECT 758.625 285.655 758.915 285.700 ;
      LAYER via ;
        RECT 882.380 287.680 882.640 287.940 ;
        RECT 710.340 285.640 710.600 285.900 ;
      LAYER met2 ;
        RECT 882.380 300.000 882.660 304.000 ;
        RECT 882.440 287.970 882.580 300.000 ;
        RECT 882.380 287.650 882.640 287.970 ;
        RECT 710.340 285.610 710.600 285.930 ;
        RECT 710.400 2.400 710.540 285.610 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1531.410 287.540 1531.730 287.600 ;
        RECT 1558.550 287.540 1558.870 287.600 ;
        RECT 1531.410 287.400 1558.870 287.540 ;
        RECT 1531.410 287.340 1531.730 287.400 ;
        RECT 1558.550 287.340 1558.870 287.400 ;
      LAYER via ;
        RECT 1531.440 287.340 1531.700 287.600 ;
        RECT 1558.580 287.340 1558.840 287.600 ;
      LAYER met2 ;
        RECT 1558.580 300.000 1558.860 304.000 ;
        RECT 1558.640 287.630 1558.780 300.000 ;
        RECT 1531.440 287.310 1531.700 287.630 ;
        RECT 1558.580 287.310 1558.840 287.630 ;
        RECT 1531.500 17.410 1531.640 287.310 ;
        RECT 1531.040 17.270 1531.640 17.410 ;
        RECT 1531.040 2.400 1531.180 17.270 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1552.110 288.560 1552.430 288.620 ;
        RECT 1573.270 288.560 1573.590 288.620 ;
        RECT 1552.110 288.420 1573.590 288.560 ;
        RECT 1552.110 288.360 1552.430 288.420 ;
        RECT 1573.270 288.360 1573.590 288.420 ;
        RECT 1548.890 17.580 1549.210 17.640 ;
        RECT 1552.110 17.580 1552.430 17.640 ;
        RECT 1548.890 17.440 1552.430 17.580 ;
        RECT 1548.890 17.380 1549.210 17.440 ;
        RECT 1552.110 17.380 1552.430 17.440 ;
      LAYER via ;
        RECT 1552.140 288.360 1552.400 288.620 ;
        RECT 1573.300 288.360 1573.560 288.620 ;
        RECT 1548.920 17.380 1549.180 17.640 ;
        RECT 1552.140 17.380 1552.400 17.640 ;
      LAYER met2 ;
        RECT 1573.300 300.000 1573.580 304.000 ;
        RECT 1573.360 288.650 1573.500 300.000 ;
        RECT 1552.140 288.330 1552.400 288.650 ;
        RECT 1573.300 288.330 1573.560 288.650 ;
        RECT 1552.200 17.670 1552.340 288.330 ;
        RECT 1548.920 17.350 1549.180 17.670 ;
        RECT 1552.140 17.350 1552.400 17.670 ;
        RECT 1548.980 2.400 1549.120 17.350 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1583.390 288.220 1583.710 288.280 ;
        RECT 1587.990 288.220 1588.310 288.280 ;
        RECT 1583.390 288.080 1588.310 288.220 ;
        RECT 1583.390 288.020 1583.710 288.080 ;
        RECT 1587.990 288.020 1588.310 288.080 ;
        RECT 1566.830 19.960 1567.150 20.020 ;
        RECT 1583.390 19.960 1583.710 20.020 ;
        RECT 1566.830 19.820 1583.710 19.960 ;
        RECT 1566.830 19.760 1567.150 19.820 ;
        RECT 1583.390 19.760 1583.710 19.820 ;
      LAYER via ;
        RECT 1583.420 288.020 1583.680 288.280 ;
        RECT 1588.020 288.020 1588.280 288.280 ;
        RECT 1566.860 19.760 1567.120 20.020 ;
        RECT 1583.420 19.760 1583.680 20.020 ;
      LAYER met2 ;
        RECT 1588.020 300.000 1588.300 304.000 ;
        RECT 1588.080 288.310 1588.220 300.000 ;
        RECT 1583.420 287.990 1583.680 288.310 ;
        RECT 1588.020 287.990 1588.280 288.310 ;
        RECT 1583.480 20.050 1583.620 287.990 ;
        RECT 1566.860 19.730 1567.120 20.050 ;
        RECT 1583.420 19.730 1583.680 20.050 ;
        RECT 1566.920 2.400 1567.060 19.730 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1586.610 287.880 1586.930 287.940 ;
        RECT 1602.710 287.880 1603.030 287.940 ;
        RECT 1586.610 287.740 1603.030 287.880 ;
        RECT 1586.610 287.680 1586.930 287.740 ;
        RECT 1602.710 287.680 1603.030 287.740 ;
        RECT 1584.770 2.960 1585.090 3.020 ;
        RECT 1586.610 2.960 1586.930 3.020 ;
        RECT 1584.770 2.820 1586.930 2.960 ;
        RECT 1584.770 2.760 1585.090 2.820 ;
        RECT 1586.610 2.760 1586.930 2.820 ;
      LAYER via ;
        RECT 1586.640 287.680 1586.900 287.940 ;
        RECT 1602.740 287.680 1603.000 287.940 ;
        RECT 1584.800 2.760 1585.060 3.020 ;
        RECT 1586.640 2.760 1586.900 3.020 ;
      LAYER met2 ;
        RECT 1602.740 300.000 1603.020 304.000 ;
        RECT 1602.800 287.970 1602.940 300.000 ;
        RECT 1586.640 287.650 1586.900 287.970 ;
        RECT 1602.740 287.650 1603.000 287.970 ;
        RECT 1586.700 3.050 1586.840 287.650 ;
        RECT 1584.800 2.730 1585.060 3.050 ;
        RECT 1586.640 2.730 1586.900 3.050 ;
        RECT 1584.860 2.400 1585.000 2.730 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1607.310 288.560 1607.630 288.620 ;
        RECT 1617.430 288.560 1617.750 288.620 ;
        RECT 1607.310 288.420 1617.750 288.560 ;
        RECT 1607.310 288.360 1607.630 288.420 ;
        RECT 1617.430 288.360 1617.750 288.420 ;
        RECT 1602.250 17.580 1602.570 17.640 ;
        RECT 1607.310 17.580 1607.630 17.640 ;
        RECT 1602.250 17.440 1607.630 17.580 ;
        RECT 1602.250 17.380 1602.570 17.440 ;
        RECT 1607.310 17.380 1607.630 17.440 ;
      LAYER via ;
        RECT 1607.340 288.360 1607.600 288.620 ;
        RECT 1617.460 288.360 1617.720 288.620 ;
        RECT 1602.280 17.380 1602.540 17.640 ;
        RECT 1607.340 17.380 1607.600 17.640 ;
      LAYER met2 ;
        RECT 1617.460 300.000 1617.740 304.000 ;
        RECT 1617.520 288.650 1617.660 300.000 ;
        RECT 1607.340 288.330 1607.600 288.650 ;
        RECT 1617.460 288.330 1617.720 288.650 ;
        RECT 1607.400 17.670 1607.540 288.330 ;
        RECT 1602.280 17.350 1602.540 17.670 ;
        RECT 1607.340 17.350 1607.600 17.670 ;
        RECT 1602.340 2.400 1602.480 17.350 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1621.110 283.460 1621.430 283.520 ;
        RECT 1631.690 283.460 1632.010 283.520 ;
        RECT 1621.110 283.320 1632.010 283.460 ;
        RECT 1621.110 283.260 1621.430 283.320 ;
        RECT 1631.690 283.260 1632.010 283.320 ;
      LAYER via ;
        RECT 1621.140 283.260 1621.400 283.520 ;
        RECT 1631.720 283.260 1631.980 283.520 ;
      LAYER met2 ;
        RECT 1631.720 300.000 1632.000 304.000 ;
        RECT 1631.780 283.550 1631.920 300.000 ;
        RECT 1621.140 283.230 1621.400 283.550 ;
        RECT 1631.720 283.230 1631.980 283.550 ;
        RECT 1621.200 17.410 1621.340 283.230 ;
        RECT 1620.280 17.270 1621.340 17.410 ;
        RECT 1620.280 2.400 1620.420 17.270 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1641.810 288.220 1642.130 288.280 ;
        RECT 1646.410 288.220 1646.730 288.280 ;
        RECT 1641.810 288.080 1646.730 288.220 ;
        RECT 1641.810 288.020 1642.130 288.080 ;
        RECT 1646.410 288.020 1646.730 288.080 ;
        RECT 1638.130 17.580 1638.450 17.640 ;
        RECT 1641.810 17.580 1642.130 17.640 ;
        RECT 1638.130 17.440 1642.130 17.580 ;
        RECT 1638.130 17.380 1638.450 17.440 ;
        RECT 1641.810 17.380 1642.130 17.440 ;
      LAYER via ;
        RECT 1641.840 288.020 1642.100 288.280 ;
        RECT 1646.440 288.020 1646.700 288.280 ;
        RECT 1638.160 17.380 1638.420 17.640 ;
        RECT 1641.840 17.380 1642.100 17.640 ;
      LAYER met2 ;
        RECT 1646.440 300.000 1646.720 304.000 ;
        RECT 1646.500 288.310 1646.640 300.000 ;
        RECT 1641.840 287.990 1642.100 288.310 ;
        RECT 1646.440 287.990 1646.700 288.310 ;
        RECT 1641.900 17.670 1642.040 287.990 ;
        RECT 1638.160 17.350 1638.420 17.670 ;
        RECT 1641.840 17.350 1642.100 17.670 ;
        RECT 1638.220 2.400 1638.360 17.350 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1661.160 300.290 1661.440 304.000 ;
        RECT 1657.080 300.150 1661.440 300.290 ;
        RECT 1657.080 12.650 1657.220 300.150 ;
        RECT 1661.160 300.000 1661.440 300.150 ;
        RECT 1656.160 12.510 1657.220 12.650 ;
        RECT 1656.160 2.400 1656.300 12.510 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1670.865 241.485 1671.035 278.035 ;
        RECT 1669.945 41.565 1670.115 89.675 ;
      LAYER mcon ;
        RECT 1670.865 277.865 1671.035 278.035 ;
        RECT 1669.945 89.505 1670.115 89.675 ;
      LAYER met1 ;
        RECT 1670.805 278.020 1671.095 278.065 ;
        RECT 1671.710 278.020 1672.030 278.080 ;
        RECT 1670.805 277.880 1672.030 278.020 ;
        RECT 1670.805 277.835 1671.095 277.880 ;
        RECT 1671.710 277.820 1672.030 277.880 ;
        RECT 1670.790 241.640 1671.110 241.700 ;
        RECT 1670.595 241.500 1671.110 241.640 ;
        RECT 1670.790 241.440 1671.110 241.500 ;
        RECT 1669.870 158.820 1670.190 159.080 ;
        RECT 1669.960 158.340 1670.100 158.820 ;
        RECT 1670.330 158.340 1670.650 158.400 ;
        RECT 1669.960 158.200 1670.650 158.340 ;
        RECT 1670.330 158.140 1670.650 158.200 ;
        RECT 1669.870 89.660 1670.190 89.720 ;
        RECT 1669.675 89.520 1670.190 89.660 ;
        RECT 1669.870 89.460 1670.190 89.520 ;
        RECT 1669.885 41.720 1670.175 41.765 ;
        RECT 1670.330 41.720 1670.650 41.780 ;
        RECT 1669.885 41.580 1670.650 41.720 ;
        RECT 1669.885 41.535 1670.175 41.580 ;
        RECT 1670.330 41.520 1670.650 41.580 ;
        RECT 1670.330 16.560 1670.650 16.620 ;
        RECT 1673.550 16.560 1673.870 16.620 ;
        RECT 1670.330 16.420 1673.870 16.560 ;
        RECT 1670.330 16.360 1670.650 16.420 ;
        RECT 1673.550 16.360 1673.870 16.420 ;
      LAYER via ;
        RECT 1671.740 277.820 1672.000 278.080 ;
        RECT 1670.820 241.440 1671.080 241.700 ;
        RECT 1669.900 158.820 1670.160 159.080 ;
        RECT 1670.360 158.140 1670.620 158.400 ;
        RECT 1669.900 89.460 1670.160 89.720 ;
        RECT 1670.360 41.520 1670.620 41.780 ;
        RECT 1670.360 16.360 1670.620 16.620 ;
        RECT 1673.580 16.360 1673.840 16.620 ;
      LAYER met2 ;
        RECT 1675.880 300.970 1676.160 304.000 ;
        RECT 1671.800 300.830 1676.160 300.970 ;
        RECT 1671.800 278.110 1671.940 300.830 ;
        RECT 1675.880 300.000 1676.160 300.830 ;
        RECT 1671.740 277.790 1672.000 278.110 ;
        RECT 1670.820 241.410 1671.080 241.730 ;
        RECT 1670.880 207.130 1671.020 241.410 ;
        RECT 1669.960 206.990 1671.020 207.130 ;
        RECT 1669.960 159.110 1670.100 206.990 ;
        RECT 1669.900 158.790 1670.160 159.110 ;
        RECT 1670.360 158.110 1670.620 158.430 ;
        RECT 1670.420 90.965 1670.560 158.110 ;
        RECT 1670.350 90.595 1670.630 90.965 ;
        RECT 1669.890 89.915 1670.170 90.285 ;
        RECT 1669.960 89.750 1670.100 89.915 ;
        RECT 1669.900 89.430 1670.160 89.750 ;
        RECT 1670.360 41.490 1670.620 41.810 ;
        RECT 1670.420 16.650 1670.560 41.490 ;
        RECT 1670.360 16.330 1670.620 16.650 ;
        RECT 1673.580 16.330 1673.840 16.650 ;
        RECT 1673.640 2.400 1673.780 16.330 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
      LAYER via2 ;
        RECT 1670.350 90.640 1670.630 90.920 ;
        RECT 1669.890 89.960 1670.170 90.240 ;
      LAYER met3 ;
        RECT 1670.325 90.930 1670.655 90.945 ;
        RECT 1669.190 90.630 1670.655 90.930 ;
        RECT 1669.190 90.250 1669.490 90.630 ;
        RECT 1670.325 90.615 1670.655 90.630 ;
        RECT 1669.865 90.250 1670.195 90.265 ;
        RECT 1669.190 89.950 1670.195 90.250 ;
        RECT 1669.865 89.935 1670.195 89.950 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1690.645 186.405 1690.815 234.515 ;
        RECT 1690.645 48.365 1690.815 137.955 ;
      LAYER mcon ;
        RECT 1690.645 234.345 1690.815 234.515 ;
        RECT 1690.645 137.785 1690.815 137.955 ;
      LAYER met1 ;
        RECT 1690.570 283.120 1690.890 283.180 ;
        RECT 1691.030 283.120 1691.350 283.180 ;
        RECT 1690.570 282.980 1691.350 283.120 ;
        RECT 1690.570 282.920 1690.890 282.980 ;
        RECT 1691.030 282.920 1691.350 282.980 ;
        RECT 1690.570 234.500 1690.890 234.560 ;
        RECT 1690.375 234.360 1690.890 234.500 ;
        RECT 1690.570 234.300 1690.890 234.360 ;
        RECT 1690.570 186.560 1690.890 186.620 ;
        RECT 1690.375 186.420 1690.890 186.560 ;
        RECT 1690.570 186.360 1690.890 186.420 ;
        RECT 1690.570 137.940 1690.890 138.000 ;
        RECT 1690.375 137.800 1690.890 137.940 ;
        RECT 1690.570 137.740 1690.890 137.800 ;
        RECT 1690.585 48.520 1690.875 48.565 ;
        RECT 1691.490 48.520 1691.810 48.580 ;
        RECT 1690.585 48.380 1691.810 48.520 ;
        RECT 1690.585 48.335 1690.875 48.380 ;
        RECT 1691.490 48.320 1691.810 48.380 ;
      LAYER via ;
        RECT 1690.600 282.920 1690.860 283.180 ;
        RECT 1691.060 282.920 1691.320 283.180 ;
        RECT 1690.600 234.300 1690.860 234.560 ;
        RECT 1690.600 186.360 1690.860 186.620 ;
        RECT 1690.600 137.740 1690.860 138.000 ;
        RECT 1691.520 48.320 1691.780 48.580 ;
      LAYER met2 ;
        RECT 1690.600 300.290 1690.880 304.000 ;
        RECT 1690.600 300.150 1691.260 300.290 ;
        RECT 1690.600 300.000 1690.880 300.150 ;
        RECT 1691.120 283.210 1691.260 300.150 ;
        RECT 1690.600 282.890 1690.860 283.210 ;
        RECT 1691.060 282.890 1691.320 283.210 ;
        RECT 1690.660 234.590 1690.800 282.890 ;
        RECT 1690.600 234.270 1690.860 234.590 ;
        RECT 1690.600 186.330 1690.860 186.650 ;
        RECT 1690.660 138.030 1690.800 186.330 ;
        RECT 1690.600 137.710 1690.860 138.030 ;
        RECT 1691.520 48.290 1691.780 48.610 ;
        RECT 1691.580 2.400 1691.720 48.290 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 728.250 20.640 728.570 20.700 ;
        RECT 731.010 20.640 731.330 20.700 ;
        RECT 728.250 20.500 731.330 20.640 ;
        RECT 728.250 20.440 728.570 20.500 ;
        RECT 731.010 20.440 731.330 20.500 ;
      LAYER via ;
        RECT 728.280 20.440 728.540 20.700 ;
        RECT 731.040 20.440 731.300 20.700 ;
      LAYER met2 ;
        RECT 897.100 300.000 897.380 304.000 ;
        RECT 897.160 286.125 897.300 300.000 ;
        RECT 731.030 285.755 731.310 286.125 ;
        RECT 897.090 285.755 897.370 286.125 ;
        RECT 731.100 20.730 731.240 285.755 ;
        RECT 728.280 20.410 728.540 20.730 ;
        RECT 731.040 20.410 731.300 20.730 ;
        RECT 728.340 2.400 728.480 20.410 ;
        RECT 728.130 -4.800 728.690 2.400 ;
      LAYER via2 ;
        RECT 731.030 285.800 731.310 286.080 ;
        RECT 897.090 285.800 897.370 286.080 ;
      LAYER met3 ;
        RECT 731.005 286.090 731.335 286.105 ;
        RECT 897.065 286.090 897.395 286.105 ;
        RECT 731.005 285.790 897.395 286.090 ;
        RECT 731.005 285.775 731.335 285.790 ;
        RECT 897.065 285.775 897.395 285.790 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1704.370 17.580 1704.690 17.640 ;
        RECT 1709.430 17.580 1709.750 17.640 ;
        RECT 1704.370 17.440 1709.750 17.580 ;
        RECT 1704.370 17.380 1704.690 17.440 ;
        RECT 1709.430 17.380 1709.750 17.440 ;
      LAYER via ;
        RECT 1704.400 17.380 1704.660 17.640 ;
        RECT 1709.460 17.380 1709.720 17.640 ;
      LAYER met2 ;
        RECT 1705.320 300.290 1705.600 304.000 ;
        RECT 1704.460 300.150 1705.600 300.290 ;
        RECT 1704.460 17.670 1704.600 300.150 ;
        RECT 1705.320 300.000 1705.600 300.150 ;
        RECT 1704.400 17.350 1704.660 17.670 ;
        RECT 1709.460 17.350 1709.720 17.670 ;
        RECT 1709.520 2.400 1709.660 17.350 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1720.010 288.220 1720.330 288.280 ;
        RECT 1724.610 288.220 1724.930 288.280 ;
        RECT 1720.010 288.080 1724.930 288.220 ;
        RECT 1720.010 288.020 1720.330 288.080 ;
        RECT 1724.610 288.020 1724.930 288.080 ;
        RECT 1724.610 20.640 1724.930 20.700 ;
        RECT 1727.370 20.640 1727.690 20.700 ;
        RECT 1724.610 20.500 1727.690 20.640 ;
        RECT 1724.610 20.440 1724.930 20.500 ;
        RECT 1727.370 20.440 1727.690 20.500 ;
      LAYER via ;
        RECT 1720.040 288.020 1720.300 288.280 ;
        RECT 1724.640 288.020 1724.900 288.280 ;
        RECT 1724.640 20.440 1724.900 20.700 ;
        RECT 1727.400 20.440 1727.660 20.700 ;
      LAYER met2 ;
        RECT 1720.040 300.000 1720.320 304.000 ;
        RECT 1720.100 288.310 1720.240 300.000 ;
        RECT 1720.040 287.990 1720.300 288.310 ;
        RECT 1724.640 287.990 1724.900 288.310 ;
        RECT 1724.700 20.730 1724.840 287.990 ;
        RECT 1724.640 20.410 1724.900 20.730 ;
        RECT 1727.400 20.410 1727.660 20.730 ;
        RECT 1727.460 2.400 1727.600 20.410 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1734.730 288.220 1735.050 288.280 ;
        RECT 1739.790 288.220 1740.110 288.280 ;
        RECT 1734.730 288.080 1740.110 288.220 ;
        RECT 1734.730 288.020 1735.050 288.080 ;
        RECT 1739.790 288.020 1740.110 288.080 ;
      LAYER via ;
        RECT 1734.760 288.020 1735.020 288.280 ;
        RECT 1739.820 288.020 1740.080 288.280 ;
      LAYER met2 ;
        RECT 1734.760 300.000 1735.040 304.000 ;
        RECT 1734.820 288.310 1734.960 300.000 ;
        RECT 1734.760 287.990 1735.020 288.310 ;
        RECT 1739.820 287.990 1740.080 288.310 ;
        RECT 1739.880 3.130 1740.020 287.990 ;
        RECT 1739.880 2.990 1745.540 3.130 ;
        RECT 1745.400 2.400 1745.540 2.990 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1749.450 287.880 1749.770 287.940 ;
        RECT 1760.030 287.880 1760.350 287.940 ;
        RECT 1749.450 287.740 1760.350 287.880 ;
        RECT 1749.450 287.680 1749.770 287.740 ;
        RECT 1760.030 287.680 1760.350 287.740 ;
      LAYER via ;
        RECT 1749.480 287.680 1749.740 287.940 ;
        RECT 1760.060 287.680 1760.320 287.940 ;
      LAYER met2 ;
        RECT 1749.480 300.000 1749.760 304.000 ;
        RECT 1749.540 287.970 1749.680 300.000 ;
        RECT 1749.480 287.650 1749.740 287.970 ;
        RECT 1760.060 287.650 1760.320 287.970 ;
        RECT 1760.120 17.410 1760.260 287.650 ;
        RECT 1760.120 17.270 1763.020 17.410 ;
        RECT 1762.880 2.400 1763.020 17.270 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1766.010 20.640 1766.330 20.700 ;
        RECT 1780.730 20.640 1781.050 20.700 ;
        RECT 1766.010 20.500 1781.050 20.640 ;
        RECT 1766.010 20.440 1766.330 20.500 ;
        RECT 1780.730 20.440 1781.050 20.500 ;
      LAYER via ;
        RECT 1766.040 20.440 1766.300 20.700 ;
        RECT 1780.760 20.440 1781.020 20.700 ;
      LAYER met2 ;
        RECT 1764.200 300.290 1764.480 304.000 ;
        RECT 1764.200 300.150 1766.240 300.290 ;
        RECT 1764.200 300.000 1764.480 300.150 ;
        RECT 1766.100 20.730 1766.240 300.150 ;
        RECT 1766.040 20.410 1766.300 20.730 ;
        RECT 1780.760 20.410 1781.020 20.730 ;
        RECT 1780.820 2.400 1780.960 20.410 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1779.810 17.240 1780.130 17.300 ;
        RECT 1798.670 17.240 1798.990 17.300 ;
        RECT 1779.810 17.100 1798.990 17.240 ;
        RECT 1779.810 17.040 1780.130 17.100 ;
        RECT 1798.670 17.040 1798.990 17.100 ;
      LAYER via ;
        RECT 1779.840 17.040 1780.100 17.300 ;
        RECT 1798.700 17.040 1798.960 17.300 ;
      LAYER met2 ;
        RECT 1778.920 300.290 1779.200 304.000 ;
        RECT 1778.920 300.150 1780.040 300.290 ;
        RECT 1778.920 300.000 1779.200 300.150 ;
        RECT 1779.900 17.330 1780.040 300.150 ;
        RECT 1779.840 17.010 1780.100 17.330 ;
        RECT 1798.700 17.010 1798.960 17.330 ;
        RECT 1798.760 2.400 1798.900 17.010 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1793.610 17.920 1793.930 17.980 ;
        RECT 1816.610 17.920 1816.930 17.980 ;
        RECT 1793.610 17.780 1816.930 17.920 ;
        RECT 1793.610 17.720 1793.930 17.780 ;
        RECT 1816.610 17.720 1816.930 17.780 ;
      LAYER via ;
        RECT 1793.640 17.720 1793.900 17.980 ;
        RECT 1816.640 17.720 1816.900 17.980 ;
      LAYER met2 ;
        RECT 1793.640 300.000 1793.920 304.000 ;
        RECT 1793.700 18.010 1793.840 300.000 ;
        RECT 1793.640 17.690 1793.900 18.010 ;
        RECT 1816.640 17.690 1816.900 18.010 ;
        RECT 1816.700 2.400 1816.840 17.690 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1808.330 287.880 1808.650 287.940 ;
        RECT 1813.850 287.880 1814.170 287.940 ;
        RECT 1808.330 287.740 1814.170 287.880 ;
        RECT 1808.330 287.680 1808.650 287.740 ;
        RECT 1813.850 287.680 1814.170 287.740 ;
        RECT 1813.850 20.300 1814.170 20.360 ;
        RECT 1834.550 20.300 1834.870 20.360 ;
        RECT 1813.850 20.160 1834.870 20.300 ;
        RECT 1813.850 20.100 1814.170 20.160 ;
        RECT 1834.550 20.100 1834.870 20.160 ;
      LAYER via ;
        RECT 1808.360 287.680 1808.620 287.940 ;
        RECT 1813.880 287.680 1814.140 287.940 ;
        RECT 1813.880 20.100 1814.140 20.360 ;
        RECT 1834.580 20.100 1834.840 20.360 ;
      LAYER met2 ;
        RECT 1808.360 300.000 1808.640 304.000 ;
        RECT 1808.420 287.970 1808.560 300.000 ;
        RECT 1808.360 287.650 1808.620 287.970 ;
        RECT 1813.880 287.650 1814.140 287.970 ;
        RECT 1813.940 20.390 1814.080 287.650 ;
        RECT 1813.880 20.070 1814.140 20.390 ;
        RECT 1834.580 20.070 1834.840 20.390 ;
        RECT 1834.640 2.400 1834.780 20.070 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1823.050 287.880 1823.370 287.940 ;
        RECT 1849.730 287.880 1850.050 287.940 ;
        RECT 1823.050 287.740 1850.050 287.880 ;
        RECT 1823.050 287.680 1823.370 287.740 ;
        RECT 1849.730 287.680 1850.050 287.740 ;
        RECT 1849.730 2.960 1850.050 3.020 ;
        RECT 1852.030 2.960 1852.350 3.020 ;
        RECT 1849.730 2.820 1852.350 2.960 ;
        RECT 1849.730 2.760 1850.050 2.820 ;
        RECT 1852.030 2.760 1852.350 2.820 ;
      LAYER via ;
        RECT 1823.080 287.680 1823.340 287.940 ;
        RECT 1849.760 287.680 1850.020 287.940 ;
        RECT 1849.760 2.760 1850.020 3.020 ;
        RECT 1852.060 2.760 1852.320 3.020 ;
      LAYER met2 ;
        RECT 1823.080 300.000 1823.360 304.000 ;
        RECT 1823.140 287.970 1823.280 300.000 ;
        RECT 1823.080 287.650 1823.340 287.970 ;
        RECT 1849.760 287.650 1850.020 287.970 ;
        RECT 1849.820 3.050 1849.960 287.650 ;
        RECT 1849.760 2.730 1850.020 3.050 ;
        RECT 1852.060 2.730 1852.320 3.050 ;
        RECT 1852.120 2.400 1852.260 2.730 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1837.770 288.220 1838.090 288.280 ;
        RECT 1841.910 288.220 1842.230 288.280 ;
        RECT 1837.770 288.080 1842.230 288.220 ;
        RECT 1837.770 288.020 1838.090 288.080 ;
        RECT 1841.910 288.020 1842.230 288.080 ;
        RECT 1841.910 15.540 1842.230 15.600 ;
        RECT 1869.970 15.540 1870.290 15.600 ;
        RECT 1841.910 15.400 1870.290 15.540 ;
        RECT 1841.910 15.340 1842.230 15.400 ;
        RECT 1869.970 15.340 1870.290 15.400 ;
      LAYER via ;
        RECT 1837.800 288.020 1838.060 288.280 ;
        RECT 1841.940 288.020 1842.200 288.280 ;
        RECT 1841.940 15.340 1842.200 15.600 ;
        RECT 1870.000 15.340 1870.260 15.600 ;
      LAYER met2 ;
        RECT 1837.800 300.000 1838.080 304.000 ;
        RECT 1837.860 288.310 1838.000 300.000 ;
        RECT 1837.800 287.990 1838.060 288.310 ;
        RECT 1841.940 287.990 1842.200 288.310 ;
        RECT 1842.000 15.630 1842.140 287.990 ;
        RECT 1841.940 15.310 1842.200 15.630 ;
        RECT 1870.000 15.310 1870.260 15.630 ;
        RECT 1870.060 2.400 1870.200 15.310 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 751.710 289.240 752.030 289.300 ;
        RECT 911.790 289.240 912.110 289.300 ;
        RECT 751.710 289.100 912.110 289.240 ;
        RECT 751.710 289.040 752.030 289.100 ;
        RECT 911.790 289.040 912.110 289.100 ;
        RECT 746.190 19.620 746.510 19.680 ;
        RECT 751.710 19.620 752.030 19.680 ;
        RECT 746.190 19.480 752.030 19.620 ;
        RECT 746.190 19.420 746.510 19.480 ;
        RECT 751.710 19.420 752.030 19.480 ;
      LAYER via ;
        RECT 751.740 289.040 752.000 289.300 ;
        RECT 911.820 289.040 912.080 289.300 ;
        RECT 746.220 19.420 746.480 19.680 ;
        RECT 751.740 19.420 752.000 19.680 ;
      LAYER met2 ;
        RECT 911.820 300.000 912.100 304.000 ;
        RECT 911.880 289.330 912.020 300.000 ;
        RECT 751.740 289.010 752.000 289.330 ;
        RECT 911.820 289.010 912.080 289.330 ;
        RECT 751.800 19.710 751.940 289.010 ;
        RECT 746.220 19.390 746.480 19.710 ;
        RECT 751.740 19.390 752.000 19.710 ;
        RECT 746.280 2.400 746.420 19.390 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1855.710 18.940 1856.030 19.000 ;
        RECT 1887.910 18.940 1888.230 19.000 ;
        RECT 1855.710 18.800 1888.230 18.940 ;
        RECT 1855.710 18.740 1856.030 18.800 ;
        RECT 1887.910 18.740 1888.230 18.800 ;
      LAYER via ;
        RECT 1855.740 18.740 1856.000 19.000 ;
        RECT 1887.940 18.740 1888.200 19.000 ;
      LAYER met2 ;
        RECT 1852.520 300.290 1852.800 304.000 ;
        RECT 1852.520 300.150 1855.940 300.290 ;
        RECT 1852.520 300.000 1852.800 300.150 ;
        RECT 1855.800 19.030 1855.940 300.150 ;
        RECT 1855.740 18.710 1856.000 19.030 ;
        RECT 1887.940 18.710 1888.200 19.030 ;
        RECT 1888.000 2.400 1888.140 18.710 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1869.510 17.920 1869.830 17.980 ;
        RECT 1905.850 17.920 1906.170 17.980 ;
        RECT 1869.510 17.780 1906.170 17.920 ;
        RECT 1869.510 17.720 1869.830 17.780 ;
        RECT 1905.850 17.720 1906.170 17.780 ;
      LAYER via ;
        RECT 1869.540 17.720 1869.800 17.980 ;
        RECT 1905.880 17.720 1906.140 17.980 ;
      LAYER met2 ;
        RECT 1867.240 300.290 1867.520 304.000 ;
        RECT 1867.240 300.150 1869.740 300.290 ;
        RECT 1867.240 300.000 1867.520 300.150 ;
        RECT 1869.600 18.010 1869.740 300.150 ;
        RECT 1869.540 17.690 1869.800 18.010 ;
        RECT 1905.880 17.690 1906.140 18.010 ;
        RECT 1905.940 2.400 1906.080 17.690 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1883.310 17.580 1883.630 17.640 ;
        RECT 1923.330 17.580 1923.650 17.640 ;
        RECT 1883.310 17.440 1923.650 17.580 ;
        RECT 1883.310 17.380 1883.630 17.440 ;
        RECT 1923.330 17.380 1923.650 17.440 ;
      LAYER via ;
        RECT 1883.340 17.380 1883.600 17.640 ;
        RECT 1923.360 17.380 1923.620 17.640 ;
      LAYER met2 ;
        RECT 1881.500 300.290 1881.780 304.000 ;
        RECT 1881.500 300.150 1883.540 300.290 ;
        RECT 1881.500 300.000 1881.780 300.150 ;
        RECT 1883.400 17.670 1883.540 300.150 ;
        RECT 1883.340 17.350 1883.600 17.670 ;
        RECT 1923.360 17.350 1923.620 17.670 ;
        RECT 1923.420 2.400 1923.560 17.350 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1896.190 288.220 1896.510 288.280 ;
        RECT 1900.790 288.220 1901.110 288.280 ;
        RECT 1896.190 288.080 1901.110 288.220 ;
        RECT 1896.190 288.020 1896.510 288.080 ;
        RECT 1900.790 288.020 1901.110 288.080 ;
        RECT 1900.790 17.240 1901.110 17.300 ;
        RECT 1941.270 17.240 1941.590 17.300 ;
        RECT 1900.790 17.100 1941.590 17.240 ;
        RECT 1900.790 17.040 1901.110 17.100 ;
        RECT 1941.270 17.040 1941.590 17.100 ;
      LAYER via ;
        RECT 1896.220 288.020 1896.480 288.280 ;
        RECT 1900.820 288.020 1901.080 288.280 ;
        RECT 1900.820 17.040 1901.080 17.300 ;
        RECT 1941.300 17.040 1941.560 17.300 ;
      LAYER met2 ;
        RECT 1896.220 300.000 1896.500 304.000 ;
        RECT 1896.280 288.310 1896.420 300.000 ;
        RECT 1896.220 287.990 1896.480 288.310 ;
        RECT 1900.820 287.990 1901.080 288.310 ;
        RECT 1900.880 17.330 1901.020 287.990 ;
        RECT 1900.820 17.010 1901.080 17.330 ;
        RECT 1941.300 17.010 1941.560 17.330 ;
        RECT 1941.360 2.400 1941.500 17.010 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1910.910 19.620 1911.230 19.680 ;
        RECT 1958.750 19.620 1959.070 19.680 ;
        RECT 1910.910 19.480 1959.070 19.620 ;
        RECT 1910.910 19.420 1911.230 19.480 ;
        RECT 1958.750 19.420 1959.070 19.480 ;
      LAYER via ;
        RECT 1910.940 19.420 1911.200 19.680 ;
        RECT 1958.780 19.420 1959.040 19.680 ;
      LAYER met2 ;
        RECT 1910.940 300.000 1911.220 304.000 ;
        RECT 1911.000 19.710 1911.140 300.000 ;
        RECT 1910.940 19.390 1911.200 19.710 ;
        RECT 1958.780 19.390 1959.040 19.710 ;
        RECT 1958.840 16.050 1958.980 19.390 ;
        RECT 1958.840 15.910 1959.440 16.050 ;
        RECT 1959.300 2.400 1959.440 15.910 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1925.630 286.180 1925.950 286.240 ;
        RECT 1931.610 286.180 1931.930 286.240 ;
        RECT 1925.630 286.040 1931.930 286.180 ;
        RECT 1925.630 285.980 1925.950 286.040 ;
        RECT 1931.610 285.980 1931.930 286.040 ;
        RECT 1931.610 19.960 1931.930 20.020 ;
        RECT 1977.150 19.960 1977.470 20.020 ;
        RECT 1931.610 19.820 1977.470 19.960 ;
        RECT 1931.610 19.760 1931.930 19.820 ;
        RECT 1977.150 19.760 1977.470 19.820 ;
      LAYER via ;
        RECT 1925.660 285.980 1925.920 286.240 ;
        RECT 1931.640 285.980 1931.900 286.240 ;
        RECT 1931.640 19.760 1931.900 20.020 ;
        RECT 1977.180 19.760 1977.440 20.020 ;
      LAYER met2 ;
        RECT 1925.660 300.000 1925.940 304.000 ;
        RECT 1925.720 286.270 1925.860 300.000 ;
        RECT 1925.660 285.950 1925.920 286.270 ;
        RECT 1931.640 285.950 1931.900 286.270 ;
        RECT 1931.700 20.050 1931.840 285.950 ;
        RECT 1931.640 19.730 1931.900 20.050 ;
        RECT 1977.180 19.730 1977.440 20.050 ;
        RECT 1977.240 2.400 1977.380 19.730 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1940.350 288.220 1940.670 288.280 ;
        RECT 1945.410 288.220 1945.730 288.280 ;
        RECT 1940.350 288.080 1945.730 288.220 ;
        RECT 1940.350 288.020 1940.670 288.080 ;
        RECT 1945.410 288.020 1945.730 288.080 ;
        RECT 1945.410 18.600 1945.730 18.660 ;
        RECT 1995.090 18.600 1995.410 18.660 ;
        RECT 1945.410 18.460 1995.410 18.600 ;
        RECT 1945.410 18.400 1945.730 18.460 ;
        RECT 1995.090 18.400 1995.410 18.460 ;
      LAYER via ;
        RECT 1940.380 288.020 1940.640 288.280 ;
        RECT 1945.440 288.020 1945.700 288.280 ;
        RECT 1945.440 18.400 1945.700 18.660 ;
        RECT 1995.120 18.400 1995.380 18.660 ;
      LAYER met2 ;
        RECT 1940.380 300.000 1940.660 304.000 ;
        RECT 1940.440 288.310 1940.580 300.000 ;
        RECT 1940.380 287.990 1940.640 288.310 ;
        RECT 1945.440 287.990 1945.700 288.310 ;
        RECT 1945.500 18.690 1945.640 287.990 ;
        RECT 1945.440 18.370 1945.700 18.690 ;
        RECT 1995.120 18.370 1995.380 18.690 ;
        RECT 1995.180 2.400 1995.320 18.370 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1955.070 288.220 1955.390 288.280 ;
        RECT 1959.210 288.220 1959.530 288.280 ;
        RECT 1955.070 288.080 1959.530 288.220 ;
        RECT 1955.070 288.020 1955.390 288.080 ;
        RECT 1959.210 288.020 1959.530 288.080 ;
        RECT 1959.210 16.900 1959.530 16.960 ;
        RECT 2012.570 16.900 2012.890 16.960 ;
        RECT 1959.210 16.760 2012.890 16.900 ;
        RECT 1959.210 16.700 1959.530 16.760 ;
        RECT 2012.570 16.700 2012.890 16.760 ;
      LAYER via ;
        RECT 1955.100 288.020 1955.360 288.280 ;
        RECT 1959.240 288.020 1959.500 288.280 ;
        RECT 1959.240 16.700 1959.500 16.960 ;
        RECT 2012.600 16.700 2012.860 16.960 ;
      LAYER met2 ;
        RECT 1955.100 300.000 1955.380 304.000 ;
        RECT 1955.160 288.310 1955.300 300.000 ;
        RECT 1955.100 287.990 1955.360 288.310 ;
        RECT 1959.240 287.990 1959.500 288.310 ;
        RECT 1959.300 16.990 1959.440 287.990 ;
        RECT 1959.240 16.670 1959.500 16.990 ;
        RECT 2012.600 16.670 2012.860 16.990 ;
        RECT 2012.660 2.400 2012.800 16.670 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1973.010 16.220 1973.330 16.280 ;
        RECT 2030.510 16.220 2030.830 16.280 ;
        RECT 1973.010 16.080 2030.830 16.220 ;
        RECT 1973.010 16.020 1973.330 16.080 ;
        RECT 2030.510 16.020 2030.830 16.080 ;
      LAYER via ;
        RECT 1973.040 16.020 1973.300 16.280 ;
        RECT 2030.540 16.020 2030.800 16.280 ;
      LAYER met2 ;
        RECT 1969.820 300.290 1970.100 304.000 ;
        RECT 1969.820 300.150 1973.240 300.290 ;
        RECT 1969.820 300.000 1970.100 300.150 ;
        RECT 1973.100 16.310 1973.240 300.150 ;
        RECT 1973.040 15.990 1973.300 16.310 ;
        RECT 2030.540 15.990 2030.800 16.310 ;
        RECT 2030.600 2.400 2030.740 15.990 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1986.810 20.640 1987.130 20.700 ;
        RECT 2047.990 20.640 2048.310 20.700 ;
        RECT 1986.810 20.500 2048.310 20.640 ;
        RECT 1986.810 20.440 1987.130 20.500 ;
        RECT 2047.990 20.440 2048.310 20.500 ;
      LAYER via ;
        RECT 1986.840 20.440 1987.100 20.700 ;
        RECT 2048.020 20.440 2048.280 20.700 ;
      LAYER met2 ;
        RECT 1984.540 300.290 1984.820 304.000 ;
        RECT 1984.540 300.150 1987.040 300.290 ;
        RECT 1984.540 300.000 1984.820 300.150 ;
        RECT 1986.900 20.730 1987.040 300.150 ;
        RECT 1986.840 20.410 1987.100 20.730 ;
        RECT 2048.020 20.410 2048.280 20.730 ;
        RECT 2048.080 20.130 2048.220 20.410 ;
        RECT 2048.080 19.990 2048.680 20.130 ;
        RECT 2048.540 2.400 2048.680 19.990 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 780.305 285.685 780.475 288.915 ;
      LAYER mcon ;
        RECT 780.305 288.745 780.475 288.915 ;
      LAYER met1 ;
        RECT 780.245 288.900 780.535 288.945 ;
        RECT 926.510 288.900 926.830 288.960 ;
        RECT 780.245 288.760 926.830 288.900 ;
        RECT 780.245 288.715 780.535 288.760 ;
        RECT 926.510 288.700 926.830 288.760 ;
        RECT 765.510 285.840 765.830 285.900 ;
        RECT 780.245 285.840 780.535 285.885 ;
        RECT 765.510 285.700 780.535 285.840 ;
        RECT 765.510 285.640 765.830 285.700 ;
        RECT 780.245 285.655 780.535 285.700 ;
      LAYER via ;
        RECT 926.540 288.700 926.800 288.960 ;
        RECT 765.540 285.640 765.800 285.900 ;
      LAYER met2 ;
        RECT 926.540 300.000 926.820 304.000 ;
        RECT 926.600 288.990 926.740 300.000 ;
        RECT 926.540 288.670 926.800 288.990 ;
        RECT 765.540 285.610 765.800 285.930 ;
        RECT 765.600 16.730 765.740 285.610 ;
        RECT 763.760 16.590 765.740 16.730 ;
        RECT 763.760 2.400 763.900 16.590 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2000.610 18.600 2000.930 18.660 ;
        RECT 2066.390 18.600 2066.710 18.660 ;
        RECT 2000.610 18.460 2066.710 18.600 ;
        RECT 2000.610 18.400 2000.930 18.460 ;
        RECT 2066.390 18.400 2066.710 18.460 ;
      LAYER via ;
        RECT 2000.640 18.400 2000.900 18.660 ;
        RECT 2066.420 18.400 2066.680 18.660 ;
      LAYER met2 ;
        RECT 1999.260 300.290 1999.540 304.000 ;
        RECT 1999.260 300.150 2000.840 300.290 ;
        RECT 1999.260 300.000 1999.540 300.150 ;
        RECT 2000.700 18.690 2000.840 300.150 ;
        RECT 2000.640 18.370 2000.900 18.690 ;
        RECT 2066.420 18.370 2066.680 18.690 ;
        RECT 2066.480 2.400 2066.620 18.370 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2014.410 17.580 2014.730 17.640 ;
        RECT 2084.330 17.580 2084.650 17.640 ;
        RECT 2014.410 17.440 2084.650 17.580 ;
        RECT 2014.410 17.380 2014.730 17.440 ;
        RECT 2084.330 17.380 2084.650 17.440 ;
      LAYER via ;
        RECT 2014.440 17.380 2014.700 17.640 ;
        RECT 2084.360 17.380 2084.620 17.640 ;
      LAYER met2 ;
        RECT 2013.980 300.290 2014.260 304.000 ;
        RECT 2013.980 300.150 2014.640 300.290 ;
        RECT 2013.980 300.000 2014.260 300.150 ;
        RECT 2014.500 17.670 2014.640 300.150 ;
        RECT 2014.440 17.350 2014.700 17.670 ;
        RECT 2084.360 17.350 2084.620 17.670 ;
        RECT 2084.420 2.400 2084.560 17.350 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2028.670 285.500 2028.990 285.560 ;
        RECT 2034.650 285.500 2034.970 285.560 ;
        RECT 2028.670 285.360 2034.970 285.500 ;
        RECT 2028.670 285.300 2028.990 285.360 ;
        RECT 2034.650 285.300 2034.970 285.360 ;
        RECT 2034.650 16.220 2034.970 16.280 ;
        RECT 2101.810 16.220 2102.130 16.280 ;
        RECT 2034.650 16.080 2102.130 16.220 ;
        RECT 2034.650 16.020 2034.970 16.080 ;
        RECT 2101.810 16.020 2102.130 16.080 ;
      LAYER via ;
        RECT 2028.700 285.300 2028.960 285.560 ;
        RECT 2034.680 285.300 2034.940 285.560 ;
        RECT 2034.680 16.020 2034.940 16.280 ;
        RECT 2101.840 16.020 2102.100 16.280 ;
      LAYER met2 ;
        RECT 2028.700 300.000 2028.980 304.000 ;
        RECT 2028.760 285.590 2028.900 300.000 ;
        RECT 2028.700 285.270 2028.960 285.590 ;
        RECT 2034.680 285.270 2034.940 285.590 ;
        RECT 2034.740 16.310 2034.880 285.270 ;
        RECT 2034.680 15.990 2034.940 16.310 ;
        RECT 2101.840 15.990 2102.100 16.310 ;
        RECT 2101.900 2.400 2102.040 15.990 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2043.390 288.220 2043.710 288.280 ;
        RECT 2048.450 288.220 2048.770 288.280 ;
        RECT 2043.390 288.080 2048.770 288.220 ;
        RECT 2043.390 288.020 2043.710 288.080 ;
        RECT 2048.450 288.020 2048.770 288.080 ;
        RECT 2048.450 20.640 2048.770 20.700 ;
        RECT 2119.750 20.640 2120.070 20.700 ;
        RECT 2048.450 20.500 2120.070 20.640 ;
        RECT 2048.450 20.440 2048.770 20.500 ;
        RECT 2119.750 20.440 2120.070 20.500 ;
      LAYER via ;
        RECT 2043.420 288.020 2043.680 288.280 ;
        RECT 2048.480 288.020 2048.740 288.280 ;
        RECT 2048.480 20.440 2048.740 20.700 ;
        RECT 2119.780 20.440 2120.040 20.700 ;
      LAYER met2 ;
        RECT 2043.420 300.000 2043.700 304.000 ;
        RECT 2043.480 288.310 2043.620 300.000 ;
        RECT 2043.420 287.990 2043.680 288.310 ;
        RECT 2048.480 287.990 2048.740 288.310 ;
        RECT 2048.540 20.730 2048.680 287.990 ;
        RECT 2048.480 20.410 2048.740 20.730 ;
        RECT 2119.780 20.410 2120.040 20.730 ;
        RECT 2119.840 2.400 2119.980 20.410 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2058.110 288.220 2058.430 288.280 ;
        RECT 2062.250 288.220 2062.570 288.280 ;
        RECT 2058.110 288.080 2062.570 288.220 ;
        RECT 2058.110 288.020 2058.430 288.080 ;
        RECT 2062.250 288.020 2062.570 288.080 ;
        RECT 2062.250 20.300 2062.570 20.360 ;
        RECT 2137.690 20.300 2138.010 20.360 ;
        RECT 2062.250 20.160 2138.010 20.300 ;
        RECT 2062.250 20.100 2062.570 20.160 ;
        RECT 2137.690 20.100 2138.010 20.160 ;
      LAYER via ;
        RECT 2058.140 288.020 2058.400 288.280 ;
        RECT 2062.280 288.020 2062.540 288.280 ;
        RECT 2062.280 20.100 2062.540 20.360 ;
        RECT 2137.720 20.100 2137.980 20.360 ;
      LAYER met2 ;
        RECT 2058.140 300.000 2058.420 304.000 ;
        RECT 2058.200 288.310 2058.340 300.000 ;
        RECT 2058.140 287.990 2058.400 288.310 ;
        RECT 2062.280 287.990 2062.540 288.310 ;
        RECT 2062.340 20.390 2062.480 287.990 ;
        RECT 2062.280 20.070 2062.540 20.390 ;
        RECT 2137.720 20.070 2137.980 20.390 ;
        RECT 2137.780 2.400 2137.920 20.070 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2072.830 286.860 2073.150 286.920 ;
        RECT 2076.510 286.860 2076.830 286.920 ;
        RECT 2072.830 286.720 2076.830 286.860 ;
        RECT 2072.830 286.660 2073.150 286.720 ;
        RECT 2076.510 286.660 2076.830 286.720 ;
        RECT 2076.510 18.940 2076.830 19.000 ;
        RECT 2155.630 18.940 2155.950 19.000 ;
        RECT 2076.510 18.800 2155.950 18.940 ;
        RECT 2076.510 18.740 2076.830 18.800 ;
        RECT 2155.630 18.740 2155.950 18.800 ;
      LAYER via ;
        RECT 2072.860 286.660 2073.120 286.920 ;
        RECT 2076.540 286.660 2076.800 286.920 ;
        RECT 2076.540 18.740 2076.800 19.000 ;
        RECT 2155.660 18.740 2155.920 19.000 ;
      LAYER met2 ;
        RECT 2072.860 300.000 2073.140 304.000 ;
        RECT 2072.920 286.950 2073.060 300.000 ;
        RECT 2072.860 286.630 2073.120 286.950 ;
        RECT 2076.540 286.630 2076.800 286.950 ;
        RECT 2076.600 19.030 2076.740 286.630 ;
        RECT 2076.540 18.710 2076.800 19.030 ;
        RECT 2155.660 18.710 2155.920 19.030 ;
        RECT 2155.720 2.400 2155.860 18.710 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2090.310 19.280 2090.630 19.340 ;
        RECT 2172.650 19.280 2172.970 19.340 ;
        RECT 2090.310 19.140 2172.970 19.280 ;
        RECT 2090.310 19.080 2090.630 19.140 ;
        RECT 2172.650 19.080 2172.970 19.140 ;
      LAYER via ;
        RECT 2090.340 19.080 2090.600 19.340 ;
        RECT 2172.680 19.080 2172.940 19.340 ;
      LAYER met2 ;
        RECT 2087.580 300.290 2087.860 304.000 ;
        RECT 2087.580 300.150 2090.540 300.290 ;
        RECT 2087.580 300.000 2087.860 300.150 ;
        RECT 2090.400 19.370 2090.540 300.150 ;
        RECT 2090.340 19.050 2090.600 19.370 ;
        RECT 2172.680 19.050 2172.940 19.370 ;
        RECT 2172.740 18.770 2172.880 19.050 ;
        RECT 2172.740 18.630 2173.340 18.770 ;
        RECT 2173.200 2.400 2173.340 18.630 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2104.110 14.860 2104.430 14.920 ;
        RECT 2191.050 14.860 2191.370 14.920 ;
        RECT 2104.110 14.720 2191.370 14.860 ;
        RECT 2104.110 14.660 2104.430 14.720 ;
        RECT 2191.050 14.660 2191.370 14.720 ;
      LAYER via ;
        RECT 2104.140 14.660 2104.400 14.920 ;
        RECT 2191.080 14.660 2191.340 14.920 ;
      LAYER met2 ;
        RECT 2102.300 300.290 2102.580 304.000 ;
        RECT 2102.300 300.150 2104.340 300.290 ;
        RECT 2102.300 300.000 2102.580 300.150 ;
        RECT 2104.200 14.950 2104.340 300.150 ;
        RECT 2104.140 14.630 2104.400 14.950 ;
        RECT 2191.080 14.630 2191.340 14.950 ;
        RECT 2191.140 2.400 2191.280 14.630 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2117.910 17.240 2118.230 17.300 ;
        RECT 2208.990 17.240 2209.310 17.300 ;
        RECT 2117.910 17.100 2209.310 17.240 ;
        RECT 2117.910 17.040 2118.230 17.100 ;
        RECT 2208.990 17.040 2209.310 17.100 ;
      LAYER via ;
        RECT 2117.940 17.040 2118.200 17.300 ;
        RECT 2209.020 17.040 2209.280 17.300 ;
      LAYER met2 ;
        RECT 2117.020 300.290 2117.300 304.000 ;
        RECT 2117.020 300.150 2118.140 300.290 ;
        RECT 2117.020 300.000 2117.300 300.150 ;
        RECT 2118.000 17.330 2118.140 300.150 ;
        RECT 2117.940 17.010 2118.200 17.330 ;
        RECT 2209.020 17.010 2209.280 17.330 ;
        RECT 2209.080 2.400 2209.220 17.010 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2131.710 17.920 2132.030 17.980 ;
        RECT 2226.930 17.920 2227.250 17.980 ;
        RECT 2131.710 17.780 2227.250 17.920 ;
        RECT 2131.710 17.720 2132.030 17.780 ;
        RECT 2226.930 17.720 2227.250 17.780 ;
      LAYER via ;
        RECT 2131.740 17.720 2132.000 17.980 ;
        RECT 2226.960 17.720 2227.220 17.980 ;
      LAYER met2 ;
        RECT 2131.280 300.290 2131.560 304.000 ;
        RECT 2131.280 300.150 2131.940 300.290 ;
        RECT 2131.280 300.000 2131.560 300.150 ;
        RECT 2131.800 18.010 2131.940 300.150 ;
        RECT 2131.740 17.690 2132.000 18.010 ;
        RECT 2226.960 17.690 2227.220 18.010 ;
        RECT 2227.020 2.400 2227.160 17.690 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 786.210 285.840 786.530 285.900 ;
        RECT 941.230 285.840 941.550 285.900 ;
        RECT 786.210 285.700 941.550 285.840 ;
        RECT 786.210 285.640 786.530 285.700 ;
        RECT 941.230 285.640 941.550 285.700 ;
        RECT 781.610 17.240 781.930 17.300 ;
        RECT 786.210 17.240 786.530 17.300 ;
        RECT 781.610 17.100 786.530 17.240 ;
        RECT 781.610 17.040 781.930 17.100 ;
        RECT 786.210 17.040 786.530 17.100 ;
      LAYER via ;
        RECT 786.240 285.640 786.500 285.900 ;
        RECT 941.260 285.640 941.520 285.900 ;
        RECT 781.640 17.040 781.900 17.300 ;
        RECT 786.240 17.040 786.500 17.300 ;
      LAYER met2 ;
        RECT 941.260 300.000 941.540 304.000 ;
        RECT 941.320 285.930 941.460 300.000 ;
        RECT 786.240 285.610 786.500 285.930 ;
        RECT 941.260 285.610 941.520 285.930 ;
        RECT 786.300 17.330 786.440 285.610 ;
        RECT 781.640 17.010 781.900 17.330 ;
        RECT 786.240 17.010 786.500 17.330 ;
        RECT 781.700 2.400 781.840 17.010 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2145.970 287.880 2146.290 287.940 ;
        RECT 2152.410 287.880 2152.730 287.940 ;
        RECT 2145.970 287.740 2152.730 287.880 ;
        RECT 2145.970 287.680 2146.290 287.740 ;
        RECT 2152.410 287.680 2152.730 287.740 ;
        RECT 2152.410 20.300 2152.730 20.360 ;
        RECT 2244.870 20.300 2245.190 20.360 ;
        RECT 2152.410 20.160 2245.190 20.300 ;
        RECT 2152.410 20.100 2152.730 20.160 ;
        RECT 2244.870 20.100 2245.190 20.160 ;
      LAYER via ;
        RECT 2146.000 287.680 2146.260 287.940 ;
        RECT 2152.440 287.680 2152.700 287.940 ;
        RECT 2152.440 20.100 2152.700 20.360 ;
        RECT 2244.900 20.100 2245.160 20.360 ;
      LAYER met2 ;
        RECT 2146.000 300.000 2146.280 304.000 ;
        RECT 2146.060 287.970 2146.200 300.000 ;
        RECT 2146.000 287.650 2146.260 287.970 ;
        RECT 2152.440 287.650 2152.700 287.970 ;
        RECT 2152.500 20.390 2152.640 287.650 ;
        RECT 2152.440 20.070 2152.700 20.390 ;
        RECT 2244.900 20.070 2245.160 20.390 ;
        RECT 2244.960 2.400 2245.100 20.070 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2160.690 288.220 2161.010 288.280 ;
        RECT 2165.750 288.220 2166.070 288.280 ;
        RECT 2160.690 288.080 2166.070 288.220 ;
        RECT 2160.690 288.020 2161.010 288.080 ;
        RECT 2165.750 288.020 2166.070 288.080 ;
        RECT 2165.750 16.560 2166.070 16.620 ;
        RECT 2262.350 16.560 2262.670 16.620 ;
        RECT 2165.750 16.420 2262.670 16.560 ;
        RECT 2165.750 16.360 2166.070 16.420 ;
        RECT 2262.350 16.360 2262.670 16.420 ;
      LAYER via ;
        RECT 2160.720 288.020 2160.980 288.280 ;
        RECT 2165.780 288.020 2166.040 288.280 ;
        RECT 2165.780 16.360 2166.040 16.620 ;
        RECT 2262.380 16.360 2262.640 16.620 ;
      LAYER met2 ;
        RECT 2160.720 300.000 2161.000 304.000 ;
        RECT 2160.780 288.310 2160.920 300.000 ;
        RECT 2160.720 287.990 2160.980 288.310 ;
        RECT 2165.780 287.990 2166.040 288.310 ;
        RECT 2165.840 16.650 2165.980 287.990 ;
        RECT 2165.780 16.330 2166.040 16.650 ;
        RECT 2262.380 16.330 2262.640 16.650 ;
        RECT 2262.440 2.400 2262.580 16.330 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2175.410 288.220 2175.730 288.280 ;
        RECT 2180.010 288.220 2180.330 288.280 ;
        RECT 2175.410 288.080 2180.330 288.220 ;
        RECT 2175.410 288.020 2175.730 288.080 ;
        RECT 2180.010 288.020 2180.330 288.080 ;
        RECT 2180.010 14.520 2180.330 14.580 ;
        RECT 2280.290 14.520 2280.610 14.580 ;
        RECT 2180.010 14.380 2280.610 14.520 ;
        RECT 2180.010 14.320 2180.330 14.380 ;
        RECT 2280.290 14.320 2280.610 14.380 ;
      LAYER via ;
        RECT 2175.440 288.020 2175.700 288.280 ;
        RECT 2180.040 288.020 2180.300 288.280 ;
        RECT 2180.040 14.320 2180.300 14.580 ;
        RECT 2280.320 14.320 2280.580 14.580 ;
      LAYER met2 ;
        RECT 2175.440 300.000 2175.720 304.000 ;
        RECT 2175.500 288.310 2175.640 300.000 ;
        RECT 2175.440 287.990 2175.700 288.310 ;
        RECT 2180.040 287.990 2180.300 288.310 ;
        RECT 2180.100 14.610 2180.240 287.990 ;
        RECT 2180.040 14.290 2180.300 14.610 ;
        RECT 2280.320 14.290 2280.580 14.610 ;
        RECT 2280.380 2.400 2280.520 14.290 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2193.810 18.260 2194.130 18.320 ;
        RECT 2280.290 18.260 2280.610 18.320 ;
        RECT 2193.810 18.120 2280.610 18.260 ;
        RECT 2193.810 18.060 2194.130 18.120 ;
        RECT 2280.290 18.060 2280.610 18.120 ;
        RECT 2281.670 18.260 2281.990 18.320 ;
        RECT 2298.230 18.260 2298.550 18.320 ;
        RECT 2281.670 18.120 2298.550 18.260 ;
        RECT 2281.670 18.060 2281.990 18.120 ;
        RECT 2298.230 18.060 2298.550 18.120 ;
      LAYER via ;
        RECT 2193.840 18.060 2194.100 18.320 ;
        RECT 2280.320 18.060 2280.580 18.320 ;
        RECT 2281.700 18.060 2281.960 18.320 ;
        RECT 2298.260 18.060 2298.520 18.320 ;
      LAYER met2 ;
        RECT 2190.160 300.290 2190.440 304.000 ;
        RECT 2190.160 300.150 2194.040 300.290 ;
        RECT 2190.160 300.000 2190.440 300.150 ;
        RECT 2193.900 18.350 2194.040 300.150 ;
        RECT 2193.840 18.030 2194.100 18.350 ;
        RECT 2280.320 18.090 2280.580 18.350 ;
        RECT 2281.700 18.090 2281.960 18.350 ;
        RECT 2280.320 18.030 2281.960 18.090 ;
        RECT 2298.260 18.030 2298.520 18.350 ;
        RECT 2280.380 17.950 2281.900 18.030 ;
        RECT 2298.320 2.400 2298.460 18.030 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2280.825 17.425 2280.995 19.295 ;
      LAYER mcon ;
        RECT 2280.825 19.125 2280.995 19.295 ;
      LAYER met1 ;
        RECT 2207.610 19.620 2207.930 19.680 ;
        RECT 2207.610 19.480 2280.060 19.620 ;
        RECT 2207.610 19.420 2207.930 19.480 ;
        RECT 2279.920 19.280 2280.060 19.480 ;
        RECT 2280.765 19.280 2281.055 19.325 ;
        RECT 2279.920 19.140 2281.055 19.280 ;
        RECT 2280.765 19.095 2281.055 19.140 ;
        RECT 2280.765 17.580 2281.055 17.625 ;
        RECT 2316.170 17.580 2316.490 17.640 ;
        RECT 2280.765 17.440 2316.490 17.580 ;
        RECT 2280.765 17.395 2281.055 17.440 ;
        RECT 2316.170 17.380 2316.490 17.440 ;
      LAYER via ;
        RECT 2207.640 19.420 2207.900 19.680 ;
        RECT 2316.200 17.380 2316.460 17.640 ;
      LAYER met2 ;
        RECT 2204.880 300.290 2205.160 304.000 ;
        RECT 2204.880 300.150 2207.840 300.290 ;
        RECT 2204.880 300.000 2205.160 300.150 ;
        RECT 2207.700 19.710 2207.840 300.150 ;
        RECT 2207.640 19.390 2207.900 19.710 ;
        RECT 2316.200 17.350 2316.460 17.670 ;
        RECT 2316.260 2.400 2316.400 17.350 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2221.410 16.220 2221.730 16.280 ;
        RECT 2334.110 16.220 2334.430 16.280 ;
        RECT 2221.410 16.080 2334.430 16.220 ;
        RECT 2221.410 16.020 2221.730 16.080 ;
        RECT 2334.110 16.020 2334.430 16.080 ;
      LAYER via ;
        RECT 2221.440 16.020 2221.700 16.280 ;
        RECT 2334.140 16.020 2334.400 16.280 ;
      LAYER met2 ;
        RECT 2219.600 300.290 2219.880 304.000 ;
        RECT 2219.600 300.150 2221.640 300.290 ;
        RECT 2219.600 300.000 2219.880 300.150 ;
        RECT 2221.500 16.310 2221.640 300.150 ;
        RECT 2221.440 15.990 2221.700 16.310 ;
        RECT 2334.140 15.990 2334.400 16.310 ;
        RECT 2334.200 2.400 2334.340 15.990 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2235.210 18.600 2235.530 18.660 ;
        RECT 2235.210 18.460 2280.980 18.600 ;
        RECT 2235.210 18.400 2235.530 18.460 ;
        RECT 2280.840 17.920 2280.980 18.460 ;
        RECT 2351.590 17.920 2351.910 17.980 ;
        RECT 2280.840 17.780 2351.910 17.920 ;
        RECT 2351.590 17.720 2351.910 17.780 ;
      LAYER via ;
        RECT 2235.240 18.400 2235.500 18.660 ;
        RECT 2351.620 17.720 2351.880 17.980 ;
      LAYER met2 ;
        RECT 2234.320 300.290 2234.600 304.000 ;
        RECT 2234.320 300.150 2235.440 300.290 ;
        RECT 2234.320 300.000 2234.600 300.150 ;
        RECT 2235.300 18.690 2235.440 300.150 ;
        RECT 2235.240 18.370 2235.500 18.690 ;
        RECT 2351.620 17.690 2351.880 18.010 ;
        RECT 2351.680 2.400 2351.820 17.690 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2249.010 19.960 2249.330 20.020 ;
        RECT 2369.530 19.960 2369.850 20.020 ;
        RECT 2249.010 19.820 2369.850 19.960 ;
        RECT 2249.010 19.760 2249.330 19.820 ;
        RECT 2369.530 19.760 2369.850 19.820 ;
      LAYER via ;
        RECT 2249.040 19.760 2249.300 20.020 ;
        RECT 2369.560 19.760 2369.820 20.020 ;
      LAYER met2 ;
        RECT 2249.040 300.000 2249.320 304.000 ;
        RECT 2249.100 20.050 2249.240 300.000 ;
        RECT 2249.040 19.730 2249.300 20.050 ;
        RECT 2369.560 19.730 2369.820 20.050 ;
        RECT 2369.620 2.400 2369.760 19.730 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2281.285 18.445 2281.455 20.995 ;
        RECT 2286.805 16.745 2286.975 18.615 ;
        RECT 2304.285 14.025 2304.455 16.915 ;
      LAYER mcon ;
        RECT 2281.285 20.825 2281.455 20.995 ;
        RECT 2286.805 18.445 2286.975 18.615 ;
        RECT 2304.285 16.745 2304.455 16.915 ;
      LAYER met1 ;
        RECT 2263.730 288.220 2264.050 288.280 ;
        RECT 2269.710 288.220 2270.030 288.280 ;
        RECT 2263.730 288.080 2270.030 288.220 ;
        RECT 2263.730 288.020 2264.050 288.080 ;
        RECT 2269.710 288.020 2270.030 288.080 ;
        RECT 2269.710 20.980 2270.030 21.040 ;
        RECT 2281.225 20.980 2281.515 21.025 ;
        RECT 2269.710 20.840 2281.515 20.980 ;
        RECT 2269.710 20.780 2270.030 20.840 ;
        RECT 2281.225 20.795 2281.515 20.840 ;
        RECT 2281.225 18.600 2281.515 18.645 ;
        RECT 2286.745 18.600 2287.035 18.645 ;
        RECT 2281.225 18.460 2287.035 18.600 ;
        RECT 2281.225 18.415 2281.515 18.460 ;
        RECT 2286.745 18.415 2287.035 18.460 ;
        RECT 2286.745 16.900 2287.035 16.945 ;
        RECT 2304.225 16.900 2304.515 16.945 ;
        RECT 2286.745 16.760 2304.515 16.900 ;
        RECT 2286.745 16.715 2287.035 16.760 ;
        RECT 2304.225 16.715 2304.515 16.760 ;
        RECT 2304.225 14.180 2304.515 14.225 ;
        RECT 2387.470 14.180 2387.790 14.240 ;
        RECT 2304.225 14.040 2387.790 14.180 ;
        RECT 2304.225 13.995 2304.515 14.040 ;
        RECT 2387.470 13.980 2387.790 14.040 ;
      LAYER via ;
        RECT 2263.760 288.020 2264.020 288.280 ;
        RECT 2269.740 288.020 2270.000 288.280 ;
        RECT 2269.740 20.780 2270.000 21.040 ;
        RECT 2387.500 13.980 2387.760 14.240 ;
      LAYER met2 ;
        RECT 2263.760 300.000 2264.040 304.000 ;
        RECT 2263.820 288.310 2263.960 300.000 ;
        RECT 2263.760 287.990 2264.020 288.310 ;
        RECT 2269.740 287.990 2270.000 288.310 ;
        RECT 2269.800 21.070 2269.940 287.990 ;
        RECT 2269.740 20.750 2270.000 21.070 ;
        RECT 2387.500 13.950 2387.760 14.270 ;
        RECT 2387.560 2.400 2387.700 13.950 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2310.725 16.745 2310.895 19.295 ;
      LAYER mcon ;
        RECT 2310.725 19.125 2310.895 19.295 ;
      LAYER met1 ;
        RECT 2278.450 288.220 2278.770 288.280 ;
        RECT 2283.510 288.220 2283.830 288.280 ;
        RECT 2278.450 288.080 2283.830 288.220 ;
        RECT 2278.450 288.020 2278.770 288.080 ;
        RECT 2283.510 288.020 2283.830 288.080 ;
        RECT 2283.510 19.280 2283.830 19.340 ;
        RECT 2310.665 19.280 2310.955 19.325 ;
        RECT 2283.510 19.140 2310.955 19.280 ;
        RECT 2283.510 19.080 2283.830 19.140 ;
        RECT 2310.665 19.095 2310.955 19.140 ;
        RECT 2310.665 16.900 2310.955 16.945 ;
        RECT 2405.410 16.900 2405.730 16.960 ;
        RECT 2310.665 16.760 2405.730 16.900 ;
        RECT 2310.665 16.715 2310.955 16.760 ;
        RECT 2405.410 16.700 2405.730 16.760 ;
      LAYER via ;
        RECT 2278.480 288.020 2278.740 288.280 ;
        RECT 2283.540 288.020 2283.800 288.280 ;
        RECT 2283.540 19.080 2283.800 19.340 ;
        RECT 2405.440 16.700 2405.700 16.960 ;
      LAYER met2 ;
        RECT 2278.480 300.000 2278.760 304.000 ;
        RECT 2278.540 288.310 2278.680 300.000 ;
        RECT 2278.480 287.990 2278.740 288.310 ;
        RECT 2283.540 287.990 2283.800 288.310 ;
        RECT 2283.600 19.370 2283.740 287.990 ;
        RECT 2283.540 19.050 2283.800 19.370 ;
        RECT 2405.440 16.670 2405.700 16.990 ;
        RECT 2405.500 2.400 2405.640 16.670 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 800.010 285.500 800.330 285.560 ;
        RECT 955.950 285.500 956.270 285.560 ;
        RECT 800.010 285.360 956.270 285.500 ;
        RECT 800.010 285.300 800.330 285.360 ;
        RECT 955.950 285.300 956.270 285.360 ;
      LAYER via ;
        RECT 800.040 285.300 800.300 285.560 ;
        RECT 955.980 285.300 956.240 285.560 ;
      LAYER met2 ;
        RECT 955.980 300.000 956.260 304.000 ;
        RECT 956.040 285.590 956.180 300.000 ;
        RECT 800.040 285.270 800.300 285.590 ;
        RECT 955.980 285.270 956.240 285.590 ;
        RECT 800.100 17.410 800.240 285.270 ;
        RECT 799.640 17.270 800.240 17.410 ;
        RECT 799.640 2.400 799.780 17.270 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 644.990 24.040 645.310 24.100 ;
        RECT 828.530 24.040 828.850 24.100 ;
        RECT 644.990 23.900 828.850 24.040 ;
        RECT 644.990 23.840 645.310 23.900 ;
        RECT 828.530 23.840 828.850 23.900 ;
      LAYER via ;
        RECT 645.020 23.840 645.280 24.100 ;
        RECT 828.560 23.840 828.820 24.100 ;
      LAYER met2 ;
        RECT 828.560 300.000 828.840 304.000 ;
        RECT 828.620 24.130 828.760 300.000 ;
        RECT 645.020 23.810 645.280 24.130 ;
        RECT 828.560 23.810 828.820 24.130 ;
        RECT 645.080 2.400 645.220 23.810 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2297.770 288.220 2298.090 288.280 ;
        RECT 2304.210 288.220 2304.530 288.280 ;
        RECT 2297.770 288.080 2304.530 288.220 ;
        RECT 2297.770 288.020 2298.090 288.080 ;
        RECT 2304.210 288.020 2304.530 288.080 ;
        RECT 2304.210 18.260 2304.530 18.320 ;
        RECT 2428.870 18.260 2429.190 18.320 ;
        RECT 2304.210 18.120 2429.190 18.260 ;
        RECT 2304.210 18.060 2304.530 18.120 ;
        RECT 2428.870 18.060 2429.190 18.120 ;
      LAYER via ;
        RECT 2297.800 288.020 2298.060 288.280 ;
        RECT 2304.240 288.020 2304.500 288.280 ;
        RECT 2304.240 18.060 2304.500 18.320 ;
        RECT 2428.900 18.060 2429.160 18.320 ;
      LAYER met2 ;
        RECT 2297.800 300.000 2298.080 304.000 ;
        RECT 2297.860 288.310 2298.000 300.000 ;
        RECT 2297.800 287.990 2298.060 288.310 ;
        RECT 2304.240 287.990 2304.500 288.310 ;
        RECT 2304.300 18.350 2304.440 287.990 ;
        RECT 2304.240 18.030 2304.500 18.350 ;
        RECT 2428.900 18.030 2429.160 18.350 ;
        RECT 2428.960 2.400 2429.100 18.030 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2329.125 15.725 2329.295 17.255 ;
        RECT 2346.605 14.705 2346.775 16.235 ;
      LAYER mcon ;
        RECT 2329.125 17.085 2329.295 17.255 ;
        RECT 2346.605 16.065 2346.775 16.235 ;
      LAYER met1 ;
        RECT 2312.490 288.220 2312.810 288.280 ;
        RECT 2318.010 288.220 2318.330 288.280 ;
        RECT 2312.490 288.080 2318.330 288.220 ;
        RECT 2312.490 288.020 2312.810 288.080 ;
        RECT 2318.010 288.020 2318.330 288.080 ;
        RECT 2318.010 17.580 2318.330 17.640 ;
        RECT 2318.010 17.440 2328.820 17.580 ;
        RECT 2318.010 17.380 2318.330 17.440 ;
        RECT 2328.680 17.240 2328.820 17.440 ;
        RECT 2329.065 17.240 2329.355 17.285 ;
        RECT 2328.680 17.100 2329.355 17.240 ;
        RECT 2329.065 17.055 2329.355 17.100 ;
        RECT 2346.545 16.220 2346.835 16.265 ;
        RECT 2335.120 16.080 2346.835 16.220 ;
        RECT 2329.065 15.880 2329.355 15.925 ;
        RECT 2335.120 15.880 2335.260 16.080 ;
        RECT 2346.545 16.035 2346.835 16.080 ;
        RECT 2329.065 15.740 2335.260 15.880 ;
        RECT 2329.065 15.695 2329.355 15.740 ;
        RECT 2346.545 14.860 2346.835 14.905 ;
        RECT 2446.810 14.860 2447.130 14.920 ;
        RECT 2346.545 14.720 2447.130 14.860 ;
        RECT 2346.545 14.675 2346.835 14.720 ;
        RECT 2446.810 14.660 2447.130 14.720 ;
      LAYER via ;
        RECT 2312.520 288.020 2312.780 288.280 ;
        RECT 2318.040 288.020 2318.300 288.280 ;
        RECT 2318.040 17.380 2318.300 17.640 ;
        RECT 2446.840 14.660 2447.100 14.920 ;
      LAYER met2 ;
        RECT 2312.520 300.000 2312.800 304.000 ;
        RECT 2312.580 288.310 2312.720 300.000 ;
        RECT 2312.520 287.990 2312.780 288.310 ;
        RECT 2318.040 287.990 2318.300 288.310 ;
        RECT 2318.100 17.670 2318.240 287.990 ;
        RECT 2318.040 17.350 2318.300 17.670 ;
        RECT 2446.840 14.630 2447.100 14.950 ;
        RECT 2446.900 2.400 2447.040 14.630 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2327.210 288.220 2327.530 288.280 ;
        RECT 2331.810 288.220 2332.130 288.280 ;
        RECT 2327.210 288.080 2332.130 288.220 ;
        RECT 2327.210 288.020 2327.530 288.080 ;
        RECT 2331.810 288.020 2332.130 288.080 ;
        RECT 2464.750 17.580 2465.070 17.640 ;
        RECT 2376.980 17.440 2465.070 17.580 ;
        RECT 2331.810 17.240 2332.130 17.300 ;
        RECT 2376.980 17.240 2377.120 17.440 ;
        RECT 2464.750 17.380 2465.070 17.440 ;
        RECT 2331.810 17.100 2377.120 17.240 ;
        RECT 2331.810 17.040 2332.130 17.100 ;
      LAYER via ;
        RECT 2327.240 288.020 2327.500 288.280 ;
        RECT 2331.840 288.020 2332.100 288.280 ;
        RECT 2331.840 17.040 2332.100 17.300 ;
        RECT 2464.780 17.380 2465.040 17.640 ;
      LAYER met2 ;
        RECT 2327.240 300.000 2327.520 304.000 ;
        RECT 2327.300 288.310 2327.440 300.000 ;
        RECT 2327.240 287.990 2327.500 288.310 ;
        RECT 2331.840 287.990 2332.100 288.310 ;
        RECT 2331.900 17.330 2332.040 287.990 ;
        RECT 2464.780 17.350 2465.040 17.670 ;
        RECT 2331.840 17.010 2332.100 17.330 ;
        RECT 2464.840 2.400 2464.980 17.350 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2345.610 15.680 2345.930 15.940 ;
        RECT 2345.700 15.540 2345.840 15.680 ;
        RECT 2482.690 15.540 2483.010 15.600 ;
        RECT 2345.700 15.400 2483.010 15.540 ;
        RECT 2482.690 15.340 2483.010 15.400 ;
      LAYER via ;
        RECT 2345.640 15.680 2345.900 15.940 ;
        RECT 2482.720 15.340 2482.980 15.600 ;
      LAYER met2 ;
        RECT 2341.960 300.290 2342.240 304.000 ;
        RECT 2341.960 300.150 2345.840 300.290 ;
        RECT 2341.960 300.000 2342.240 300.150 ;
        RECT 2345.700 15.970 2345.840 300.150 ;
        RECT 2345.640 15.650 2345.900 15.970 ;
        RECT 2482.720 15.310 2482.980 15.630 ;
        RECT 2482.780 2.400 2482.920 15.310 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2380.645 17.085 2380.815 18.955 ;
      LAYER mcon ;
        RECT 2380.645 18.785 2380.815 18.955 ;
      LAYER met1 ;
        RECT 2359.410 18.940 2359.730 19.000 ;
        RECT 2380.585 18.940 2380.875 18.985 ;
        RECT 2359.410 18.800 2380.875 18.940 ;
        RECT 2359.410 18.740 2359.730 18.800 ;
        RECT 2380.585 18.755 2380.875 18.800 ;
        RECT 2380.585 17.240 2380.875 17.285 ;
        RECT 2500.630 17.240 2500.950 17.300 ;
        RECT 2380.585 17.100 2500.950 17.240 ;
        RECT 2380.585 17.055 2380.875 17.100 ;
        RECT 2500.630 17.040 2500.950 17.100 ;
      LAYER via ;
        RECT 2359.440 18.740 2359.700 19.000 ;
        RECT 2500.660 17.040 2500.920 17.300 ;
      LAYER met2 ;
        RECT 2356.680 300.290 2356.960 304.000 ;
        RECT 2356.680 300.150 2359.640 300.290 ;
        RECT 2356.680 300.000 2356.960 300.150 ;
        RECT 2359.500 19.030 2359.640 300.150 ;
        RECT 2359.440 18.710 2359.700 19.030 ;
        RECT 2500.660 17.010 2500.920 17.330 ;
        RECT 2500.720 2.400 2500.860 17.010 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2373.210 15.880 2373.530 15.940 ;
        RECT 2518.110 15.880 2518.430 15.940 ;
        RECT 2373.210 15.740 2518.430 15.880 ;
        RECT 2373.210 15.680 2373.530 15.740 ;
        RECT 2518.110 15.680 2518.430 15.740 ;
      LAYER via ;
        RECT 2373.240 15.680 2373.500 15.940 ;
        RECT 2518.140 15.680 2518.400 15.940 ;
      LAYER met2 ;
        RECT 2371.400 300.290 2371.680 304.000 ;
        RECT 2371.400 300.150 2373.440 300.290 ;
        RECT 2371.400 300.000 2371.680 300.150 ;
        RECT 2373.300 15.970 2373.440 300.150 ;
        RECT 2373.240 15.650 2373.500 15.970 ;
        RECT 2518.140 15.650 2518.400 15.970 ;
        RECT 2518.200 2.400 2518.340 15.650 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2386.550 19.960 2386.870 20.020 ;
        RECT 2536.050 19.960 2536.370 20.020 ;
        RECT 2386.550 19.820 2536.370 19.960 ;
        RECT 2386.550 19.760 2386.870 19.820 ;
        RECT 2536.050 19.760 2536.370 19.820 ;
      LAYER via ;
        RECT 2386.580 19.760 2386.840 20.020 ;
        RECT 2536.080 19.760 2536.340 20.020 ;
      LAYER met2 ;
        RECT 2386.120 300.290 2386.400 304.000 ;
        RECT 2386.120 300.150 2386.780 300.290 ;
        RECT 2386.120 300.000 2386.400 300.150 ;
        RECT 2386.640 20.050 2386.780 300.150 ;
        RECT 2386.580 19.730 2386.840 20.050 ;
        RECT 2536.080 19.730 2536.340 20.050 ;
        RECT 2536.140 2.400 2536.280 19.730 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2400.810 289.240 2401.130 289.300 ;
        RECT 2445.890 289.240 2446.210 289.300 ;
        RECT 2400.810 289.100 2446.210 289.240 ;
        RECT 2400.810 289.040 2401.130 289.100 ;
        RECT 2445.890 289.040 2446.210 289.100 ;
        RECT 2445.890 14.180 2446.210 14.240 ;
        RECT 2553.990 14.180 2554.310 14.240 ;
        RECT 2445.890 14.040 2554.310 14.180 ;
        RECT 2445.890 13.980 2446.210 14.040 ;
        RECT 2553.990 13.980 2554.310 14.040 ;
      LAYER via ;
        RECT 2400.840 289.040 2401.100 289.300 ;
        RECT 2445.920 289.040 2446.180 289.300 ;
        RECT 2445.920 13.980 2446.180 14.240 ;
        RECT 2554.020 13.980 2554.280 14.240 ;
      LAYER met2 ;
        RECT 2400.840 300.000 2401.120 304.000 ;
        RECT 2400.900 289.330 2401.040 300.000 ;
        RECT 2400.840 289.010 2401.100 289.330 ;
        RECT 2445.920 289.010 2446.180 289.330 ;
        RECT 2445.980 14.270 2446.120 289.010 ;
        RECT 2445.920 13.950 2446.180 14.270 ;
        RECT 2554.020 13.950 2554.280 14.270 ;
        RECT 2554.080 2.400 2554.220 13.950 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2415.530 288.900 2415.850 288.960 ;
        RECT 2421.510 288.900 2421.830 288.960 ;
        RECT 2415.530 288.760 2421.830 288.900 ;
        RECT 2415.530 288.700 2415.850 288.760 ;
        RECT 2421.510 288.700 2421.830 288.760 ;
        RECT 2421.510 20.640 2421.830 20.700 ;
        RECT 2571.930 20.640 2572.250 20.700 ;
        RECT 2421.510 20.500 2572.250 20.640 ;
        RECT 2421.510 20.440 2421.830 20.500 ;
        RECT 2571.930 20.440 2572.250 20.500 ;
      LAYER via ;
        RECT 2415.560 288.700 2415.820 288.960 ;
        RECT 2421.540 288.700 2421.800 288.960 ;
        RECT 2421.540 20.440 2421.800 20.700 ;
        RECT 2571.960 20.440 2572.220 20.700 ;
      LAYER met2 ;
        RECT 2415.560 300.000 2415.840 304.000 ;
        RECT 2415.620 288.990 2415.760 300.000 ;
        RECT 2415.560 288.670 2415.820 288.990 ;
        RECT 2421.540 288.670 2421.800 288.990 ;
        RECT 2421.600 20.730 2421.740 288.670 ;
        RECT 2421.540 20.410 2421.800 20.730 ;
        RECT 2571.960 20.410 2572.220 20.730 ;
        RECT 2572.020 2.400 2572.160 20.410 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2430.250 284.820 2430.570 284.880 ;
        RECT 2459.690 284.820 2460.010 284.880 ;
        RECT 2430.250 284.680 2460.010 284.820 ;
        RECT 2430.250 284.620 2430.570 284.680 ;
        RECT 2459.690 284.620 2460.010 284.680 ;
        RECT 2459.690 14.520 2460.010 14.580 ;
        RECT 2589.410 14.520 2589.730 14.580 ;
        RECT 2459.690 14.380 2589.730 14.520 ;
        RECT 2459.690 14.320 2460.010 14.380 ;
        RECT 2589.410 14.320 2589.730 14.380 ;
      LAYER via ;
        RECT 2430.280 284.620 2430.540 284.880 ;
        RECT 2459.720 284.620 2459.980 284.880 ;
        RECT 2459.720 14.320 2459.980 14.580 ;
        RECT 2589.440 14.320 2589.700 14.580 ;
      LAYER met2 ;
        RECT 2430.280 300.000 2430.560 304.000 ;
        RECT 2430.340 284.910 2430.480 300.000 ;
        RECT 2430.280 284.590 2430.540 284.910 ;
        RECT 2459.720 284.590 2459.980 284.910 ;
        RECT 2459.780 14.610 2459.920 284.590 ;
        RECT 2459.720 14.290 2459.980 14.610 ;
        RECT 2589.440 14.290 2589.700 14.610 ;
        RECT 2589.500 2.400 2589.640 14.290 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 827.610 284.820 827.930 284.880 ;
        RECT 975.730 284.820 976.050 284.880 ;
        RECT 827.610 284.680 976.050 284.820 ;
        RECT 827.610 284.620 827.930 284.680 ;
        RECT 975.730 284.620 976.050 284.680 ;
        RECT 823.470 17.580 823.790 17.640 ;
        RECT 827.610 17.580 827.930 17.640 ;
        RECT 823.470 17.440 827.930 17.580 ;
        RECT 823.470 17.380 823.790 17.440 ;
        RECT 827.610 17.380 827.930 17.440 ;
      LAYER via ;
        RECT 827.640 284.620 827.900 284.880 ;
        RECT 975.760 284.620 976.020 284.880 ;
        RECT 823.500 17.380 823.760 17.640 ;
        RECT 827.640 17.380 827.900 17.640 ;
      LAYER met2 ;
        RECT 975.760 300.000 976.040 304.000 ;
        RECT 975.820 284.910 975.960 300.000 ;
        RECT 827.640 284.590 827.900 284.910 ;
        RECT 975.760 284.590 976.020 284.910 ;
        RECT 827.700 17.670 827.840 284.590 ;
        RECT 823.500 17.350 823.760 17.670 ;
        RECT 827.640 17.350 827.900 17.670 ;
        RECT 823.560 2.400 823.700 17.350 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2444.970 288.900 2445.290 288.960 ;
        RECT 2449.110 288.900 2449.430 288.960 ;
        RECT 2444.970 288.760 2449.430 288.900 ;
        RECT 2444.970 288.700 2445.290 288.760 ;
        RECT 2449.110 288.700 2449.430 288.760 ;
        RECT 2449.110 19.280 2449.430 19.340 ;
        RECT 2607.350 19.280 2607.670 19.340 ;
        RECT 2449.110 19.140 2607.670 19.280 ;
        RECT 2449.110 19.080 2449.430 19.140 ;
        RECT 2607.350 19.080 2607.670 19.140 ;
      LAYER via ;
        RECT 2445.000 288.700 2445.260 288.960 ;
        RECT 2449.140 288.700 2449.400 288.960 ;
        RECT 2449.140 19.080 2449.400 19.340 ;
        RECT 2607.380 19.080 2607.640 19.340 ;
      LAYER met2 ;
        RECT 2445.000 300.000 2445.280 304.000 ;
        RECT 2445.060 288.990 2445.200 300.000 ;
        RECT 2445.000 288.670 2445.260 288.990 ;
        RECT 2449.140 288.670 2449.400 288.990 ;
        RECT 2449.200 19.370 2449.340 288.670 ;
        RECT 2449.140 19.050 2449.400 19.370 ;
        RECT 2607.380 19.050 2607.640 19.370 ;
        RECT 2607.440 2.400 2607.580 19.050 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2462.910 19.620 2463.230 19.680 ;
        RECT 2625.290 19.620 2625.610 19.680 ;
        RECT 2462.910 19.480 2625.610 19.620 ;
        RECT 2462.910 19.420 2463.230 19.480 ;
        RECT 2625.290 19.420 2625.610 19.480 ;
      LAYER via ;
        RECT 2462.940 19.420 2463.200 19.680 ;
        RECT 2625.320 19.420 2625.580 19.680 ;
      LAYER met2 ;
        RECT 2459.720 300.290 2460.000 304.000 ;
        RECT 2459.720 300.150 2463.140 300.290 ;
        RECT 2459.720 300.000 2460.000 300.150 ;
        RECT 2463.000 19.710 2463.140 300.150 ;
        RECT 2462.940 19.390 2463.200 19.710 ;
        RECT 2625.320 19.390 2625.580 19.710 ;
        RECT 2625.380 2.400 2625.520 19.390 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2474.410 285.840 2474.730 285.900 ;
        RECT 2632.190 285.840 2632.510 285.900 ;
        RECT 2474.410 285.700 2632.510 285.840 ;
        RECT 2474.410 285.640 2474.730 285.700 ;
        RECT 2632.190 285.640 2632.510 285.700 ;
        RECT 2632.190 19.960 2632.510 20.020 ;
        RECT 2643.230 19.960 2643.550 20.020 ;
        RECT 2632.190 19.820 2643.550 19.960 ;
        RECT 2632.190 19.760 2632.510 19.820 ;
        RECT 2643.230 19.760 2643.550 19.820 ;
      LAYER via ;
        RECT 2474.440 285.640 2474.700 285.900 ;
        RECT 2632.220 285.640 2632.480 285.900 ;
        RECT 2632.220 19.760 2632.480 20.020 ;
        RECT 2643.260 19.760 2643.520 20.020 ;
      LAYER met2 ;
        RECT 2474.440 300.000 2474.720 304.000 ;
        RECT 2474.500 285.930 2474.640 300.000 ;
        RECT 2474.440 285.610 2474.700 285.930 ;
        RECT 2632.220 285.610 2632.480 285.930 ;
        RECT 2632.280 20.050 2632.420 285.610 ;
        RECT 2632.220 19.730 2632.480 20.050 ;
        RECT 2643.260 19.730 2643.520 20.050 ;
        RECT 2643.320 2.400 2643.460 19.730 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2489.130 289.580 2489.450 289.640 ;
        RECT 2645.990 289.580 2646.310 289.640 ;
        RECT 2489.130 289.440 2646.310 289.580 ;
        RECT 2489.130 289.380 2489.450 289.440 ;
        RECT 2645.990 289.380 2646.310 289.440 ;
        RECT 2645.990 17.920 2646.310 17.980 ;
        RECT 2661.170 17.920 2661.490 17.980 ;
        RECT 2645.990 17.780 2661.490 17.920 ;
        RECT 2645.990 17.720 2646.310 17.780 ;
        RECT 2661.170 17.720 2661.490 17.780 ;
      LAYER via ;
        RECT 2489.160 289.380 2489.420 289.640 ;
        RECT 2646.020 289.380 2646.280 289.640 ;
        RECT 2646.020 17.720 2646.280 17.980 ;
        RECT 2661.200 17.720 2661.460 17.980 ;
      LAYER met2 ;
        RECT 2489.160 300.000 2489.440 304.000 ;
        RECT 2489.220 289.670 2489.360 300.000 ;
        RECT 2489.160 289.350 2489.420 289.670 ;
        RECT 2646.020 289.350 2646.280 289.670 ;
        RECT 2646.080 18.010 2646.220 289.350 ;
        RECT 2646.020 17.690 2646.280 18.010 ;
        RECT 2661.200 17.690 2661.460 18.010 ;
        RECT 2661.260 2.400 2661.400 17.690 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2503.850 17.240 2504.170 17.300 ;
        RECT 2678.650 17.240 2678.970 17.300 ;
        RECT 2503.850 17.100 2678.970 17.240 ;
        RECT 2503.850 17.040 2504.170 17.100 ;
        RECT 2678.650 17.040 2678.970 17.100 ;
      LAYER via ;
        RECT 2503.880 17.040 2504.140 17.300 ;
        RECT 2678.680 17.040 2678.940 17.300 ;
      LAYER met2 ;
        RECT 2503.880 300.000 2504.160 304.000 ;
        RECT 2503.940 17.330 2504.080 300.000 ;
        RECT 2503.880 17.010 2504.140 17.330 ;
        RECT 2678.680 17.010 2678.940 17.330 ;
        RECT 2678.740 2.400 2678.880 17.010 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2554.525 14.025 2554.695 15.215 ;
      LAYER mcon ;
        RECT 2554.525 15.045 2554.695 15.215 ;
      LAYER met1 ;
        RECT 2520.410 283.460 2520.730 283.520 ;
        RECT 2549.390 283.460 2549.710 283.520 ;
        RECT 2520.410 283.320 2549.710 283.460 ;
        RECT 2520.410 283.260 2520.730 283.320 ;
        RECT 2549.390 283.260 2549.710 283.320 ;
        RECT 2549.390 15.200 2549.710 15.260 ;
        RECT 2554.465 15.200 2554.755 15.245 ;
        RECT 2549.390 15.060 2554.755 15.200 ;
        RECT 2549.390 15.000 2549.710 15.060 ;
        RECT 2554.465 15.015 2554.755 15.060 ;
        RECT 2554.465 14.180 2554.755 14.225 ;
        RECT 2696.590 14.180 2696.910 14.240 ;
        RECT 2554.465 14.040 2696.910 14.180 ;
        RECT 2554.465 13.995 2554.755 14.040 ;
        RECT 2696.590 13.980 2696.910 14.040 ;
      LAYER via ;
        RECT 2520.440 283.260 2520.700 283.520 ;
        RECT 2549.420 283.260 2549.680 283.520 ;
        RECT 2549.420 15.000 2549.680 15.260 ;
        RECT 2696.620 13.980 2696.880 14.240 ;
      LAYER met2 ;
        RECT 2518.600 300.290 2518.880 304.000 ;
        RECT 2518.600 300.150 2520.640 300.290 ;
        RECT 2518.600 300.000 2518.880 300.150 ;
        RECT 2520.500 283.550 2520.640 300.150 ;
        RECT 2520.440 283.230 2520.700 283.550 ;
        RECT 2549.420 283.230 2549.680 283.550 ;
        RECT 2549.480 15.290 2549.620 283.230 ;
        RECT 2549.420 14.970 2549.680 15.290 ;
        RECT 2696.620 13.950 2696.880 14.270 ;
        RECT 2696.680 2.400 2696.820 13.950 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2533.290 287.880 2533.610 287.940 ;
        RECT 2533.290 287.740 2694.520 287.880 ;
        RECT 2533.290 287.680 2533.610 287.740 ;
        RECT 2694.380 287.540 2694.520 287.740 ;
        RECT 2711.770 287.540 2712.090 287.600 ;
        RECT 2694.380 287.400 2712.090 287.540 ;
        RECT 2711.770 287.340 2712.090 287.400 ;
        RECT 2711.770 2.960 2712.090 3.020 ;
        RECT 2714.530 2.960 2714.850 3.020 ;
        RECT 2711.770 2.820 2714.850 2.960 ;
        RECT 2711.770 2.760 2712.090 2.820 ;
        RECT 2714.530 2.760 2714.850 2.820 ;
      LAYER via ;
        RECT 2533.320 287.680 2533.580 287.940 ;
        RECT 2711.800 287.340 2712.060 287.600 ;
        RECT 2711.800 2.760 2712.060 3.020 ;
        RECT 2714.560 2.760 2714.820 3.020 ;
      LAYER met2 ;
        RECT 2533.320 300.000 2533.600 304.000 ;
        RECT 2533.380 287.970 2533.520 300.000 ;
        RECT 2533.320 287.650 2533.580 287.970 ;
        RECT 2711.800 287.310 2712.060 287.630 ;
        RECT 2711.860 3.050 2712.000 287.310 ;
        RECT 2711.800 2.730 2712.060 3.050 ;
        RECT 2714.560 2.730 2714.820 3.050 ;
        RECT 2714.620 2.400 2714.760 2.730 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2693.905 285.685 2694.075 287.555 ;
      LAYER mcon ;
        RECT 2693.905 287.385 2694.075 287.555 ;
      LAYER met1 ;
        RECT 2547.550 287.540 2547.870 287.600 ;
        RECT 2693.845 287.540 2694.135 287.585 ;
        RECT 2547.550 287.400 2694.135 287.540 ;
        RECT 2547.550 287.340 2547.870 287.400 ;
        RECT 2693.845 287.355 2694.135 287.400 ;
        RECT 2693.845 285.840 2694.135 285.885 ;
        RECT 2728.790 285.840 2729.110 285.900 ;
        RECT 2693.845 285.700 2729.110 285.840 ;
        RECT 2693.845 285.655 2694.135 285.700 ;
        RECT 2728.790 285.640 2729.110 285.700 ;
        RECT 2728.790 15.880 2729.110 15.940 ;
        RECT 2732.470 15.880 2732.790 15.940 ;
        RECT 2728.790 15.740 2732.790 15.880 ;
        RECT 2728.790 15.680 2729.110 15.740 ;
        RECT 2732.470 15.680 2732.790 15.740 ;
      LAYER via ;
        RECT 2547.580 287.340 2547.840 287.600 ;
        RECT 2728.820 285.640 2729.080 285.900 ;
        RECT 2728.820 15.680 2729.080 15.940 ;
        RECT 2732.500 15.680 2732.760 15.940 ;
      LAYER met2 ;
        RECT 2547.580 300.000 2547.860 304.000 ;
        RECT 2547.640 287.630 2547.780 300.000 ;
        RECT 2547.580 287.310 2547.840 287.630 ;
        RECT 2728.820 285.610 2729.080 285.930 ;
        RECT 2728.880 15.970 2729.020 285.610 ;
        RECT 2728.820 15.650 2729.080 15.970 ;
        RECT 2732.500 15.650 2732.760 15.970 ;
        RECT 2732.560 2.400 2732.700 15.650 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2562.270 288.560 2562.590 288.620 ;
        RECT 2735.690 288.560 2736.010 288.620 ;
        RECT 2562.270 288.420 2736.010 288.560 ;
        RECT 2562.270 288.360 2562.590 288.420 ;
        RECT 2735.690 288.360 2736.010 288.420 ;
        RECT 2735.690 15.880 2736.010 15.940 ;
        RECT 2750.410 15.880 2750.730 15.940 ;
        RECT 2735.690 15.740 2750.730 15.880 ;
        RECT 2735.690 15.680 2736.010 15.740 ;
        RECT 2750.410 15.680 2750.730 15.740 ;
      LAYER via ;
        RECT 2562.300 288.360 2562.560 288.620 ;
        RECT 2735.720 288.360 2735.980 288.620 ;
        RECT 2735.720 15.680 2735.980 15.940 ;
        RECT 2750.440 15.680 2750.700 15.940 ;
      LAYER met2 ;
        RECT 2562.300 300.000 2562.580 304.000 ;
        RECT 2562.360 288.650 2562.500 300.000 ;
        RECT 2562.300 288.330 2562.560 288.650 ;
        RECT 2735.720 288.330 2735.980 288.650 ;
        RECT 2735.780 15.970 2735.920 288.330 ;
        RECT 2735.720 15.650 2735.980 15.970 ;
        RECT 2750.440 15.650 2750.700 15.970 ;
        RECT 2750.500 2.400 2750.640 15.650 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2576.990 288.220 2577.310 288.280 ;
        RECT 2749.490 288.220 2749.810 288.280 ;
        RECT 2576.990 288.080 2749.810 288.220 ;
        RECT 2576.990 288.020 2577.310 288.080 ;
        RECT 2749.490 288.020 2749.810 288.080 ;
        RECT 2749.490 16.900 2749.810 16.960 ;
        RECT 2767.890 16.900 2768.210 16.960 ;
        RECT 2749.490 16.760 2768.210 16.900 ;
        RECT 2749.490 16.700 2749.810 16.760 ;
        RECT 2767.890 16.700 2768.210 16.760 ;
      LAYER via ;
        RECT 2577.020 288.020 2577.280 288.280 ;
        RECT 2749.520 288.020 2749.780 288.280 ;
        RECT 2749.520 16.700 2749.780 16.960 ;
        RECT 2767.920 16.700 2768.180 16.960 ;
      LAYER met2 ;
        RECT 2577.020 300.000 2577.300 304.000 ;
        RECT 2577.080 288.310 2577.220 300.000 ;
        RECT 2577.020 287.990 2577.280 288.310 ;
        RECT 2749.520 287.990 2749.780 288.310 ;
        RECT 2749.580 16.990 2749.720 287.990 ;
        RECT 2749.520 16.670 2749.780 16.990 ;
        RECT 2767.920 16.670 2768.180 16.990 ;
        RECT 2767.980 2.400 2768.120 16.670 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 840.950 286.180 841.270 286.240 ;
        RECT 990.450 286.180 990.770 286.240 ;
        RECT 840.950 286.040 990.770 286.180 ;
        RECT 840.950 285.980 841.270 286.040 ;
        RECT 990.450 285.980 990.770 286.040 ;
      LAYER via ;
        RECT 840.980 285.980 841.240 286.240 ;
        RECT 990.480 285.980 990.740 286.240 ;
      LAYER met2 ;
        RECT 990.480 300.000 990.760 304.000 ;
        RECT 990.540 286.270 990.680 300.000 ;
        RECT 840.980 285.950 841.240 286.270 ;
        RECT 990.480 285.950 990.740 286.270 ;
        RECT 841.040 2.400 841.180 285.950 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2594.010 16.560 2594.330 16.620 ;
        RECT 2785.830 16.560 2786.150 16.620 ;
        RECT 2594.010 16.420 2786.150 16.560 ;
        RECT 2594.010 16.360 2594.330 16.420 ;
        RECT 2785.830 16.360 2786.150 16.420 ;
      LAYER via ;
        RECT 2594.040 16.360 2594.300 16.620 ;
        RECT 2785.860 16.360 2786.120 16.620 ;
      LAYER met2 ;
        RECT 2591.740 300.290 2592.020 304.000 ;
        RECT 2591.740 300.150 2594.240 300.290 ;
        RECT 2591.740 300.000 2592.020 300.150 ;
        RECT 2594.100 16.650 2594.240 300.150 ;
        RECT 2594.040 16.330 2594.300 16.650 ;
        RECT 2785.860 16.330 2786.120 16.650 ;
        RECT 2785.920 2.400 2786.060 16.330 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2607.810 18.940 2608.130 19.000 ;
        RECT 2803.770 18.940 2804.090 19.000 ;
        RECT 2607.810 18.800 2804.090 18.940 ;
        RECT 2607.810 18.740 2608.130 18.800 ;
        RECT 2803.770 18.740 2804.090 18.800 ;
      LAYER via ;
        RECT 2607.840 18.740 2608.100 19.000 ;
        RECT 2803.800 18.740 2804.060 19.000 ;
      LAYER met2 ;
        RECT 2606.460 300.290 2606.740 304.000 ;
        RECT 2606.460 300.150 2607.580 300.290 ;
        RECT 2606.460 300.000 2606.740 300.150 ;
        RECT 2607.440 26.930 2607.580 300.150 ;
        RECT 2607.440 26.790 2608.040 26.930 ;
        RECT 2607.900 19.030 2608.040 26.790 ;
        RECT 2607.840 18.710 2608.100 19.030 ;
        RECT 2803.800 18.710 2804.060 19.030 ;
        RECT 2803.860 2.400 2804.000 18.710 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2666.765 18.445 2666.935 19.295 ;
      LAYER mcon ;
        RECT 2666.765 19.125 2666.935 19.295 ;
      LAYER met1 ;
        RECT 2666.705 19.280 2666.995 19.325 ;
        RECT 2821.710 19.280 2822.030 19.340 ;
        RECT 2666.705 19.140 2822.030 19.280 ;
        RECT 2666.705 19.095 2666.995 19.140 ;
        RECT 2821.710 19.080 2822.030 19.140 ;
        RECT 2621.150 18.600 2621.470 18.660 ;
        RECT 2666.705 18.600 2666.995 18.645 ;
        RECT 2621.150 18.460 2666.995 18.600 ;
        RECT 2621.150 18.400 2621.470 18.460 ;
        RECT 2666.705 18.415 2666.995 18.460 ;
      LAYER via ;
        RECT 2821.740 19.080 2822.000 19.340 ;
        RECT 2621.180 18.400 2621.440 18.660 ;
      LAYER met2 ;
        RECT 2621.180 300.000 2621.460 304.000 ;
        RECT 2621.240 18.690 2621.380 300.000 ;
        RECT 2821.740 19.050 2822.000 19.370 ;
        RECT 2621.180 18.370 2621.440 18.690 ;
        RECT 2821.800 2.400 2821.940 19.050 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2635.870 289.240 2636.190 289.300 ;
        RECT 2642.310 289.240 2642.630 289.300 ;
        RECT 2635.870 289.100 2642.630 289.240 ;
        RECT 2635.870 289.040 2636.190 289.100 ;
        RECT 2642.310 289.040 2642.630 289.100 ;
        RECT 2642.310 19.620 2642.630 19.680 ;
        RECT 2839.190 19.620 2839.510 19.680 ;
        RECT 2642.310 19.480 2839.510 19.620 ;
        RECT 2642.310 19.420 2642.630 19.480 ;
        RECT 2839.190 19.420 2839.510 19.480 ;
      LAYER via ;
        RECT 2635.900 289.040 2636.160 289.300 ;
        RECT 2642.340 289.040 2642.600 289.300 ;
        RECT 2642.340 19.420 2642.600 19.680 ;
        RECT 2839.220 19.420 2839.480 19.680 ;
      LAYER met2 ;
        RECT 2635.900 300.000 2636.180 304.000 ;
        RECT 2635.960 289.330 2636.100 300.000 ;
        RECT 2635.900 289.010 2636.160 289.330 ;
        RECT 2642.340 289.010 2642.600 289.330 ;
        RECT 2642.400 19.710 2642.540 289.010 ;
        RECT 2642.340 19.390 2642.600 19.710 ;
        RECT 2839.220 19.390 2839.480 19.710 ;
        RECT 2839.280 2.400 2839.420 19.390 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2667.225 18.445 2667.395 20.315 ;
      LAYER mcon ;
        RECT 2667.225 20.145 2667.395 20.315 ;
      LAYER met1 ;
        RECT 2650.590 288.900 2650.910 288.960 ;
        RECT 2656.110 288.900 2656.430 288.960 ;
        RECT 2650.590 288.760 2656.430 288.900 ;
        RECT 2650.590 288.700 2650.910 288.760 ;
        RECT 2656.110 288.700 2656.430 288.760 ;
        RECT 2656.110 20.300 2656.430 20.360 ;
        RECT 2667.165 20.300 2667.455 20.345 ;
        RECT 2656.110 20.160 2667.455 20.300 ;
        RECT 2656.110 20.100 2656.430 20.160 ;
        RECT 2667.165 20.115 2667.455 20.160 ;
        RECT 2667.165 18.600 2667.455 18.645 ;
        RECT 2857.130 18.600 2857.450 18.660 ;
        RECT 2667.165 18.460 2857.450 18.600 ;
        RECT 2667.165 18.415 2667.455 18.460 ;
        RECT 2857.130 18.400 2857.450 18.460 ;
      LAYER via ;
        RECT 2650.620 288.700 2650.880 288.960 ;
        RECT 2656.140 288.700 2656.400 288.960 ;
        RECT 2656.140 20.100 2656.400 20.360 ;
        RECT 2857.160 18.400 2857.420 18.660 ;
      LAYER met2 ;
        RECT 2650.620 300.000 2650.900 304.000 ;
        RECT 2650.680 288.990 2650.820 300.000 ;
        RECT 2650.620 288.670 2650.880 288.990 ;
        RECT 2656.140 288.670 2656.400 288.990 ;
        RECT 2656.200 20.390 2656.340 288.670 ;
        RECT 2656.140 20.070 2656.400 20.390 ;
        RECT 2857.160 18.370 2857.420 18.690 ;
        RECT 2857.220 2.400 2857.360 18.370 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2665.310 289.240 2665.630 289.300 ;
        RECT 2665.310 289.100 2678.420 289.240 ;
        RECT 2665.310 289.040 2665.630 289.100 ;
        RECT 2678.280 288.900 2678.420 289.100 ;
        RECT 2708.090 288.900 2708.410 288.960 ;
        RECT 2678.280 288.760 2708.410 288.900 ;
        RECT 2708.090 288.700 2708.410 288.760 ;
        RECT 2709.470 15.880 2709.790 15.940 ;
        RECT 2709.470 15.740 2727.180 15.880 ;
        RECT 2709.470 15.680 2709.790 15.740 ;
        RECT 2727.040 15.540 2727.180 15.740 ;
        RECT 2727.040 15.400 2780.540 15.540 ;
        RECT 2780.400 14.860 2780.540 15.400 ;
        RECT 2875.070 14.860 2875.390 14.920 ;
        RECT 2780.400 14.720 2875.390 14.860 ;
        RECT 2875.070 14.660 2875.390 14.720 ;
      LAYER via ;
        RECT 2665.340 289.040 2665.600 289.300 ;
        RECT 2708.120 288.700 2708.380 288.960 ;
        RECT 2709.500 15.680 2709.760 15.940 ;
        RECT 2875.100 14.660 2875.360 14.920 ;
      LAYER met2 ;
        RECT 2665.340 300.000 2665.620 304.000 ;
        RECT 2665.400 289.330 2665.540 300.000 ;
        RECT 2665.340 289.010 2665.600 289.330 ;
        RECT 2708.120 288.670 2708.380 288.990 ;
        RECT 2708.180 24.890 2708.320 288.670 ;
        RECT 2708.180 24.750 2709.700 24.890 ;
        RECT 2709.560 15.970 2709.700 24.750 ;
        RECT 2709.500 15.650 2709.760 15.970 ;
        RECT 2875.100 14.630 2875.360 14.950 ;
        RECT 2875.160 2.400 2875.300 14.630 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2680.030 284.140 2680.350 284.200 ;
        RECT 2683.710 284.140 2684.030 284.200 ;
        RECT 2680.030 284.000 2684.030 284.140 ;
        RECT 2680.030 283.940 2680.350 284.000 ;
        RECT 2683.710 283.940 2684.030 284.000 ;
        RECT 2683.710 17.580 2684.030 17.640 ;
        RECT 2893.010 17.580 2893.330 17.640 ;
        RECT 2683.710 17.440 2893.330 17.580 ;
        RECT 2683.710 17.380 2684.030 17.440 ;
        RECT 2893.010 17.380 2893.330 17.440 ;
      LAYER via ;
        RECT 2680.060 283.940 2680.320 284.200 ;
        RECT 2683.740 283.940 2684.000 284.200 ;
        RECT 2683.740 17.380 2684.000 17.640 ;
        RECT 2893.040 17.380 2893.300 17.640 ;
      LAYER met2 ;
        RECT 2680.060 300.000 2680.340 304.000 ;
        RECT 2680.120 284.230 2680.260 300.000 ;
        RECT 2680.060 283.910 2680.320 284.230 ;
        RECT 2683.740 283.910 2684.000 284.230 ;
        RECT 2683.800 17.670 2683.940 283.910 ;
        RECT 2683.740 17.350 2684.000 17.670 ;
        RECT 2893.040 17.350 2893.300 17.670 ;
        RECT 2893.100 2.400 2893.240 17.350 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2763.365 14.705 2763.535 15.895 ;
      LAYER mcon ;
        RECT 2763.365 15.725 2763.535 15.895 ;
      LAYER met1 ;
        RECT 2694.750 287.880 2695.070 287.940 ;
        RECT 2721.890 287.880 2722.210 287.940 ;
        RECT 2694.750 287.740 2722.210 287.880 ;
        RECT 2694.750 287.680 2695.070 287.740 ;
        RECT 2721.890 287.680 2722.210 287.740 ;
        RECT 2763.305 15.880 2763.595 15.925 ;
        RECT 2910.950 15.880 2911.270 15.940 ;
        RECT 2763.305 15.740 2911.270 15.880 ;
        RECT 2763.305 15.695 2763.595 15.740 ;
        RECT 2910.950 15.680 2911.270 15.740 ;
        RECT 2721.890 14.860 2722.210 14.920 ;
        RECT 2763.305 14.860 2763.595 14.905 ;
        RECT 2721.890 14.720 2763.595 14.860 ;
        RECT 2721.890 14.660 2722.210 14.720 ;
        RECT 2763.305 14.675 2763.595 14.720 ;
      LAYER via ;
        RECT 2694.780 287.680 2695.040 287.940 ;
        RECT 2721.920 287.680 2722.180 287.940 ;
        RECT 2910.980 15.680 2911.240 15.940 ;
        RECT 2721.920 14.660 2722.180 14.920 ;
      LAYER met2 ;
        RECT 2694.780 300.000 2695.060 304.000 ;
        RECT 2694.840 287.970 2694.980 300.000 ;
        RECT 2694.780 287.650 2695.040 287.970 ;
        RECT 2721.920 287.650 2722.180 287.970 ;
        RECT 2721.980 14.950 2722.120 287.650 ;
        RECT 2910.980 15.650 2911.240 15.970 ;
        RECT 2721.920 14.630 2722.180 14.950 ;
        RECT 2911.040 2.400 2911.180 15.650 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 862.110 284.480 862.430 284.540 ;
        RECT 1005.170 284.480 1005.490 284.540 ;
        RECT 862.110 284.340 1005.490 284.480 ;
        RECT 862.110 284.280 862.430 284.340 ;
        RECT 1005.170 284.280 1005.490 284.340 ;
        RECT 858.890 15.200 859.210 15.260 ;
        RECT 862.110 15.200 862.430 15.260 ;
        RECT 858.890 15.060 862.430 15.200 ;
        RECT 858.890 15.000 859.210 15.060 ;
        RECT 862.110 15.000 862.430 15.060 ;
      LAYER via ;
        RECT 862.140 284.280 862.400 284.540 ;
        RECT 1005.200 284.280 1005.460 284.540 ;
        RECT 858.920 15.000 859.180 15.260 ;
        RECT 862.140 15.000 862.400 15.260 ;
      LAYER met2 ;
        RECT 1005.200 300.000 1005.480 304.000 ;
        RECT 1005.260 284.570 1005.400 300.000 ;
        RECT 862.140 284.250 862.400 284.570 ;
        RECT 1005.200 284.250 1005.460 284.570 ;
        RECT 862.200 15.290 862.340 284.250 ;
        RECT 858.920 14.970 859.180 15.290 ;
        RECT 862.140 14.970 862.400 15.290 ;
        RECT 858.980 2.400 859.120 14.970 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.810 288.220 883.130 288.280 ;
        RECT 1019.890 288.220 1020.210 288.280 ;
        RECT 882.810 288.080 1020.210 288.220 ;
        RECT 882.810 288.020 883.130 288.080 ;
        RECT 1019.890 288.020 1020.210 288.080 ;
        RECT 876.830 16.900 877.150 16.960 ;
        RECT 882.810 16.900 883.130 16.960 ;
        RECT 876.830 16.760 883.130 16.900 ;
        RECT 876.830 16.700 877.150 16.760 ;
        RECT 882.810 16.700 883.130 16.760 ;
      LAYER via ;
        RECT 882.840 288.020 883.100 288.280 ;
        RECT 1019.920 288.020 1020.180 288.280 ;
        RECT 876.860 16.700 877.120 16.960 ;
        RECT 882.840 16.700 883.100 16.960 ;
      LAYER met2 ;
        RECT 1019.920 300.000 1020.200 304.000 ;
        RECT 1019.980 288.310 1020.120 300.000 ;
        RECT 882.840 287.990 883.100 288.310 ;
        RECT 1019.920 287.990 1020.180 288.310 ;
        RECT 882.900 16.990 883.040 287.990 ;
        RECT 876.860 16.670 877.120 16.990 ;
        RECT 882.840 16.670 883.100 16.990 ;
        RECT 876.920 2.400 877.060 16.670 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 927.505 283.305 927.675 286.875 ;
      LAYER mcon ;
        RECT 927.505 286.705 927.675 286.875 ;
      LAYER met1 ;
        RECT 896.610 286.860 896.930 286.920 ;
        RECT 927.445 286.860 927.735 286.905 ;
        RECT 896.610 286.720 927.735 286.860 ;
        RECT 896.610 286.660 896.930 286.720 ;
        RECT 927.445 286.675 927.735 286.720 ;
        RECT 927.445 283.460 927.735 283.505 ;
        RECT 1034.610 283.460 1034.930 283.520 ;
        RECT 927.445 283.320 1034.930 283.460 ;
        RECT 927.445 283.275 927.735 283.320 ;
        RECT 1034.610 283.260 1034.930 283.320 ;
      LAYER via ;
        RECT 896.640 286.660 896.900 286.920 ;
        RECT 1034.640 283.260 1034.900 283.520 ;
      LAYER met2 ;
        RECT 1034.640 300.000 1034.920 304.000 ;
        RECT 896.640 286.630 896.900 286.950 ;
        RECT 896.700 16.730 896.840 286.630 ;
        RECT 1034.700 283.550 1034.840 300.000 ;
        RECT 1034.640 283.230 1034.900 283.550 ;
        RECT 894.860 16.590 896.840 16.730 ;
        RECT 894.860 2.400 895.000 16.590 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 956.025 288.405 956.195 289.255 ;
      LAYER mcon ;
        RECT 956.025 289.085 956.195 289.255 ;
      LAYER met1 ;
        RECT 917.310 289.240 917.630 289.300 ;
        RECT 955.965 289.240 956.255 289.285 ;
        RECT 917.310 289.100 956.255 289.240 ;
        RECT 917.310 289.040 917.630 289.100 ;
        RECT 955.965 289.055 956.255 289.100 ;
        RECT 955.965 288.560 956.255 288.605 ;
        RECT 1048.870 288.560 1049.190 288.620 ;
        RECT 955.965 288.420 1049.190 288.560 ;
        RECT 955.965 288.375 956.255 288.420 ;
        RECT 1048.870 288.360 1049.190 288.420 ;
        RECT 912.710 16.900 913.030 16.960 ;
        RECT 917.310 16.900 917.630 16.960 ;
        RECT 912.710 16.760 917.630 16.900 ;
        RECT 912.710 16.700 913.030 16.760 ;
        RECT 917.310 16.700 917.630 16.760 ;
      LAYER via ;
        RECT 917.340 289.040 917.600 289.300 ;
        RECT 1048.900 288.360 1049.160 288.620 ;
        RECT 912.740 16.700 913.000 16.960 ;
        RECT 917.340 16.700 917.600 16.960 ;
      LAYER met2 ;
        RECT 1048.900 300.000 1049.180 304.000 ;
        RECT 917.340 289.010 917.600 289.330 ;
        RECT 917.400 16.990 917.540 289.010 ;
        RECT 1048.960 288.650 1049.100 300.000 ;
        RECT 1048.900 288.330 1049.160 288.650 ;
        RECT 912.740 16.670 913.000 16.990 ;
        RECT 917.340 16.670 917.600 16.990 ;
        RECT 912.800 2.400 912.940 16.670 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 931.110 288.900 931.430 288.960 ;
        RECT 1063.590 288.900 1063.910 288.960 ;
        RECT 931.110 288.760 1063.910 288.900 ;
        RECT 931.110 288.700 931.430 288.760 ;
        RECT 1063.590 288.700 1063.910 288.760 ;
      LAYER via ;
        RECT 931.140 288.700 931.400 288.960 ;
        RECT 1063.620 288.700 1063.880 288.960 ;
      LAYER met2 ;
        RECT 1063.620 300.000 1063.900 304.000 ;
        RECT 1063.680 288.990 1063.820 300.000 ;
        RECT 931.140 288.670 931.400 288.990 ;
        RECT 1063.620 288.670 1063.880 288.990 ;
        RECT 931.200 16.730 931.340 288.670 ;
        RECT 930.280 16.590 931.340 16.730 ;
        RECT 930.280 2.400 930.420 16.590 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 951.810 289.580 952.130 289.640 ;
        RECT 1078.310 289.580 1078.630 289.640 ;
        RECT 951.810 289.440 1078.630 289.580 ;
        RECT 951.810 289.380 952.130 289.440 ;
        RECT 1078.310 289.380 1078.630 289.440 ;
        RECT 948.130 15.540 948.450 15.600 ;
        RECT 951.810 15.540 952.130 15.600 ;
        RECT 948.130 15.400 952.130 15.540 ;
        RECT 948.130 15.340 948.450 15.400 ;
        RECT 951.810 15.340 952.130 15.400 ;
      LAYER via ;
        RECT 951.840 289.380 952.100 289.640 ;
        RECT 1078.340 289.380 1078.600 289.640 ;
        RECT 948.160 15.340 948.420 15.600 ;
        RECT 951.840 15.340 952.100 15.600 ;
      LAYER met2 ;
        RECT 1078.340 300.000 1078.620 304.000 ;
        RECT 1078.400 289.670 1078.540 300.000 ;
        RECT 951.840 289.350 952.100 289.670 ;
        RECT 1078.340 289.350 1078.600 289.670 ;
        RECT 951.900 15.630 952.040 289.350 ;
        RECT 948.160 15.310 948.420 15.630 ;
        RECT 951.840 15.310 952.100 15.630 ;
        RECT 948.220 2.400 948.360 15.310 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1059.525 283.645 1059.695 287.555 ;
      LAYER mcon ;
        RECT 1059.525 287.385 1059.695 287.555 ;
      LAYER met1 ;
        RECT 1059.465 287.540 1059.755 287.585 ;
        RECT 1093.030 287.540 1093.350 287.600 ;
        RECT 1059.465 287.400 1093.350 287.540 ;
        RECT 1059.465 287.355 1059.755 287.400 ;
        RECT 1093.030 287.340 1093.350 287.400 ;
        RECT 1059.465 283.800 1059.755 283.845 ;
        RECT 1041.140 283.660 1059.755 283.800 ;
        RECT 972.510 283.120 972.830 283.180 ;
        RECT 1041.140 283.120 1041.280 283.660 ;
        RECT 1059.465 283.615 1059.755 283.660 ;
        RECT 972.510 282.980 1041.280 283.120 ;
        RECT 972.510 282.920 972.830 282.980 ;
        RECT 966.070 20.640 966.390 20.700 ;
        RECT 972.510 20.640 972.830 20.700 ;
        RECT 966.070 20.500 972.830 20.640 ;
        RECT 966.070 20.440 966.390 20.500 ;
        RECT 972.510 20.440 972.830 20.500 ;
      LAYER via ;
        RECT 1093.060 287.340 1093.320 287.600 ;
        RECT 972.540 282.920 972.800 283.180 ;
        RECT 966.100 20.440 966.360 20.700 ;
        RECT 972.540 20.440 972.800 20.700 ;
      LAYER met2 ;
        RECT 1093.060 300.000 1093.340 304.000 ;
        RECT 1093.120 287.630 1093.260 300.000 ;
        RECT 1093.060 287.310 1093.320 287.630 ;
        RECT 972.540 282.890 972.800 283.210 ;
        RECT 972.600 20.730 972.740 282.890 ;
        RECT 966.100 20.410 966.360 20.730 ;
        RECT 972.540 20.410 972.800 20.730 ;
        RECT 966.160 2.400 966.300 20.410 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1064.125 285.005 1064.295 288.915 ;
      LAYER mcon ;
        RECT 1064.125 288.745 1064.295 288.915 ;
      LAYER met1 ;
        RECT 1064.065 288.900 1064.355 288.945 ;
        RECT 1107.750 288.900 1108.070 288.960 ;
        RECT 1064.065 288.760 1108.070 288.900 ;
        RECT 1064.065 288.715 1064.355 288.760 ;
        RECT 1107.750 288.700 1108.070 288.760 ;
        RECT 986.310 285.160 986.630 285.220 ;
        RECT 1064.065 285.160 1064.355 285.205 ;
        RECT 986.310 285.020 1064.355 285.160 ;
        RECT 986.310 284.960 986.630 285.020 ;
        RECT 1064.065 284.975 1064.355 285.020 ;
        RECT 984.010 20.640 984.330 20.700 ;
        RECT 986.310 20.640 986.630 20.700 ;
        RECT 984.010 20.500 986.630 20.640 ;
        RECT 984.010 20.440 984.330 20.500 ;
        RECT 986.310 20.440 986.630 20.500 ;
      LAYER via ;
        RECT 1107.780 288.700 1108.040 288.960 ;
        RECT 986.340 284.960 986.600 285.220 ;
        RECT 984.040 20.440 984.300 20.700 ;
        RECT 986.340 20.440 986.600 20.700 ;
      LAYER met2 ;
        RECT 1107.780 300.000 1108.060 304.000 ;
        RECT 1107.840 288.990 1107.980 300.000 ;
        RECT 1107.780 288.670 1108.040 288.990 ;
        RECT 986.340 284.930 986.600 285.250 ;
        RECT 986.400 20.730 986.540 284.930 ;
        RECT 984.040 20.410 984.300 20.730 ;
        RECT 986.340 20.410 986.600 20.730 ;
        RECT 984.100 2.400 984.240 20.410 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 662.930 24.720 663.250 24.780 ;
        RECT 842.330 24.720 842.650 24.780 ;
        RECT 662.930 24.580 842.650 24.720 ;
        RECT 662.930 24.520 663.250 24.580 ;
        RECT 842.330 24.520 842.650 24.580 ;
      LAYER via ;
        RECT 662.960 24.520 663.220 24.780 ;
        RECT 842.360 24.520 842.620 24.780 ;
      LAYER met2 ;
        RECT 843.280 300.290 843.560 304.000 ;
        RECT 842.420 300.150 843.560 300.290 ;
        RECT 842.420 24.810 842.560 300.150 ;
        RECT 843.280 300.000 843.560 300.150 ;
        RECT 662.960 24.490 663.220 24.810 ;
        RECT 842.360 24.490 842.620 24.810 ;
        RECT 663.020 2.400 663.160 24.490 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.010 284.480 1007.330 284.540 ;
        RECT 1122.470 284.480 1122.790 284.540 ;
        RECT 1007.010 284.340 1122.790 284.480 ;
        RECT 1007.010 284.280 1007.330 284.340 ;
        RECT 1122.470 284.280 1122.790 284.340 ;
        RECT 1001.950 16.900 1002.270 16.960 ;
        RECT 1007.010 16.900 1007.330 16.960 ;
        RECT 1001.950 16.760 1007.330 16.900 ;
        RECT 1001.950 16.700 1002.270 16.760 ;
        RECT 1007.010 16.700 1007.330 16.760 ;
      LAYER via ;
        RECT 1007.040 284.280 1007.300 284.540 ;
        RECT 1122.500 284.280 1122.760 284.540 ;
        RECT 1001.980 16.700 1002.240 16.960 ;
        RECT 1007.040 16.700 1007.300 16.960 ;
      LAYER met2 ;
        RECT 1122.500 300.000 1122.780 304.000 ;
        RECT 1122.560 284.570 1122.700 300.000 ;
        RECT 1007.040 284.250 1007.300 284.570 ;
        RECT 1122.500 284.250 1122.760 284.570 ;
        RECT 1007.100 16.990 1007.240 284.250 ;
        RECT 1001.980 16.670 1002.240 16.990 ;
        RECT 1007.040 16.670 1007.300 16.990 ;
        RECT 1002.040 2.400 1002.180 16.670 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1020.810 288.220 1021.130 288.280 ;
        RECT 1137.190 288.220 1137.510 288.280 ;
        RECT 1020.810 288.080 1137.510 288.220 ;
        RECT 1020.810 288.020 1021.130 288.080 ;
        RECT 1137.190 288.020 1137.510 288.080 ;
        RECT 1018.510 65.860 1018.830 65.920 ;
        RECT 1020.810 65.860 1021.130 65.920 ;
        RECT 1018.510 65.720 1021.130 65.860 ;
        RECT 1018.510 65.660 1018.830 65.720 ;
        RECT 1020.810 65.660 1021.130 65.720 ;
        RECT 1018.510 2.960 1018.830 3.020 ;
        RECT 1019.430 2.960 1019.750 3.020 ;
        RECT 1018.510 2.820 1019.750 2.960 ;
        RECT 1018.510 2.760 1018.830 2.820 ;
        RECT 1019.430 2.760 1019.750 2.820 ;
      LAYER via ;
        RECT 1020.840 288.020 1021.100 288.280 ;
        RECT 1137.220 288.020 1137.480 288.280 ;
        RECT 1018.540 65.660 1018.800 65.920 ;
        RECT 1020.840 65.660 1021.100 65.920 ;
        RECT 1018.540 2.760 1018.800 3.020 ;
        RECT 1019.460 2.760 1019.720 3.020 ;
      LAYER met2 ;
        RECT 1137.220 300.000 1137.500 304.000 ;
        RECT 1137.280 288.310 1137.420 300.000 ;
        RECT 1020.840 287.990 1021.100 288.310 ;
        RECT 1137.220 287.990 1137.480 288.310 ;
        RECT 1020.900 65.950 1021.040 287.990 ;
        RECT 1018.540 65.630 1018.800 65.950 ;
        RECT 1020.840 65.630 1021.100 65.950 ;
        RECT 1018.600 3.050 1018.740 65.630 ;
        RECT 1018.540 2.730 1018.800 3.050 ;
        RECT 1019.460 2.730 1019.720 3.050 ;
        RECT 1019.520 2.400 1019.660 2.730 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1121.165 283.305 1121.335 286.535 ;
      LAYER mcon ;
        RECT 1121.165 286.365 1121.335 286.535 ;
      LAYER met1 ;
        RECT 1151.910 286.860 1152.230 286.920 ;
        RECT 1142.800 286.720 1152.230 286.860 ;
        RECT 1121.105 286.520 1121.395 286.565 ;
        RECT 1142.800 286.520 1142.940 286.720 ;
        RECT 1151.910 286.660 1152.230 286.720 ;
        RECT 1121.105 286.380 1142.940 286.520 ;
        RECT 1121.105 286.335 1121.395 286.380 ;
        RECT 1041.510 283.460 1041.830 283.520 ;
        RECT 1121.105 283.460 1121.395 283.505 ;
        RECT 1041.510 283.320 1121.395 283.460 ;
        RECT 1041.510 283.260 1041.830 283.320 ;
        RECT 1121.105 283.275 1121.395 283.320 ;
        RECT 1037.370 20.640 1037.690 20.700 ;
        RECT 1041.510 20.640 1041.830 20.700 ;
        RECT 1037.370 20.500 1041.830 20.640 ;
        RECT 1037.370 20.440 1037.690 20.500 ;
        RECT 1041.510 20.440 1041.830 20.500 ;
      LAYER via ;
        RECT 1151.940 286.660 1152.200 286.920 ;
        RECT 1041.540 283.260 1041.800 283.520 ;
        RECT 1037.400 20.440 1037.660 20.700 ;
        RECT 1041.540 20.440 1041.800 20.700 ;
      LAYER met2 ;
        RECT 1151.940 300.000 1152.220 304.000 ;
        RECT 1152.000 286.950 1152.140 300.000 ;
        RECT 1151.940 286.630 1152.200 286.950 ;
        RECT 1041.540 283.230 1041.800 283.550 ;
        RECT 1041.600 20.730 1041.740 283.230 ;
        RECT 1037.400 20.410 1037.660 20.730 ;
        RECT 1041.540 20.410 1041.800 20.730 ;
        RECT 1037.460 2.400 1037.600 20.410 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1055.310 287.880 1055.630 287.940 ;
        RECT 1166.630 287.880 1166.950 287.940 ;
        RECT 1055.310 287.740 1166.950 287.880 ;
        RECT 1055.310 287.680 1055.630 287.740 ;
        RECT 1166.630 287.680 1166.950 287.740 ;
      LAYER via ;
        RECT 1055.340 287.680 1055.600 287.940 ;
        RECT 1166.660 287.680 1166.920 287.940 ;
      LAYER met2 ;
        RECT 1166.660 300.000 1166.940 304.000 ;
        RECT 1166.720 287.970 1166.860 300.000 ;
        RECT 1055.340 287.650 1055.600 287.970 ;
        RECT 1166.660 287.650 1166.920 287.970 ;
        RECT 1055.400 2.400 1055.540 287.650 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1076.010 289.240 1076.330 289.300 ;
        RECT 1181.350 289.240 1181.670 289.300 ;
        RECT 1076.010 289.100 1181.670 289.240 ;
        RECT 1076.010 289.040 1076.330 289.100 ;
        RECT 1181.350 289.040 1181.670 289.100 ;
        RECT 1073.250 20.640 1073.570 20.700 ;
        RECT 1076.010 20.640 1076.330 20.700 ;
        RECT 1073.250 20.500 1076.330 20.640 ;
        RECT 1073.250 20.440 1073.570 20.500 ;
        RECT 1076.010 20.440 1076.330 20.500 ;
      LAYER via ;
        RECT 1076.040 289.040 1076.300 289.300 ;
        RECT 1181.380 289.040 1181.640 289.300 ;
        RECT 1073.280 20.440 1073.540 20.700 ;
        RECT 1076.040 20.440 1076.300 20.700 ;
      LAYER met2 ;
        RECT 1181.380 300.000 1181.660 304.000 ;
        RECT 1181.440 289.330 1181.580 300.000 ;
        RECT 1076.040 289.010 1076.300 289.330 ;
        RECT 1181.380 289.010 1181.640 289.330 ;
        RECT 1076.100 20.730 1076.240 289.010 ;
        RECT 1073.280 20.410 1073.540 20.730 ;
        RECT 1076.040 20.410 1076.300 20.730 ;
        RECT 1073.340 2.400 1073.480 20.410 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.710 285.500 1097.030 285.560 ;
        RECT 1196.070 285.500 1196.390 285.560 ;
        RECT 1096.710 285.360 1196.390 285.500 ;
        RECT 1096.710 285.300 1097.030 285.360 ;
        RECT 1196.070 285.300 1196.390 285.360 ;
        RECT 1090.730 17.920 1091.050 17.980 ;
        RECT 1096.710 17.920 1097.030 17.980 ;
        RECT 1090.730 17.780 1097.030 17.920 ;
        RECT 1090.730 17.720 1091.050 17.780 ;
        RECT 1096.710 17.720 1097.030 17.780 ;
      LAYER via ;
        RECT 1096.740 285.300 1097.000 285.560 ;
        RECT 1196.100 285.300 1196.360 285.560 ;
        RECT 1090.760 17.720 1091.020 17.980 ;
        RECT 1096.740 17.720 1097.000 17.980 ;
      LAYER met2 ;
        RECT 1196.100 300.000 1196.380 304.000 ;
        RECT 1196.160 285.590 1196.300 300.000 ;
        RECT 1096.740 285.270 1097.000 285.590 ;
        RECT 1196.100 285.270 1196.360 285.590 ;
        RECT 1096.800 18.010 1096.940 285.270 ;
        RECT 1090.760 17.690 1091.020 18.010 ;
        RECT 1096.740 17.690 1097.000 18.010 ;
        RECT 1090.820 2.400 1090.960 17.690 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1120.705 288.745 1120.875 289.935 ;
      LAYER mcon ;
        RECT 1120.705 289.765 1120.875 289.935 ;
      LAYER met1 ;
        RECT 1120.645 289.920 1120.935 289.965 ;
        RECT 1120.645 289.780 1121.780 289.920 ;
        RECT 1120.645 289.735 1120.935 289.780 ;
        RECT 1121.640 289.580 1121.780 289.780 ;
        RECT 1210.790 289.580 1211.110 289.640 ;
        RECT 1121.640 289.440 1211.110 289.580 ;
        RECT 1210.790 289.380 1211.110 289.440 ;
        RECT 1110.510 288.900 1110.830 288.960 ;
        RECT 1120.645 288.900 1120.935 288.945 ;
        RECT 1110.510 288.760 1120.935 288.900 ;
        RECT 1110.510 288.700 1110.830 288.760 ;
        RECT 1120.645 288.715 1120.935 288.760 ;
      LAYER via ;
        RECT 1210.820 289.380 1211.080 289.640 ;
        RECT 1110.540 288.700 1110.800 288.960 ;
      LAYER met2 ;
        RECT 1210.820 300.000 1211.100 304.000 ;
        RECT 1210.880 289.670 1211.020 300.000 ;
        RECT 1210.820 289.350 1211.080 289.670 ;
        RECT 1110.540 288.670 1110.800 288.990 ;
        RECT 1110.600 17.410 1110.740 288.670 ;
        RECT 1108.760 17.270 1110.740 17.410 ;
        RECT 1108.760 2.400 1108.900 17.270 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1131.210 283.460 1131.530 283.520 ;
        RECT 1225.510 283.460 1225.830 283.520 ;
        RECT 1131.210 283.320 1225.830 283.460 ;
        RECT 1131.210 283.260 1131.530 283.320 ;
        RECT 1225.510 283.260 1225.830 283.320 ;
        RECT 1126.610 17.580 1126.930 17.640 ;
        RECT 1131.210 17.580 1131.530 17.640 ;
        RECT 1126.610 17.440 1131.530 17.580 ;
        RECT 1126.610 17.380 1126.930 17.440 ;
        RECT 1131.210 17.380 1131.530 17.440 ;
      LAYER via ;
        RECT 1131.240 283.260 1131.500 283.520 ;
        RECT 1225.540 283.260 1225.800 283.520 ;
        RECT 1126.640 17.380 1126.900 17.640 ;
        RECT 1131.240 17.380 1131.500 17.640 ;
      LAYER met2 ;
        RECT 1225.540 300.000 1225.820 304.000 ;
        RECT 1225.600 283.550 1225.740 300.000 ;
        RECT 1131.240 283.230 1131.500 283.550 ;
        RECT 1225.540 283.230 1225.800 283.550 ;
        RECT 1131.300 17.670 1131.440 283.230 ;
        RECT 1126.640 17.350 1126.900 17.670 ;
        RECT 1131.240 17.350 1131.500 17.670 ;
        RECT 1126.700 2.400 1126.840 17.350 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1144.550 286.520 1144.870 286.580 ;
        RECT 1240.230 286.520 1240.550 286.580 ;
        RECT 1144.550 286.380 1240.550 286.520 ;
        RECT 1144.550 286.320 1144.870 286.380 ;
        RECT 1240.230 286.320 1240.550 286.380 ;
      LAYER via ;
        RECT 1144.580 286.320 1144.840 286.580 ;
        RECT 1240.260 286.320 1240.520 286.580 ;
      LAYER met2 ;
        RECT 1240.260 300.000 1240.540 304.000 ;
        RECT 1240.320 286.610 1240.460 300.000 ;
        RECT 1144.580 286.290 1144.840 286.610 ;
        RECT 1240.260 286.290 1240.520 286.610 ;
        RECT 1144.640 2.400 1144.780 286.290 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1165.710 288.560 1166.030 288.620 ;
        RECT 1254.950 288.560 1255.270 288.620 ;
        RECT 1165.710 288.420 1255.270 288.560 ;
        RECT 1165.710 288.360 1166.030 288.420 ;
        RECT 1254.950 288.360 1255.270 288.420 ;
        RECT 1162.490 17.580 1162.810 17.640 ;
        RECT 1165.710 17.580 1166.030 17.640 ;
        RECT 1162.490 17.440 1166.030 17.580 ;
        RECT 1162.490 17.380 1162.810 17.440 ;
        RECT 1165.710 17.380 1166.030 17.440 ;
      LAYER via ;
        RECT 1165.740 288.360 1166.000 288.620 ;
        RECT 1254.980 288.360 1255.240 288.620 ;
        RECT 1162.520 17.380 1162.780 17.640 ;
        RECT 1165.740 17.380 1166.000 17.640 ;
      LAYER met2 ;
        RECT 1254.980 300.000 1255.260 304.000 ;
        RECT 1255.040 288.650 1255.180 300.000 ;
        RECT 1165.740 288.330 1166.000 288.650 ;
        RECT 1254.980 288.330 1255.240 288.650 ;
        RECT 1165.800 17.670 1165.940 288.330 ;
        RECT 1162.520 17.350 1162.780 17.670 ;
        RECT 1165.740 17.350 1166.000 17.670 ;
        RECT 1162.580 2.400 1162.720 17.350 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 682.710 287.200 683.030 287.260 ;
        RECT 682.710 287.060 714.220 287.200 ;
        RECT 682.710 287.000 683.030 287.060 ;
        RECT 714.080 286.860 714.220 287.060 ;
        RECT 857.970 286.860 858.290 286.920 ;
        RECT 714.080 286.720 858.290 286.860 ;
        RECT 857.970 286.660 858.290 286.720 ;
        RECT 680.410 20.640 680.730 20.700 ;
        RECT 682.710 20.640 683.030 20.700 ;
        RECT 680.410 20.500 683.030 20.640 ;
        RECT 680.410 20.440 680.730 20.500 ;
        RECT 682.710 20.440 683.030 20.500 ;
      LAYER via ;
        RECT 682.740 287.000 683.000 287.260 ;
        RECT 858.000 286.660 858.260 286.920 ;
        RECT 680.440 20.440 680.700 20.700 ;
        RECT 682.740 20.440 683.000 20.700 ;
      LAYER met2 ;
        RECT 858.000 300.000 858.280 304.000 ;
        RECT 682.740 286.970 683.000 287.290 ;
        RECT 682.800 20.730 682.940 286.970 ;
        RECT 858.060 286.950 858.200 300.000 ;
        RECT 858.000 286.630 858.260 286.950 ;
        RECT 680.440 20.410 680.700 20.730 ;
        RECT 682.740 20.410 683.000 20.730 ;
        RECT 680.500 2.400 680.640 20.410 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 288.900 1186.730 288.960 ;
        RECT 1269.670 288.900 1269.990 288.960 ;
        RECT 1186.410 288.760 1269.990 288.900 ;
        RECT 1186.410 288.700 1186.730 288.760 ;
        RECT 1269.670 288.700 1269.990 288.760 ;
        RECT 1179.970 16.220 1180.290 16.280 ;
        RECT 1186.410 16.220 1186.730 16.280 ;
        RECT 1179.970 16.080 1186.730 16.220 ;
        RECT 1179.970 16.020 1180.290 16.080 ;
        RECT 1186.410 16.020 1186.730 16.080 ;
      LAYER via ;
        RECT 1186.440 288.700 1186.700 288.960 ;
        RECT 1269.700 288.700 1269.960 288.960 ;
        RECT 1180.000 16.020 1180.260 16.280 ;
        RECT 1186.440 16.020 1186.700 16.280 ;
      LAYER met2 ;
        RECT 1269.700 300.000 1269.980 304.000 ;
        RECT 1269.760 288.990 1269.900 300.000 ;
        RECT 1186.440 288.670 1186.700 288.990 ;
        RECT 1269.700 288.670 1269.960 288.990 ;
        RECT 1186.500 16.310 1186.640 288.670 ;
        RECT 1180.000 15.990 1180.260 16.310 ;
        RECT 1186.440 15.990 1186.700 16.310 ;
        RECT 1180.060 2.400 1180.200 15.990 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1200.210 289.240 1200.530 289.300 ;
        RECT 1284.390 289.240 1284.710 289.300 ;
        RECT 1200.210 289.100 1284.710 289.240 ;
        RECT 1200.210 289.040 1200.530 289.100 ;
        RECT 1284.390 289.040 1284.710 289.100 ;
        RECT 1197.910 17.580 1198.230 17.640 ;
        RECT 1200.210 17.580 1200.530 17.640 ;
        RECT 1197.910 17.440 1200.530 17.580 ;
        RECT 1197.910 17.380 1198.230 17.440 ;
        RECT 1200.210 17.380 1200.530 17.440 ;
      LAYER via ;
        RECT 1200.240 289.040 1200.500 289.300 ;
        RECT 1284.420 289.040 1284.680 289.300 ;
        RECT 1197.940 17.380 1198.200 17.640 ;
        RECT 1200.240 17.380 1200.500 17.640 ;
      LAYER met2 ;
        RECT 1284.420 300.000 1284.700 304.000 ;
        RECT 1284.480 289.330 1284.620 300.000 ;
        RECT 1200.240 289.010 1200.500 289.330 ;
        RECT 1284.420 289.010 1284.680 289.330 ;
        RECT 1200.300 17.670 1200.440 289.010 ;
        RECT 1197.940 17.350 1198.200 17.670 ;
        RECT 1200.240 17.350 1200.500 17.670 ;
        RECT 1198.000 2.400 1198.140 17.350 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1220.910 286.180 1221.230 286.240 ;
        RECT 1298.650 286.180 1298.970 286.240 ;
        RECT 1220.910 286.040 1298.970 286.180 ;
        RECT 1220.910 285.980 1221.230 286.040 ;
        RECT 1298.650 285.980 1298.970 286.040 ;
        RECT 1215.850 17.580 1216.170 17.640 ;
        RECT 1220.910 17.580 1221.230 17.640 ;
        RECT 1215.850 17.440 1221.230 17.580 ;
        RECT 1215.850 17.380 1216.170 17.440 ;
        RECT 1220.910 17.380 1221.230 17.440 ;
      LAYER via ;
        RECT 1220.940 285.980 1221.200 286.240 ;
        RECT 1298.680 285.980 1298.940 286.240 ;
        RECT 1215.880 17.380 1216.140 17.640 ;
        RECT 1220.940 17.380 1221.200 17.640 ;
      LAYER met2 ;
        RECT 1298.680 300.000 1298.960 304.000 ;
        RECT 1298.740 286.270 1298.880 300.000 ;
        RECT 1220.940 285.950 1221.200 286.270 ;
        RECT 1298.680 285.950 1298.940 286.270 ;
        RECT 1221.000 17.670 1221.140 285.950 ;
        RECT 1215.880 17.350 1216.140 17.670 ;
        RECT 1220.940 17.350 1221.200 17.670 ;
        RECT 1215.940 2.400 1216.080 17.350 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1234.710 285.840 1235.030 285.900 ;
        RECT 1313.370 285.840 1313.690 285.900 ;
        RECT 1234.710 285.700 1313.690 285.840 ;
        RECT 1234.710 285.640 1235.030 285.700 ;
        RECT 1313.370 285.640 1313.690 285.700 ;
      LAYER via ;
        RECT 1234.740 285.640 1235.000 285.900 ;
        RECT 1313.400 285.640 1313.660 285.900 ;
      LAYER met2 ;
        RECT 1313.400 300.000 1313.680 304.000 ;
        RECT 1313.460 285.930 1313.600 300.000 ;
        RECT 1234.740 285.610 1235.000 285.930 ;
        RECT 1313.400 285.610 1313.660 285.930 ;
        RECT 1234.800 17.410 1234.940 285.610 ;
        RECT 1233.880 17.270 1234.940 17.410 ;
        RECT 1233.880 2.400 1234.020 17.270 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1255.410 287.200 1255.730 287.260 ;
        RECT 1328.090 287.200 1328.410 287.260 ;
        RECT 1255.410 287.060 1328.410 287.200 ;
        RECT 1255.410 287.000 1255.730 287.060 ;
        RECT 1328.090 287.000 1328.410 287.060 ;
        RECT 1251.730 17.580 1252.050 17.640 ;
        RECT 1255.410 17.580 1255.730 17.640 ;
        RECT 1251.730 17.440 1255.730 17.580 ;
        RECT 1251.730 17.380 1252.050 17.440 ;
        RECT 1255.410 17.380 1255.730 17.440 ;
      LAYER via ;
        RECT 1255.440 287.000 1255.700 287.260 ;
        RECT 1328.120 287.000 1328.380 287.260 ;
        RECT 1251.760 17.380 1252.020 17.640 ;
        RECT 1255.440 17.380 1255.700 17.640 ;
      LAYER met2 ;
        RECT 1328.120 300.000 1328.400 304.000 ;
        RECT 1328.180 287.290 1328.320 300.000 ;
        RECT 1255.440 286.970 1255.700 287.290 ;
        RECT 1328.120 286.970 1328.380 287.290 ;
        RECT 1255.500 17.670 1255.640 286.970 ;
        RECT 1251.760 17.350 1252.020 17.670 ;
        RECT 1255.440 17.350 1255.700 17.670 ;
        RECT 1251.820 2.400 1251.960 17.350 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1268.750 286.860 1269.070 286.920 ;
        RECT 1342.810 286.860 1343.130 286.920 ;
        RECT 1268.750 286.720 1343.130 286.860 ;
        RECT 1268.750 286.660 1269.070 286.720 ;
        RECT 1342.810 286.660 1343.130 286.720 ;
      LAYER via ;
        RECT 1268.780 286.660 1269.040 286.920 ;
        RECT 1342.840 286.660 1343.100 286.920 ;
      LAYER met2 ;
        RECT 1342.840 300.000 1343.120 304.000 ;
        RECT 1342.900 286.950 1343.040 300.000 ;
        RECT 1268.780 286.630 1269.040 286.950 ;
        RECT 1342.840 286.630 1343.100 286.950 ;
        RECT 1268.840 17.410 1268.980 286.630 ;
        RECT 1268.840 17.270 1269.440 17.410 ;
        RECT 1269.300 2.400 1269.440 17.270 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1289.910 288.900 1290.230 288.960 ;
        RECT 1357.530 288.900 1357.850 288.960 ;
        RECT 1289.910 288.760 1357.850 288.900 ;
        RECT 1289.910 288.700 1290.230 288.760 ;
        RECT 1357.530 288.700 1357.850 288.760 ;
        RECT 1287.150 17.580 1287.470 17.640 ;
        RECT 1289.910 17.580 1290.230 17.640 ;
        RECT 1287.150 17.440 1290.230 17.580 ;
        RECT 1287.150 17.380 1287.470 17.440 ;
        RECT 1289.910 17.380 1290.230 17.440 ;
      LAYER via ;
        RECT 1289.940 288.700 1290.200 288.960 ;
        RECT 1357.560 288.700 1357.820 288.960 ;
        RECT 1287.180 17.380 1287.440 17.640 ;
        RECT 1289.940 17.380 1290.200 17.640 ;
      LAYER met2 ;
        RECT 1357.560 300.000 1357.840 304.000 ;
        RECT 1357.620 288.990 1357.760 300.000 ;
        RECT 1289.940 288.670 1290.200 288.990 ;
        RECT 1357.560 288.670 1357.820 288.990 ;
        RECT 1290.000 17.670 1290.140 288.670 ;
        RECT 1287.180 17.350 1287.440 17.670 ;
        RECT 1289.940 17.350 1290.200 17.670 ;
        RECT 1287.240 2.400 1287.380 17.350 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1310.610 285.500 1310.930 285.560 ;
        RECT 1372.250 285.500 1372.570 285.560 ;
        RECT 1310.610 285.360 1372.570 285.500 ;
        RECT 1310.610 285.300 1310.930 285.360 ;
        RECT 1372.250 285.300 1372.570 285.360 ;
        RECT 1305.090 16.220 1305.410 16.280 ;
        RECT 1310.610 16.220 1310.930 16.280 ;
        RECT 1305.090 16.080 1310.930 16.220 ;
        RECT 1305.090 16.020 1305.410 16.080 ;
        RECT 1310.610 16.020 1310.930 16.080 ;
      LAYER via ;
        RECT 1310.640 285.300 1310.900 285.560 ;
        RECT 1372.280 285.300 1372.540 285.560 ;
        RECT 1305.120 16.020 1305.380 16.280 ;
        RECT 1310.640 16.020 1310.900 16.280 ;
      LAYER met2 ;
        RECT 1372.280 300.000 1372.560 304.000 ;
        RECT 1372.340 285.590 1372.480 300.000 ;
        RECT 1310.640 285.270 1310.900 285.590 ;
        RECT 1372.280 285.270 1372.540 285.590 ;
        RECT 1310.700 16.310 1310.840 285.270 ;
        RECT 1305.120 15.990 1305.380 16.310 ;
        RECT 1310.640 15.990 1310.900 16.310 ;
        RECT 1305.180 2.400 1305.320 15.990 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1324.410 286.520 1324.730 286.580 ;
        RECT 1386.970 286.520 1387.290 286.580 ;
        RECT 1324.410 286.380 1387.290 286.520 ;
        RECT 1324.410 286.320 1324.730 286.380 ;
        RECT 1386.970 286.320 1387.290 286.380 ;
      LAYER via ;
        RECT 1324.440 286.320 1324.700 286.580 ;
        RECT 1387.000 286.320 1387.260 286.580 ;
      LAYER met2 ;
        RECT 1387.000 300.000 1387.280 304.000 ;
        RECT 1387.060 286.610 1387.200 300.000 ;
        RECT 1324.440 286.290 1324.700 286.610 ;
        RECT 1387.000 286.290 1387.260 286.610 ;
        RECT 1324.500 17.410 1324.640 286.290 ;
        RECT 1323.120 17.270 1324.640 17.410 ;
        RECT 1323.120 2.400 1323.260 17.270 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1345.110 285.840 1345.430 285.900 ;
        RECT 1401.690 285.840 1402.010 285.900 ;
        RECT 1345.110 285.700 1402.010 285.840 ;
        RECT 1345.110 285.640 1345.430 285.700 ;
        RECT 1401.690 285.640 1402.010 285.700 ;
        RECT 1340.510 15.200 1340.830 15.260 ;
        RECT 1345.110 15.200 1345.430 15.260 ;
        RECT 1340.510 15.060 1345.430 15.200 ;
        RECT 1340.510 15.000 1340.830 15.060 ;
        RECT 1345.110 15.000 1345.430 15.060 ;
      LAYER via ;
        RECT 1345.140 285.640 1345.400 285.900 ;
        RECT 1401.720 285.640 1401.980 285.900 ;
        RECT 1340.540 15.000 1340.800 15.260 ;
        RECT 1345.140 15.000 1345.400 15.260 ;
      LAYER met2 ;
        RECT 1401.720 300.000 1402.000 304.000 ;
        RECT 1401.780 285.930 1401.920 300.000 ;
        RECT 1345.140 285.610 1345.400 285.930 ;
        RECT 1401.720 285.610 1401.980 285.930 ;
        RECT 1345.200 15.290 1345.340 285.610 ;
        RECT 1340.540 14.970 1340.800 15.290 ;
        RECT 1345.140 14.970 1345.400 15.290 ;
        RECT 1340.600 2.400 1340.740 14.970 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 703.410 288.220 703.730 288.280 ;
        RECT 703.410 288.080 736.300 288.220 ;
        RECT 703.410 288.020 703.730 288.080 ;
        RECT 736.160 287.200 736.300 288.080 ;
        RECT 872.690 287.200 873.010 287.260 ;
        RECT 736.160 287.060 873.010 287.200 ;
        RECT 872.690 287.000 873.010 287.060 ;
        RECT 698.350 14.860 698.670 14.920 ;
        RECT 703.410 14.860 703.730 14.920 ;
        RECT 698.350 14.720 703.730 14.860 ;
        RECT 698.350 14.660 698.670 14.720 ;
        RECT 703.410 14.660 703.730 14.720 ;
      LAYER via ;
        RECT 703.440 288.020 703.700 288.280 ;
        RECT 872.720 287.000 872.980 287.260 ;
        RECT 698.380 14.660 698.640 14.920 ;
        RECT 703.440 14.660 703.700 14.920 ;
      LAYER met2 ;
        RECT 872.720 300.000 873.000 304.000 ;
        RECT 703.440 287.990 703.700 288.310 ;
        RECT 703.500 14.950 703.640 287.990 ;
        RECT 872.780 287.290 872.920 300.000 ;
        RECT 872.720 286.970 872.980 287.290 ;
        RECT 698.380 14.630 698.640 14.950 ;
        RECT 703.440 14.630 703.700 14.950 ;
        RECT 698.440 2.400 698.580 14.630 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1358.910 286.860 1359.230 286.920 ;
        RECT 1416.410 286.860 1416.730 286.920 ;
        RECT 1358.910 286.720 1416.730 286.860 ;
        RECT 1358.910 286.660 1359.230 286.720 ;
        RECT 1416.410 286.660 1416.730 286.720 ;
      LAYER via ;
        RECT 1358.940 286.660 1359.200 286.920 ;
        RECT 1416.440 286.660 1416.700 286.920 ;
      LAYER met2 ;
        RECT 1416.440 300.000 1416.720 304.000 ;
        RECT 1416.500 286.950 1416.640 300.000 ;
        RECT 1358.940 286.630 1359.200 286.950 ;
        RECT 1416.440 286.630 1416.700 286.950 ;
        RECT 1359.000 17.410 1359.140 286.630 ;
        RECT 1358.540 17.270 1359.140 17.410 ;
        RECT 1358.540 2.400 1358.680 17.270 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1379.610 288.900 1379.930 288.960 ;
        RECT 1431.130 288.900 1431.450 288.960 ;
        RECT 1379.610 288.760 1431.450 288.900 ;
        RECT 1379.610 288.700 1379.930 288.760 ;
        RECT 1431.130 288.700 1431.450 288.760 ;
        RECT 1376.390 17.580 1376.710 17.640 ;
        RECT 1379.610 17.580 1379.930 17.640 ;
        RECT 1376.390 17.440 1379.930 17.580 ;
        RECT 1376.390 17.380 1376.710 17.440 ;
        RECT 1379.610 17.380 1379.930 17.440 ;
      LAYER via ;
        RECT 1379.640 288.700 1379.900 288.960 ;
        RECT 1431.160 288.700 1431.420 288.960 ;
        RECT 1376.420 17.380 1376.680 17.640 ;
        RECT 1379.640 17.380 1379.900 17.640 ;
      LAYER met2 ;
        RECT 1431.160 300.000 1431.440 304.000 ;
        RECT 1431.220 288.990 1431.360 300.000 ;
        RECT 1379.640 288.670 1379.900 288.990 ;
        RECT 1431.160 288.670 1431.420 288.990 ;
        RECT 1379.700 17.670 1379.840 288.670 ;
        RECT 1376.420 17.350 1376.680 17.670 ;
        RECT 1379.640 17.350 1379.900 17.670 ;
        RECT 1376.480 2.400 1376.620 17.350 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.310 289.580 1400.630 289.640 ;
        RECT 1445.850 289.580 1446.170 289.640 ;
        RECT 1400.310 289.440 1446.170 289.580 ;
        RECT 1400.310 289.380 1400.630 289.440 ;
        RECT 1445.850 289.380 1446.170 289.440 ;
        RECT 1394.330 17.920 1394.650 17.980 ;
        RECT 1400.310 17.920 1400.630 17.980 ;
        RECT 1394.330 17.780 1400.630 17.920 ;
        RECT 1394.330 17.720 1394.650 17.780 ;
        RECT 1400.310 17.720 1400.630 17.780 ;
      LAYER via ;
        RECT 1400.340 289.380 1400.600 289.640 ;
        RECT 1445.880 289.380 1446.140 289.640 ;
        RECT 1394.360 17.720 1394.620 17.980 ;
        RECT 1400.340 17.720 1400.600 17.980 ;
      LAYER met2 ;
        RECT 1445.880 300.000 1446.160 304.000 ;
        RECT 1445.940 289.670 1446.080 300.000 ;
        RECT 1400.340 289.350 1400.600 289.670 ;
        RECT 1445.880 289.350 1446.140 289.670 ;
        RECT 1400.400 18.010 1400.540 289.350 ;
        RECT 1394.360 17.690 1394.620 18.010 ;
        RECT 1400.340 17.690 1400.600 18.010 ;
        RECT 1394.420 2.400 1394.560 17.690 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1414.110 287.200 1414.430 287.260 ;
        RECT 1460.570 287.200 1460.890 287.260 ;
        RECT 1414.110 287.060 1460.890 287.200 ;
        RECT 1414.110 287.000 1414.430 287.060 ;
        RECT 1460.570 287.000 1460.890 287.060 ;
      LAYER via ;
        RECT 1414.140 287.000 1414.400 287.260 ;
        RECT 1460.600 287.000 1460.860 287.260 ;
      LAYER met2 ;
        RECT 1460.600 300.000 1460.880 304.000 ;
        RECT 1460.660 287.290 1460.800 300.000 ;
        RECT 1414.140 286.970 1414.400 287.290 ;
        RECT 1460.600 286.970 1460.860 287.290 ;
        RECT 1414.200 17.580 1414.340 286.970 ;
        RECT 1412.360 17.440 1414.340 17.580 ;
        RECT 1412.360 2.400 1412.500 17.440 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1434.810 287.880 1435.130 287.940 ;
        RECT 1475.290 287.880 1475.610 287.940 ;
        RECT 1434.810 287.740 1475.610 287.880 ;
        RECT 1434.810 287.680 1435.130 287.740 ;
        RECT 1475.290 287.680 1475.610 287.740 ;
        RECT 1429.750 17.580 1430.070 17.640 ;
        RECT 1434.810 17.580 1435.130 17.640 ;
        RECT 1429.750 17.440 1435.130 17.580 ;
        RECT 1429.750 17.380 1430.070 17.440 ;
        RECT 1434.810 17.380 1435.130 17.440 ;
      LAYER via ;
        RECT 1434.840 287.680 1435.100 287.940 ;
        RECT 1475.320 287.680 1475.580 287.940 ;
        RECT 1429.780 17.380 1430.040 17.640 ;
        RECT 1434.840 17.380 1435.100 17.640 ;
      LAYER met2 ;
        RECT 1475.320 300.000 1475.600 304.000 ;
        RECT 1475.380 287.970 1475.520 300.000 ;
        RECT 1434.840 287.650 1435.100 287.970 ;
        RECT 1475.320 287.650 1475.580 287.970 ;
        RECT 1434.900 17.670 1435.040 287.650 ;
        RECT 1429.780 17.350 1430.040 17.670 ;
        RECT 1434.840 17.350 1435.100 17.670 ;
        RECT 1429.840 2.400 1429.980 17.350 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1448.610 287.540 1448.930 287.600 ;
        RECT 1490.010 287.540 1490.330 287.600 ;
        RECT 1448.610 287.400 1490.330 287.540 ;
        RECT 1448.610 287.340 1448.930 287.400 ;
        RECT 1490.010 287.340 1490.330 287.400 ;
      LAYER via ;
        RECT 1448.640 287.340 1448.900 287.600 ;
        RECT 1490.040 287.340 1490.300 287.600 ;
      LAYER met2 ;
        RECT 1490.040 300.000 1490.320 304.000 ;
        RECT 1490.100 287.630 1490.240 300.000 ;
        RECT 1448.640 287.310 1448.900 287.630 ;
        RECT 1490.040 287.310 1490.300 287.630 ;
        RECT 1448.700 17.410 1448.840 287.310 ;
        RECT 1447.780 17.270 1448.840 17.410 ;
        RECT 1447.780 2.400 1447.920 17.270 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1469.310 286.180 1469.630 286.240 ;
        RECT 1504.730 286.180 1505.050 286.240 ;
        RECT 1469.310 286.040 1505.050 286.180 ;
        RECT 1469.310 285.980 1469.630 286.040 ;
        RECT 1504.730 285.980 1505.050 286.040 ;
        RECT 1465.630 17.580 1465.950 17.640 ;
        RECT 1469.310 17.580 1469.630 17.640 ;
        RECT 1465.630 17.440 1469.630 17.580 ;
        RECT 1465.630 17.380 1465.950 17.440 ;
        RECT 1469.310 17.380 1469.630 17.440 ;
      LAYER via ;
        RECT 1469.340 285.980 1469.600 286.240 ;
        RECT 1504.760 285.980 1505.020 286.240 ;
        RECT 1465.660 17.380 1465.920 17.640 ;
        RECT 1469.340 17.380 1469.600 17.640 ;
      LAYER met2 ;
        RECT 1504.760 300.000 1505.040 304.000 ;
        RECT 1504.820 286.270 1504.960 300.000 ;
        RECT 1469.340 285.950 1469.600 286.270 ;
        RECT 1504.760 285.950 1505.020 286.270 ;
        RECT 1469.400 17.670 1469.540 285.950 ;
        RECT 1465.660 17.350 1465.920 17.670 ;
        RECT 1469.340 17.350 1469.600 17.670 ;
        RECT 1465.720 2.400 1465.860 17.350 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1489.550 285.500 1489.870 285.560 ;
        RECT 1519.450 285.500 1519.770 285.560 ;
        RECT 1489.550 285.360 1519.770 285.500 ;
        RECT 1489.550 285.300 1489.870 285.360 ;
        RECT 1519.450 285.300 1519.770 285.360 ;
        RECT 1483.570 17.920 1483.890 17.980 ;
        RECT 1489.550 17.920 1489.870 17.980 ;
        RECT 1483.570 17.780 1489.870 17.920 ;
        RECT 1483.570 17.720 1483.890 17.780 ;
        RECT 1489.550 17.720 1489.870 17.780 ;
      LAYER via ;
        RECT 1489.580 285.300 1489.840 285.560 ;
        RECT 1519.480 285.300 1519.740 285.560 ;
        RECT 1483.600 17.720 1483.860 17.980 ;
        RECT 1489.580 17.720 1489.840 17.980 ;
      LAYER met2 ;
        RECT 1519.480 300.000 1519.760 304.000 ;
        RECT 1519.540 285.590 1519.680 300.000 ;
        RECT 1489.580 285.270 1489.840 285.590 ;
        RECT 1519.480 285.270 1519.740 285.590 ;
        RECT 1489.640 18.010 1489.780 285.270 ;
        RECT 1483.600 17.690 1483.860 18.010 ;
        RECT 1489.580 17.690 1489.840 18.010 ;
        RECT 1483.660 2.400 1483.800 17.690 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1521.290 283.120 1521.610 283.180 ;
        RECT 1534.170 283.120 1534.490 283.180 ;
        RECT 1521.290 282.980 1534.490 283.120 ;
        RECT 1521.290 282.920 1521.610 282.980 ;
        RECT 1534.170 282.920 1534.490 282.980 ;
        RECT 1501.510 16.560 1501.830 16.620 ;
        RECT 1521.290 16.560 1521.610 16.620 ;
        RECT 1501.510 16.420 1521.610 16.560 ;
        RECT 1501.510 16.360 1501.830 16.420 ;
        RECT 1521.290 16.360 1521.610 16.420 ;
      LAYER via ;
        RECT 1521.320 282.920 1521.580 283.180 ;
        RECT 1534.200 282.920 1534.460 283.180 ;
        RECT 1501.540 16.360 1501.800 16.620 ;
        RECT 1521.320 16.360 1521.580 16.620 ;
      LAYER met2 ;
        RECT 1534.200 300.000 1534.480 304.000 ;
        RECT 1534.260 283.210 1534.400 300.000 ;
        RECT 1521.320 282.890 1521.580 283.210 ;
        RECT 1534.200 282.890 1534.460 283.210 ;
        RECT 1521.380 16.650 1521.520 282.890 ;
        RECT 1501.540 16.330 1501.800 16.650 ;
        RECT 1521.320 16.330 1521.580 16.650 ;
        RECT 1501.600 2.400 1501.740 16.330 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.510 286.860 1524.830 286.920 ;
        RECT 1548.430 286.860 1548.750 286.920 ;
        RECT 1524.510 286.720 1548.750 286.860 ;
        RECT 1524.510 286.660 1524.830 286.720 ;
        RECT 1548.430 286.660 1548.750 286.720 ;
        RECT 1518.990 17.580 1519.310 17.640 ;
        RECT 1524.510 17.580 1524.830 17.640 ;
        RECT 1518.990 17.440 1524.830 17.580 ;
        RECT 1518.990 17.380 1519.310 17.440 ;
        RECT 1524.510 17.380 1524.830 17.440 ;
      LAYER via ;
        RECT 1524.540 286.660 1524.800 286.920 ;
        RECT 1548.460 286.660 1548.720 286.920 ;
        RECT 1519.020 17.380 1519.280 17.640 ;
        RECT 1524.540 17.380 1524.800 17.640 ;
      LAYER met2 ;
        RECT 1548.460 300.000 1548.740 304.000 ;
        RECT 1548.520 286.950 1548.660 300.000 ;
        RECT 1524.540 286.630 1524.800 286.950 ;
        RECT 1548.460 286.630 1548.720 286.950 ;
        RECT 1524.600 17.670 1524.740 286.630 ;
        RECT 1519.020 17.350 1519.280 17.670 ;
        RECT 1524.540 17.350 1524.800 17.670 ;
        RECT 1519.080 2.400 1519.220 17.350 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 738.445 283.985 738.615 287.555 ;
        RECT 716.365 2.805 716.535 14.195 ;
      LAYER mcon ;
        RECT 738.445 287.385 738.615 287.555 ;
        RECT 716.365 14.025 716.535 14.195 ;
      LAYER met1 ;
        RECT 738.385 287.540 738.675 287.585 ;
        RECT 887.410 287.540 887.730 287.600 ;
        RECT 738.385 287.400 887.730 287.540 ;
        RECT 738.385 287.355 738.675 287.400 ;
        RECT 887.410 287.340 887.730 287.400 ;
        RECT 717.210 284.140 717.530 284.200 ;
        RECT 738.385 284.140 738.675 284.185 ;
        RECT 717.210 284.000 738.675 284.140 ;
        RECT 717.210 283.940 717.530 284.000 ;
        RECT 738.385 283.955 738.675 284.000 ;
        RECT 716.305 14.180 716.595 14.225 ;
        RECT 717.210 14.180 717.530 14.240 ;
        RECT 716.305 14.040 717.530 14.180 ;
        RECT 716.305 13.995 716.595 14.040 ;
        RECT 717.210 13.980 717.530 14.040 ;
        RECT 716.290 2.960 716.610 3.020 ;
        RECT 716.095 2.820 716.610 2.960 ;
        RECT 716.290 2.760 716.610 2.820 ;
      LAYER via ;
        RECT 887.440 287.340 887.700 287.600 ;
        RECT 717.240 283.940 717.500 284.200 ;
        RECT 717.240 13.980 717.500 14.240 ;
        RECT 716.320 2.760 716.580 3.020 ;
      LAYER met2 ;
        RECT 887.440 300.000 887.720 304.000 ;
        RECT 887.500 287.630 887.640 300.000 ;
        RECT 887.440 287.310 887.700 287.630 ;
        RECT 717.240 283.910 717.500 284.230 ;
        RECT 717.300 14.270 717.440 283.910 ;
        RECT 717.240 13.950 717.500 14.270 ;
        RECT 716.320 2.730 716.580 3.050 ;
        RECT 716.380 2.400 716.520 2.730 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1538.310 284.480 1538.630 284.540 ;
        RECT 1563.150 284.480 1563.470 284.540 ;
        RECT 1538.310 284.340 1563.470 284.480 ;
        RECT 1538.310 284.280 1538.630 284.340 ;
        RECT 1563.150 284.280 1563.470 284.340 ;
      LAYER via ;
        RECT 1538.340 284.280 1538.600 284.540 ;
        RECT 1563.180 284.280 1563.440 284.540 ;
      LAYER met2 ;
        RECT 1563.180 300.000 1563.460 304.000 ;
        RECT 1563.240 284.570 1563.380 300.000 ;
        RECT 1538.340 284.250 1538.600 284.570 ;
        RECT 1563.180 284.250 1563.440 284.570 ;
        RECT 1538.400 17.410 1538.540 284.250 ;
        RECT 1537.020 17.270 1538.540 17.410 ;
        RECT 1537.020 2.400 1537.160 17.270 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1559.010 288.220 1559.330 288.280 ;
        RECT 1577.870 288.220 1578.190 288.280 ;
        RECT 1559.010 288.080 1578.190 288.220 ;
        RECT 1559.010 288.020 1559.330 288.080 ;
        RECT 1577.870 288.020 1578.190 288.080 ;
        RECT 1554.870 17.580 1555.190 17.640 ;
        RECT 1559.010 17.580 1559.330 17.640 ;
        RECT 1554.870 17.440 1559.330 17.580 ;
        RECT 1554.870 17.380 1555.190 17.440 ;
        RECT 1559.010 17.380 1559.330 17.440 ;
      LAYER via ;
        RECT 1559.040 288.020 1559.300 288.280 ;
        RECT 1577.900 288.020 1578.160 288.280 ;
        RECT 1554.900 17.380 1555.160 17.640 ;
        RECT 1559.040 17.380 1559.300 17.640 ;
      LAYER met2 ;
        RECT 1577.900 300.000 1578.180 304.000 ;
        RECT 1577.960 288.310 1578.100 300.000 ;
        RECT 1559.040 287.990 1559.300 288.310 ;
        RECT 1577.900 287.990 1578.160 288.310 ;
        RECT 1559.100 17.670 1559.240 287.990 ;
        RECT 1554.900 17.350 1555.160 17.670 ;
        RECT 1559.040 17.350 1559.300 17.670 ;
        RECT 1554.960 2.400 1555.100 17.350 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1576.490 283.460 1576.810 283.520 ;
        RECT 1592.590 283.460 1592.910 283.520 ;
        RECT 1576.490 283.320 1592.910 283.460 ;
        RECT 1576.490 283.260 1576.810 283.320 ;
        RECT 1592.590 283.260 1592.910 283.320 ;
        RECT 1572.810 17.580 1573.130 17.640 ;
        RECT 1576.490 17.580 1576.810 17.640 ;
        RECT 1572.810 17.440 1576.810 17.580 ;
        RECT 1572.810 17.380 1573.130 17.440 ;
        RECT 1576.490 17.380 1576.810 17.440 ;
      LAYER via ;
        RECT 1576.520 283.260 1576.780 283.520 ;
        RECT 1592.620 283.260 1592.880 283.520 ;
        RECT 1572.840 17.380 1573.100 17.640 ;
        RECT 1576.520 17.380 1576.780 17.640 ;
      LAYER met2 ;
        RECT 1592.620 300.000 1592.900 304.000 ;
        RECT 1592.680 283.550 1592.820 300.000 ;
        RECT 1576.520 283.230 1576.780 283.550 ;
        RECT 1592.620 283.230 1592.880 283.550 ;
        RECT 1576.580 17.670 1576.720 283.230 ;
        RECT 1572.840 17.350 1573.100 17.670 ;
        RECT 1576.520 17.350 1576.780 17.670 ;
        RECT 1572.900 2.400 1573.040 17.350 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1597.190 289.240 1597.510 289.300 ;
        RECT 1607.310 289.240 1607.630 289.300 ;
        RECT 1597.190 289.100 1607.630 289.240 ;
        RECT 1597.190 289.040 1597.510 289.100 ;
        RECT 1607.310 289.040 1607.630 289.100 ;
        RECT 1590.290 17.580 1590.610 17.640 ;
        RECT 1597.190 17.580 1597.510 17.640 ;
        RECT 1590.290 17.440 1597.510 17.580 ;
        RECT 1590.290 17.380 1590.610 17.440 ;
        RECT 1597.190 17.380 1597.510 17.440 ;
      LAYER via ;
        RECT 1597.220 289.040 1597.480 289.300 ;
        RECT 1607.340 289.040 1607.600 289.300 ;
        RECT 1590.320 17.380 1590.580 17.640 ;
        RECT 1597.220 17.380 1597.480 17.640 ;
      LAYER met2 ;
        RECT 1607.340 300.000 1607.620 304.000 ;
        RECT 1607.400 289.330 1607.540 300.000 ;
        RECT 1597.220 289.010 1597.480 289.330 ;
        RECT 1607.340 289.010 1607.600 289.330 ;
        RECT 1597.280 17.670 1597.420 289.010 ;
        RECT 1590.320 17.350 1590.580 17.670 ;
        RECT 1597.220 17.350 1597.480 17.670 ;
        RECT 1590.380 2.400 1590.520 17.350 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1613.750 287.880 1614.070 287.940 ;
        RECT 1622.030 287.880 1622.350 287.940 ;
        RECT 1613.750 287.740 1622.350 287.880 ;
        RECT 1613.750 287.680 1614.070 287.740 ;
        RECT 1622.030 287.680 1622.350 287.740 ;
        RECT 1608.230 17.580 1608.550 17.640 ;
        RECT 1613.750 17.580 1614.070 17.640 ;
        RECT 1608.230 17.440 1614.070 17.580 ;
        RECT 1608.230 17.380 1608.550 17.440 ;
        RECT 1613.750 17.380 1614.070 17.440 ;
      LAYER via ;
        RECT 1613.780 287.680 1614.040 287.940 ;
        RECT 1622.060 287.680 1622.320 287.940 ;
        RECT 1608.260 17.380 1608.520 17.640 ;
        RECT 1613.780 17.380 1614.040 17.640 ;
      LAYER met2 ;
        RECT 1622.060 300.000 1622.340 304.000 ;
        RECT 1622.120 287.970 1622.260 300.000 ;
        RECT 1613.780 287.650 1614.040 287.970 ;
        RECT 1622.060 287.650 1622.320 287.970 ;
        RECT 1613.840 17.670 1613.980 287.650 ;
        RECT 1608.260 17.350 1608.520 17.670 ;
        RECT 1613.780 17.350 1614.040 17.670 ;
        RECT 1608.320 2.400 1608.460 17.350 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1636.750 283.120 1637.070 283.180 ;
        RECT 1631.780 282.980 1637.070 283.120 ;
        RECT 1631.780 282.840 1631.920 282.980 ;
        RECT 1636.750 282.920 1637.070 282.980 ;
        RECT 1631.690 282.580 1632.010 282.840 ;
        RECT 1626.170 16.900 1626.490 16.960 ;
        RECT 1631.690 16.900 1632.010 16.960 ;
        RECT 1626.170 16.760 1632.010 16.900 ;
        RECT 1626.170 16.700 1626.490 16.760 ;
        RECT 1631.690 16.700 1632.010 16.760 ;
      LAYER via ;
        RECT 1636.780 282.920 1637.040 283.180 ;
        RECT 1631.720 282.580 1631.980 282.840 ;
        RECT 1626.200 16.700 1626.460 16.960 ;
        RECT 1631.720 16.700 1631.980 16.960 ;
      LAYER met2 ;
        RECT 1636.780 300.000 1637.060 304.000 ;
        RECT 1636.840 283.210 1636.980 300.000 ;
        RECT 1636.780 282.890 1637.040 283.210 ;
        RECT 1631.720 282.550 1631.980 282.870 ;
        RECT 1631.780 16.990 1631.920 282.550 ;
        RECT 1626.200 16.670 1626.460 16.990 ;
        RECT 1631.720 16.670 1631.980 16.990 ;
        RECT 1626.260 2.400 1626.400 16.670 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1644.110 17.580 1644.430 17.640 ;
        RECT 1649.630 17.580 1649.950 17.640 ;
        RECT 1644.110 17.440 1649.950 17.580 ;
        RECT 1644.110 17.380 1644.430 17.440 ;
        RECT 1649.630 17.380 1649.950 17.440 ;
      LAYER via ;
        RECT 1644.140 17.380 1644.400 17.640 ;
        RECT 1649.660 17.380 1649.920 17.640 ;
      LAYER met2 ;
        RECT 1651.500 300.290 1651.780 304.000 ;
        RECT 1649.720 300.150 1651.780 300.290 ;
        RECT 1649.720 17.670 1649.860 300.150 ;
        RECT 1651.500 300.000 1651.780 300.150 ;
        RECT 1644.140 17.350 1644.400 17.670 ;
        RECT 1649.660 17.350 1649.920 17.670 ;
        RECT 1644.200 2.400 1644.340 17.350 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1662.050 20.640 1662.370 20.700 ;
        RECT 1663.430 20.640 1663.750 20.700 ;
        RECT 1662.050 20.500 1663.750 20.640 ;
        RECT 1662.050 20.440 1662.370 20.500 ;
        RECT 1663.430 20.440 1663.750 20.500 ;
      LAYER via ;
        RECT 1662.080 20.440 1662.340 20.700 ;
        RECT 1663.460 20.440 1663.720 20.700 ;
      LAYER met2 ;
        RECT 1666.220 300.290 1666.500 304.000 ;
        RECT 1663.520 300.150 1666.500 300.290 ;
        RECT 1663.520 20.730 1663.660 300.150 ;
        RECT 1666.220 300.000 1666.500 300.150 ;
        RECT 1662.080 20.410 1662.340 20.730 ;
        RECT 1663.460 20.410 1663.720 20.730 ;
        RECT 1662.140 2.400 1662.280 20.410 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1676.770 20.640 1677.090 20.700 ;
        RECT 1679.530 20.640 1679.850 20.700 ;
        RECT 1676.770 20.500 1679.850 20.640 ;
        RECT 1676.770 20.440 1677.090 20.500 ;
        RECT 1679.530 20.440 1679.850 20.500 ;
      LAYER via ;
        RECT 1676.800 20.440 1677.060 20.700 ;
        RECT 1679.560 20.440 1679.820 20.700 ;
      LAYER met2 ;
        RECT 1680.940 300.290 1681.220 304.000 ;
        RECT 1676.860 300.150 1681.220 300.290 ;
        RECT 1676.860 20.730 1677.000 300.150 ;
        RECT 1680.940 300.000 1681.220 300.150 ;
        RECT 1676.800 20.410 1677.060 20.730 ;
        RECT 1679.560 20.410 1679.820 20.730 ;
        RECT 1679.620 2.400 1679.760 20.410 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1695.660 300.290 1695.940 304.000 ;
        RECT 1695.660 300.150 1697.240 300.290 ;
        RECT 1695.660 300.000 1695.940 300.150 ;
        RECT 1697.100 20.130 1697.240 300.150 ;
        RECT 1697.100 19.990 1697.700 20.130 ;
        RECT 1697.560 2.400 1697.700 19.990 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 737.910 288.560 738.230 288.620 ;
        RECT 902.130 288.560 902.450 288.620 ;
        RECT 737.910 288.420 902.450 288.560 ;
        RECT 737.910 288.360 738.230 288.420 ;
        RECT 902.130 288.360 902.450 288.420 ;
        RECT 734.230 16.900 734.550 16.960 ;
        RECT 737.910 16.900 738.230 16.960 ;
        RECT 734.230 16.760 738.230 16.900 ;
        RECT 734.230 16.700 734.550 16.760 ;
        RECT 737.910 16.700 738.230 16.760 ;
      LAYER via ;
        RECT 737.940 288.360 738.200 288.620 ;
        RECT 902.160 288.360 902.420 288.620 ;
        RECT 734.260 16.700 734.520 16.960 ;
        RECT 737.940 16.700 738.200 16.960 ;
      LAYER met2 ;
        RECT 902.160 300.000 902.440 304.000 ;
        RECT 902.220 288.650 902.360 300.000 ;
        RECT 737.940 288.330 738.200 288.650 ;
        RECT 902.160 288.330 902.420 288.650 ;
        RECT 738.000 16.990 738.140 288.330 ;
        RECT 734.260 16.670 734.520 16.990 ;
        RECT 737.940 16.670 738.200 16.990 ;
        RECT 734.320 2.400 734.460 16.670 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1710.810 17.580 1711.130 17.640 ;
        RECT 1715.410 17.580 1715.730 17.640 ;
        RECT 1710.810 17.440 1715.730 17.580 ;
        RECT 1710.810 17.380 1711.130 17.440 ;
        RECT 1715.410 17.380 1715.730 17.440 ;
      LAYER via ;
        RECT 1710.840 17.380 1711.100 17.640 ;
        RECT 1715.440 17.380 1715.700 17.640 ;
      LAYER met2 ;
        RECT 1710.380 300.290 1710.660 304.000 ;
        RECT 1710.380 300.150 1711.040 300.290 ;
        RECT 1710.380 300.000 1710.660 300.150 ;
        RECT 1710.900 17.670 1711.040 300.150 ;
        RECT 1710.840 17.350 1711.100 17.670 ;
        RECT 1715.440 17.350 1715.700 17.670 ;
        RECT 1715.500 2.400 1715.640 17.350 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1725.070 284.820 1725.390 284.880 ;
        RECT 1731.510 284.820 1731.830 284.880 ;
        RECT 1725.070 284.680 1731.830 284.820 ;
        RECT 1725.070 284.620 1725.390 284.680 ;
        RECT 1731.510 284.620 1731.830 284.680 ;
      LAYER via ;
        RECT 1725.100 284.620 1725.360 284.880 ;
        RECT 1731.540 284.620 1731.800 284.880 ;
      LAYER met2 ;
        RECT 1725.100 300.000 1725.380 304.000 ;
        RECT 1725.160 284.910 1725.300 300.000 ;
        RECT 1725.100 284.590 1725.360 284.910 ;
        RECT 1731.540 284.590 1731.800 284.910 ;
        RECT 1731.600 17.410 1731.740 284.590 ;
        RECT 1731.600 17.270 1733.580 17.410 ;
        RECT 1733.440 2.400 1733.580 17.270 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1739.790 288.900 1740.110 288.960 ;
        RECT 1745.310 288.900 1745.630 288.960 ;
        RECT 1739.790 288.760 1745.630 288.900 ;
        RECT 1739.790 288.700 1740.110 288.760 ;
        RECT 1745.310 288.700 1745.630 288.760 ;
        RECT 1745.310 17.580 1745.630 17.640 ;
        RECT 1751.290 17.580 1751.610 17.640 ;
        RECT 1745.310 17.440 1751.610 17.580 ;
        RECT 1745.310 17.380 1745.630 17.440 ;
        RECT 1751.290 17.380 1751.610 17.440 ;
      LAYER via ;
        RECT 1739.820 288.700 1740.080 288.960 ;
        RECT 1745.340 288.700 1745.600 288.960 ;
        RECT 1745.340 17.380 1745.600 17.640 ;
        RECT 1751.320 17.380 1751.580 17.640 ;
      LAYER met2 ;
        RECT 1739.820 300.000 1740.100 304.000 ;
        RECT 1739.880 288.990 1740.020 300.000 ;
        RECT 1739.820 288.670 1740.080 288.990 ;
        RECT 1745.340 288.670 1745.600 288.990 ;
        RECT 1745.400 17.670 1745.540 288.670 ;
        RECT 1745.340 17.350 1745.600 17.670 ;
        RECT 1751.320 17.350 1751.580 17.670 ;
        RECT 1751.380 2.400 1751.520 17.350 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1754.510 288.220 1754.830 288.280 ;
        RECT 1759.110 288.220 1759.430 288.280 ;
        RECT 1754.510 288.080 1759.430 288.220 ;
        RECT 1754.510 288.020 1754.830 288.080 ;
        RECT 1759.110 288.020 1759.430 288.080 ;
        RECT 1759.110 15.200 1759.430 15.260 ;
        RECT 1768.770 15.200 1769.090 15.260 ;
        RECT 1759.110 15.060 1769.090 15.200 ;
        RECT 1759.110 15.000 1759.430 15.060 ;
        RECT 1768.770 15.000 1769.090 15.060 ;
      LAYER via ;
        RECT 1754.540 288.020 1754.800 288.280 ;
        RECT 1759.140 288.020 1759.400 288.280 ;
        RECT 1759.140 15.000 1759.400 15.260 ;
        RECT 1768.800 15.000 1769.060 15.260 ;
      LAYER met2 ;
        RECT 1754.540 300.000 1754.820 304.000 ;
        RECT 1754.600 288.310 1754.740 300.000 ;
        RECT 1754.540 287.990 1754.800 288.310 ;
        RECT 1759.140 287.990 1759.400 288.310 ;
        RECT 1759.200 15.290 1759.340 287.990 ;
        RECT 1759.140 14.970 1759.400 15.290 ;
        RECT 1768.800 14.970 1769.060 15.290 ;
        RECT 1768.860 2.400 1769.000 14.970 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1769.230 285.500 1769.550 285.560 ;
        RECT 1780.730 285.500 1781.050 285.560 ;
        RECT 1769.230 285.360 1781.050 285.500 ;
        RECT 1769.230 285.300 1769.550 285.360 ;
        RECT 1780.730 285.300 1781.050 285.360 ;
        RECT 1780.730 21.320 1781.050 21.380 ;
        RECT 1786.710 21.320 1787.030 21.380 ;
        RECT 1780.730 21.180 1787.030 21.320 ;
        RECT 1780.730 21.120 1781.050 21.180 ;
        RECT 1786.710 21.120 1787.030 21.180 ;
      LAYER via ;
        RECT 1769.260 285.300 1769.520 285.560 ;
        RECT 1780.760 285.300 1781.020 285.560 ;
        RECT 1780.760 21.120 1781.020 21.380 ;
        RECT 1786.740 21.120 1787.000 21.380 ;
      LAYER met2 ;
        RECT 1769.260 300.000 1769.540 304.000 ;
        RECT 1769.320 285.590 1769.460 300.000 ;
        RECT 1769.260 285.270 1769.520 285.590 ;
        RECT 1780.760 285.270 1781.020 285.590 ;
        RECT 1780.820 21.410 1780.960 285.270 ;
        RECT 1780.760 21.090 1781.020 21.410 ;
        RECT 1786.740 21.090 1787.000 21.410 ;
        RECT 1786.800 2.400 1786.940 21.090 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1787.170 20.640 1787.490 20.700 ;
        RECT 1804.650 20.640 1804.970 20.700 ;
        RECT 1787.170 20.500 1804.970 20.640 ;
        RECT 1787.170 20.440 1787.490 20.500 ;
        RECT 1804.650 20.440 1804.970 20.500 ;
      LAYER via ;
        RECT 1787.200 20.440 1787.460 20.700 ;
        RECT 1804.680 20.440 1804.940 20.700 ;
      LAYER met2 ;
        RECT 1783.980 300.290 1784.260 304.000 ;
        RECT 1783.980 300.150 1786.940 300.290 ;
        RECT 1783.980 300.000 1784.260 300.150 ;
        RECT 1786.800 22.170 1786.940 300.150 ;
        RECT 1786.800 22.030 1787.400 22.170 ;
        RECT 1787.260 20.730 1787.400 22.030 ;
        RECT 1787.200 20.410 1787.460 20.730 ;
        RECT 1804.680 20.410 1804.940 20.730 ;
        RECT 1804.740 2.400 1804.880 20.410 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1800.510 19.280 1800.830 19.340 ;
        RECT 1822.590 19.280 1822.910 19.340 ;
        RECT 1800.510 19.140 1822.910 19.280 ;
        RECT 1800.510 19.080 1800.830 19.140 ;
        RECT 1822.590 19.080 1822.910 19.140 ;
      LAYER via ;
        RECT 1800.540 19.080 1800.800 19.340 ;
        RECT 1822.620 19.080 1822.880 19.340 ;
      LAYER met2 ;
        RECT 1798.240 300.290 1798.520 304.000 ;
        RECT 1798.240 300.150 1800.740 300.290 ;
        RECT 1798.240 300.000 1798.520 300.150 ;
        RECT 1800.600 19.370 1800.740 300.150 ;
        RECT 1800.540 19.050 1800.800 19.370 ;
        RECT 1822.620 19.050 1822.880 19.370 ;
        RECT 1822.680 2.400 1822.820 19.050 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1814.310 18.260 1814.630 18.320 ;
        RECT 1840.070 18.260 1840.390 18.320 ;
        RECT 1814.310 18.120 1840.390 18.260 ;
        RECT 1814.310 18.060 1814.630 18.120 ;
        RECT 1840.070 18.060 1840.390 18.120 ;
      LAYER via ;
        RECT 1814.340 18.060 1814.600 18.320 ;
        RECT 1840.100 18.060 1840.360 18.320 ;
      LAYER met2 ;
        RECT 1812.960 300.290 1813.240 304.000 ;
        RECT 1812.960 300.150 1814.540 300.290 ;
        RECT 1812.960 300.000 1813.240 300.150 ;
        RECT 1814.400 18.350 1814.540 300.150 ;
        RECT 1814.340 18.030 1814.600 18.350 ;
        RECT 1840.100 18.030 1840.360 18.350 ;
        RECT 1840.160 2.400 1840.300 18.030 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1828.110 16.560 1828.430 16.620 ;
        RECT 1858.010 16.560 1858.330 16.620 ;
        RECT 1828.110 16.420 1858.330 16.560 ;
        RECT 1828.110 16.360 1828.430 16.420 ;
        RECT 1858.010 16.360 1858.330 16.420 ;
      LAYER via ;
        RECT 1828.140 16.360 1828.400 16.620 ;
        RECT 1858.040 16.360 1858.300 16.620 ;
      LAYER met2 ;
        RECT 1827.680 300.290 1827.960 304.000 ;
        RECT 1827.680 300.150 1828.340 300.290 ;
        RECT 1827.680 300.000 1827.960 300.150 ;
        RECT 1828.200 16.650 1828.340 300.150 ;
        RECT 1828.140 16.330 1828.400 16.650 ;
        RECT 1858.040 16.330 1858.300 16.650 ;
        RECT 1858.100 2.400 1858.240 16.330 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1842.370 288.220 1842.690 288.280 ;
        RECT 1848.350 288.220 1848.670 288.280 ;
        RECT 1842.370 288.080 1848.670 288.220 ;
        RECT 1842.370 288.020 1842.690 288.080 ;
        RECT 1848.350 288.020 1848.670 288.080 ;
        RECT 1848.350 14.520 1848.670 14.580 ;
        RECT 1875.950 14.520 1876.270 14.580 ;
        RECT 1848.350 14.380 1876.270 14.520 ;
        RECT 1848.350 14.320 1848.670 14.380 ;
        RECT 1875.950 14.320 1876.270 14.380 ;
      LAYER via ;
        RECT 1842.400 288.020 1842.660 288.280 ;
        RECT 1848.380 288.020 1848.640 288.280 ;
        RECT 1848.380 14.320 1848.640 14.580 ;
        RECT 1875.980 14.320 1876.240 14.580 ;
      LAYER met2 ;
        RECT 1842.400 300.000 1842.680 304.000 ;
        RECT 1842.460 288.310 1842.600 300.000 ;
        RECT 1842.400 287.990 1842.660 288.310 ;
        RECT 1848.380 287.990 1848.640 288.310 ;
        RECT 1848.440 14.610 1848.580 287.990 ;
        RECT 1848.380 14.290 1848.640 14.610 ;
        RECT 1875.980 14.290 1876.240 14.610 ;
        RECT 1876.040 2.400 1876.180 14.290 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 865.405 282.965 865.575 286.875 ;
        RECT 883.345 286.705 883.515 287.895 ;
      LAYER mcon ;
        RECT 883.345 287.725 883.515 287.895 ;
        RECT 865.405 286.705 865.575 286.875 ;
      LAYER met1 ;
        RECT 883.285 287.880 883.575 287.925 ;
        RECT 916.850 287.880 917.170 287.940 ;
        RECT 883.285 287.740 917.170 287.880 ;
        RECT 883.285 287.695 883.575 287.740 ;
        RECT 916.850 287.680 917.170 287.740 ;
        RECT 865.345 286.860 865.635 286.905 ;
        RECT 883.285 286.860 883.575 286.905 ;
        RECT 865.345 286.720 883.575 286.860 ;
        RECT 865.345 286.675 865.635 286.720 ;
        RECT 883.285 286.675 883.575 286.720 ;
        RECT 824.390 283.120 824.710 283.180 ;
        RECT 865.345 283.120 865.635 283.165 ;
        RECT 824.390 282.980 865.635 283.120 ;
        RECT 824.390 282.920 824.710 282.980 ;
        RECT 865.345 282.935 865.635 282.980 ;
        RECT 752.170 16.900 752.490 16.960 ;
        RECT 824.390 16.900 824.710 16.960 ;
        RECT 752.170 16.760 824.710 16.900 ;
        RECT 752.170 16.700 752.490 16.760 ;
        RECT 824.390 16.700 824.710 16.760 ;
      LAYER via ;
        RECT 916.880 287.680 917.140 287.940 ;
        RECT 824.420 282.920 824.680 283.180 ;
        RECT 752.200 16.700 752.460 16.960 ;
        RECT 824.420 16.700 824.680 16.960 ;
      LAYER met2 ;
        RECT 916.880 300.000 917.160 304.000 ;
        RECT 916.940 287.970 917.080 300.000 ;
        RECT 916.880 287.650 917.140 287.970 ;
        RECT 824.420 282.890 824.680 283.210 ;
        RECT 824.480 16.990 824.620 282.890 ;
        RECT 752.200 16.670 752.460 16.990 ;
        RECT 824.420 16.670 824.680 16.990 ;
        RECT 752.260 2.400 752.400 16.670 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1857.090 288.900 1857.410 288.960 ;
        RECT 1873.190 288.900 1873.510 288.960 ;
        RECT 1857.090 288.760 1873.510 288.900 ;
        RECT 1857.090 288.700 1857.410 288.760 ;
        RECT 1873.190 288.700 1873.510 288.760 ;
        RECT 1873.190 16.560 1873.510 16.620 ;
        RECT 1893.890 16.560 1894.210 16.620 ;
        RECT 1873.190 16.420 1894.210 16.560 ;
        RECT 1873.190 16.360 1873.510 16.420 ;
        RECT 1893.890 16.360 1894.210 16.420 ;
      LAYER via ;
        RECT 1857.120 288.700 1857.380 288.960 ;
        RECT 1873.220 288.700 1873.480 288.960 ;
        RECT 1873.220 16.360 1873.480 16.620 ;
        RECT 1893.920 16.360 1894.180 16.620 ;
      LAYER met2 ;
        RECT 1857.120 300.000 1857.400 304.000 ;
        RECT 1857.180 288.990 1857.320 300.000 ;
        RECT 1857.120 288.670 1857.380 288.990 ;
        RECT 1873.220 288.670 1873.480 288.990 ;
        RECT 1873.280 16.650 1873.420 288.670 ;
        RECT 1873.220 16.330 1873.480 16.650 ;
        RECT 1893.920 16.330 1894.180 16.650 ;
        RECT 1893.980 2.400 1894.120 16.330 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1871.810 288.220 1872.130 288.280 ;
        RECT 1876.410 288.220 1876.730 288.280 ;
        RECT 1871.810 288.080 1876.730 288.220 ;
        RECT 1871.810 288.020 1872.130 288.080 ;
        RECT 1876.410 288.020 1876.730 288.080 ;
        RECT 1876.410 16.900 1876.730 16.960 ;
        RECT 1911.830 16.900 1912.150 16.960 ;
        RECT 1876.410 16.760 1912.150 16.900 ;
        RECT 1876.410 16.700 1876.730 16.760 ;
        RECT 1911.830 16.700 1912.150 16.760 ;
      LAYER via ;
        RECT 1871.840 288.020 1872.100 288.280 ;
        RECT 1876.440 288.020 1876.700 288.280 ;
        RECT 1876.440 16.700 1876.700 16.960 ;
        RECT 1911.860 16.700 1912.120 16.960 ;
      LAYER met2 ;
        RECT 1871.840 300.000 1872.120 304.000 ;
        RECT 1871.900 288.310 1872.040 300.000 ;
        RECT 1871.840 287.990 1872.100 288.310 ;
        RECT 1876.440 287.990 1876.700 288.310 ;
        RECT 1876.500 16.990 1876.640 287.990 ;
        RECT 1876.440 16.670 1876.700 16.990 ;
        RECT 1911.860 16.670 1912.120 16.990 ;
        RECT 1911.920 2.400 1912.060 16.670 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1890.210 15.880 1890.530 15.940 ;
        RECT 1929.310 15.880 1929.630 15.940 ;
        RECT 1890.210 15.740 1929.630 15.880 ;
        RECT 1890.210 15.680 1890.530 15.740 ;
        RECT 1929.310 15.680 1929.630 15.740 ;
      LAYER via ;
        RECT 1890.240 15.680 1890.500 15.940 ;
        RECT 1929.340 15.680 1929.600 15.940 ;
      LAYER met2 ;
        RECT 1886.560 300.290 1886.840 304.000 ;
        RECT 1886.560 300.150 1890.440 300.290 ;
        RECT 1886.560 300.000 1886.840 300.150 ;
        RECT 1890.300 15.970 1890.440 300.150 ;
        RECT 1890.240 15.650 1890.500 15.970 ;
        RECT 1929.340 15.650 1929.600 15.970 ;
        RECT 1929.400 2.400 1929.540 15.650 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1904.010 18.940 1904.330 19.000 ;
        RECT 1947.250 18.940 1947.570 19.000 ;
        RECT 1904.010 18.800 1947.570 18.940 ;
        RECT 1904.010 18.740 1904.330 18.800 ;
        RECT 1947.250 18.740 1947.570 18.800 ;
      LAYER via ;
        RECT 1904.040 18.740 1904.300 19.000 ;
        RECT 1947.280 18.740 1947.540 19.000 ;
      LAYER met2 ;
        RECT 1901.280 300.290 1901.560 304.000 ;
        RECT 1901.280 300.150 1904.240 300.290 ;
        RECT 1901.280 300.000 1901.560 300.150 ;
        RECT 1904.100 19.030 1904.240 300.150 ;
        RECT 1904.040 18.710 1904.300 19.030 ;
        RECT 1947.280 18.710 1947.540 19.030 ;
        RECT 1947.340 2.400 1947.480 18.710 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1917.810 19.280 1918.130 19.340 ;
        RECT 1965.190 19.280 1965.510 19.340 ;
        RECT 1917.810 19.140 1965.510 19.280 ;
        RECT 1917.810 19.080 1918.130 19.140 ;
        RECT 1965.190 19.080 1965.510 19.140 ;
      LAYER via ;
        RECT 1917.840 19.080 1918.100 19.340 ;
        RECT 1965.220 19.080 1965.480 19.340 ;
      LAYER met2 ;
        RECT 1916.000 300.290 1916.280 304.000 ;
        RECT 1916.000 300.150 1918.040 300.290 ;
        RECT 1916.000 300.000 1916.280 300.150 ;
        RECT 1917.900 19.370 1918.040 300.150 ;
        RECT 1917.840 19.050 1918.100 19.370 ;
        RECT 1965.220 19.050 1965.480 19.370 ;
        RECT 1965.280 2.400 1965.420 19.050 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1931.150 17.580 1931.470 17.640 ;
        RECT 1983.130 17.580 1983.450 17.640 ;
        RECT 1931.150 17.440 1983.450 17.580 ;
        RECT 1931.150 17.380 1931.470 17.440 ;
        RECT 1983.130 17.380 1983.450 17.440 ;
      LAYER via ;
        RECT 1931.180 17.380 1931.440 17.640 ;
        RECT 1983.160 17.380 1983.420 17.640 ;
      LAYER met2 ;
        RECT 1930.720 300.290 1931.000 304.000 ;
        RECT 1930.720 300.150 1931.380 300.290 ;
        RECT 1930.720 300.000 1931.000 300.150 ;
        RECT 1931.240 17.670 1931.380 300.150 ;
        RECT 1931.180 17.350 1931.440 17.670 ;
        RECT 1983.160 17.350 1983.420 17.670 ;
        RECT 1983.220 2.400 1983.360 17.350 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1944.950 17.240 1945.270 17.300 ;
        RECT 2001.070 17.240 2001.390 17.300 ;
        RECT 1944.950 17.100 2001.390 17.240 ;
        RECT 1944.950 17.040 1945.270 17.100 ;
        RECT 2001.070 17.040 2001.390 17.100 ;
      LAYER via ;
        RECT 1944.980 17.040 1945.240 17.300 ;
        RECT 2001.100 17.040 2001.360 17.300 ;
      LAYER met2 ;
        RECT 1945.440 300.290 1945.720 304.000 ;
        RECT 1945.040 300.150 1945.720 300.290 ;
        RECT 1945.040 17.330 1945.180 300.150 ;
        RECT 1945.440 300.000 1945.720 300.150 ;
        RECT 1944.980 17.010 1945.240 17.330 ;
        RECT 2001.100 17.010 2001.360 17.330 ;
        RECT 2001.160 2.400 2001.300 17.010 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1960.130 288.220 1960.450 288.280 ;
        RECT 1966.110 288.220 1966.430 288.280 ;
        RECT 1960.130 288.080 1966.430 288.220 ;
        RECT 1960.130 288.020 1960.450 288.080 ;
        RECT 1966.110 288.020 1966.430 288.080 ;
        RECT 1966.110 19.280 1966.430 19.340 ;
        RECT 2018.550 19.280 2018.870 19.340 ;
        RECT 1966.110 19.140 2018.870 19.280 ;
        RECT 1966.110 19.080 1966.430 19.140 ;
        RECT 2018.550 19.080 2018.870 19.140 ;
      LAYER via ;
        RECT 1960.160 288.020 1960.420 288.280 ;
        RECT 1966.140 288.020 1966.400 288.280 ;
        RECT 1966.140 19.080 1966.400 19.340 ;
        RECT 2018.580 19.080 2018.840 19.340 ;
      LAYER met2 ;
        RECT 1960.160 300.000 1960.440 304.000 ;
        RECT 1960.220 288.310 1960.360 300.000 ;
        RECT 1960.160 287.990 1960.420 288.310 ;
        RECT 1966.140 287.990 1966.400 288.310 ;
        RECT 1966.200 19.370 1966.340 287.990 ;
        RECT 1966.140 19.050 1966.400 19.370 ;
        RECT 2018.580 19.050 2018.840 19.370 ;
        RECT 2018.640 2.400 2018.780 19.050 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1974.850 288.220 1975.170 288.280 ;
        RECT 1979.450 288.220 1979.770 288.280 ;
        RECT 1974.850 288.080 1979.770 288.220 ;
        RECT 1974.850 288.020 1975.170 288.080 ;
        RECT 1979.450 288.020 1979.770 288.080 ;
        RECT 1979.450 20.300 1979.770 20.360 ;
        RECT 2036.490 20.300 2036.810 20.360 ;
        RECT 1979.450 20.160 2036.810 20.300 ;
        RECT 1979.450 20.100 1979.770 20.160 ;
        RECT 2036.490 20.100 2036.810 20.160 ;
      LAYER via ;
        RECT 1974.880 288.020 1975.140 288.280 ;
        RECT 1979.480 288.020 1979.740 288.280 ;
        RECT 1979.480 20.100 1979.740 20.360 ;
        RECT 2036.520 20.100 2036.780 20.360 ;
      LAYER met2 ;
        RECT 1974.880 300.000 1975.160 304.000 ;
        RECT 1974.940 288.310 1975.080 300.000 ;
        RECT 1974.880 287.990 1975.140 288.310 ;
        RECT 1979.480 287.990 1979.740 288.310 ;
        RECT 1979.540 20.390 1979.680 287.990 ;
        RECT 1979.480 20.070 1979.740 20.390 ;
        RECT 2036.520 20.070 2036.780 20.390 ;
        RECT 2036.580 2.400 2036.720 20.070 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1989.570 288.220 1989.890 288.280 ;
        RECT 1993.710 288.220 1994.030 288.280 ;
        RECT 1989.570 288.080 1994.030 288.220 ;
        RECT 1989.570 288.020 1989.890 288.080 ;
        RECT 1993.710 288.020 1994.030 288.080 ;
        RECT 1993.710 16.560 1994.030 16.620 ;
        RECT 2054.430 16.560 2054.750 16.620 ;
        RECT 1993.710 16.420 2054.750 16.560 ;
        RECT 1993.710 16.360 1994.030 16.420 ;
        RECT 2054.430 16.360 2054.750 16.420 ;
      LAYER via ;
        RECT 1989.600 288.020 1989.860 288.280 ;
        RECT 1993.740 288.020 1994.000 288.280 ;
        RECT 1993.740 16.360 1994.000 16.620 ;
        RECT 2054.460 16.360 2054.720 16.620 ;
      LAYER met2 ;
        RECT 1989.600 300.000 1989.880 304.000 ;
        RECT 1989.660 288.310 1989.800 300.000 ;
        RECT 1989.600 287.990 1989.860 288.310 ;
        RECT 1993.740 287.990 1994.000 288.310 ;
        RECT 1993.800 16.650 1993.940 287.990 ;
        RECT 1993.740 16.330 1994.000 16.650 ;
        RECT 2054.460 16.330 2054.720 16.650 ;
        RECT 2054.520 2.400 2054.660 16.330 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 855.745 282.625 855.915 283.475 ;
      LAYER mcon ;
        RECT 855.745 283.305 855.915 283.475 ;
      LAYER met1 ;
        RECT 845.090 283.460 845.410 283.520 ;
        RECT 855.685 283.460 855.975 283.505 ;
        RECT 845.090 283.320 855.975 283.460 ;
        RECT 845.090 283.260 845.410 283.320 ;
        RECT 855.685 283.275 855.975 283.320 ;
        RECT 855.685 282.780 855.975 282.825 ;
        RECT 931.570 282.780 931.890 282.840 ;
        RECT 855.685 282.640 931.890 282.780 ;
        RECT 855.685 282.595 855.975 282.640 ;
        RECT 931.570 282.580 931.890 282.640 ;
        RECT 769.650 19.620 769.970 19.680 ;
        RECT 845.090 19.620 845.410 19.680 ;
        RECT 769.650 19.480 845.410 19.620 ;
        RECT 769.650 19.420 769.970 19.480 ;
        RECT 845.090 19.420 845.410 19.480 ;
      LAYER via ;
        RECT 845.120 283.260 845.380 283.520 ;
        RECT 931.600 282.580 931.860 282.840 ;
        RECT 769.680 19.420 769.940 19.680 ;
        RECT 845.120 19.420 845.380 19.680 ;
      LAYER met2 ;
        RECT 931.600 300.000 931.880 304.000 ;
        RECT 845.120 283.230 845.380 283.550 ;
        RECT 845.180 19.710 845.320 283.230 ;
        RECT 931.660 282.870 931.800 300.000 ;
        RECT 931.600 282.550 931.860 282.870 ;
        RECT 769.680 19.390 769.940 19.710 ;
        RECT 845.120 19.390 845.380 19.710 ;
        RECT 769.740 2.400 769.880 19.390 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2007.510 18.940 2007.830 19.000 ;
        RECT 2072.370 18.940 2072.690 19.000 ;
        RECT 2007.510 18.800 2072.690 18.940 ;
        RECT 2007.510 18.740 2007.830 18.800 ;
        RECT 2072.370 18.740 2072.690 18.800 ;
      LAYER via ;
        RECT 2007.540 18.740 2007.800 19.000 ;
        RECT 2072.400 18.740 2072.660 19.000 ;
      LAYER met2 ;
        RECT 2004.320 300.290 2004.600 304.000 ;
        RECT 2004.320 300.150 2007.740 300.290 ;
        RECT 2004.320 300.000 2004.600 300.150 ;
        RECT 2007.600 19.030 2007.740 300.150 ;
        RECT 2007.540 18.710 2007.800 19.030 ;
        RECT 2072.400 18.710 2072.660 19.030 ;
        RECT 2072.460 2.400 2072.600 18.710 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2021.310 19.280 2021.630 19.340 ;
        RECT 2089.850 19.280 2090.170 19.340 ;
        RECT 2021.310 19.140 2090.170 19.280 ;
        RECT 2021.310 19.080 2021.630 19.140 ;
        RECT 2089.850 19.080 2090.170 19.140 ;
      LAYER via ;
        RECT 2021.340 19.080 2021.600 19.340 ;
        RECT 2089.880 19.080 2090.140 19.340 ;
      LAYER met2 ;
        RECT 2019.040 300.290 2019.320 304.000 ;
        RECT 2019.040 300.150 2021.540 300.290 ;
        RECT 2019.040 300.000 2019.320 300.150 ;
        RECT 2021.400 19.370 2021.540 300.150 ;
        RECT 2021.340 19.050 2021.600 19.370 ;
        RECT 2089.880 19.050 2090.140 19.370 ;
        RECT 2089.940 2.400 2090.080 19.050 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2035.110 19.620 2035.430 19.680 ;
        RECT 2107.790 19.620 2108.110 19.680 ;
        RECT 2035.110 19.480 2108.110 19.620 ;
        RECT 2035.110 19.420 2035.430 19.480 ;
        RECT 2107.790 19.420 2108.110 19.480 ;
      LAYER via ;
        RECT 2035.140 19.420 2035.400 19.680 ;
        RECT 2107.820 19.420 2108.080 19.680 ;
      LAYER met2 ;
        RECT 2033.760 300.290 2034.040 304.000 ;
        RECT 2033.760 300.150 2035.340 300.290 ;
        RECT 2033.760 300.000 2034.040 300.150 ;
        RECT 2035.200 19.710 2035.340 300.150 ;
        RECT 2035.140 19.390 2035.400 19.710 ;
        RECT 2107.820 19.390 2108.080 19.710 ;
        RECT 2107.880 2.400 2108.020 19.390 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2048.910 17.920 2049.230 17.980 ;
        RECT 2125.730 17.920 2126.050 17.980 ;
        RECT 2048.910 17.780 2126.050 17.920 ;
        RECT 2048.910 17.720 2049.230 17.780 ;
        RECT 2125.730 17.720 2126.050 17.780 ;
      LAYER via ;
        RECT 2048.940 17.720 2049.200 17.980 ;
        RECT 2125.760 17.720 2126.020 17.980 ;
      LAYER met2 ;
        RECT 2048.020 300.290 2048.300 304.000 ;
        RECT 2048.020 300.150 2049.140 300.290 ;
        RECT 2048.020 300.000 2048.300 300.150 ;
        RECT 2049.000 18.010 2049.140 300.150 ;
        RECT 2048.940 17.690 2049.200 18.010 ;
        RECT 2125.760 17.690 2126.020 18.010 ;
        RECT 2125.820 2.400 2125.960 17.690 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2062.710 19.960 2063.030 20.020 ;
        RECT 2143.670 19.960 2143.990 20.020 ;
        RECT 2062.710 19.820 2143.990 19.960 ;
        RECT 2062.710 19.760 2063.030 19.820 ;
        RECT 2143.670 19.760 2143.990 19.820 ;
      LAYER via ;
        RECT 2062.740 19.760 2063.000 20.020 ;
        RECT 2143.700 19.760 2143.960 20.020 ;
      LAYER met2 ;
        RECT 2062.740 300.000 2063.020 304.000 ;
        RECT 2062.800 20.050 2062.940 300.000 ;
        RECT 2062.740 19.730 2063.000 20.050 ;
        RECT 2143.700 19.730 2143.960 20.050 ;
        RECT 2143.760 2.400 2143.900 19.730 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2077.430 286.180 2077.750 286.240 ;
        RECT 2083.410 286.180 2083.730 286.240 ;
        RECT 2077.430 286.040 2083.730 286.180 ;
        RECT 2077.430 285.980 2077.750 286.040 ;
        RECT 2083.410 285.980 2083.730 286.040 ;
        RECT 2083.410 16.560 2083.730 16.620 ;
        RECT 2161.610 16.560 2161.930 16.620 ;
        RECT 2083.410 16.420 2161.930 16.560 ;
        RECT 2083.410 16.360 2083.730 16.420 ;
        RECT 2161.610 16.360 2161.930 16.420 ;
      LAYER via ;
        RECT 2077.460 285.980 2077.720 286.240 ;
        RECT 2083.440 285.980 2083.700 286.240 ;
        RECT 2083.440 16.360 2083.700 16.620 ;
        RECT 2161.640 16.360 2161.900 16.620 ;
      LAYER met2 ;
        RECT 2077.460 300.000 2077.740 304.000 ;
        RECT 2077.520 286.270 2077.660 300.000 ;
        RECT 2077.460 285.950 2077.720 286.270 ;
        RECT 2083.440 285.950 2083.700 286.270 ;
        RECT 2083.500 16.650 2083.640 285.950 ;
        RECT 2083.440 16.330 2083.700 16.650 ;
        RECT 2161.640 16.330 2161.900 16.650 ;
        RECT 2161.700 2.400 2161.840 16.330 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2092.150 288.220 2092.470 288.280 ;
        RECT 2097.210 288.220 2097.530 288.280 ;
        RECT 2092.150 288.080 2097.530 288.220 ;
        RECT 2092.150 288.020 2092.470 288.080 ;
        RECT 2097.210 288.020 2097.530 288.080 ;
        RECT 2097.210 16.900 2097.530 16.960 ;
        RECT 2179.090 16.900 2179.410 16.960 ;
        RECT 2097.210 16.760 2179.410 16.900 ;
        RECT 2097.210 16.700 2097.530 16.760 ;
        RECT 2179.090 16.700 2179.410 16.760 ;
      LAYER via ;
        RECT 2092.180 288.020 2092.440 288.280 ;
        RECT 2097.240 288.020 2097.500 288.280 ;
        RECT 2097.240 16.700 2097.500 16.960 ;
        RECT 2179.120 16.700 2179.380 16.960 ;
      LAYER met2 ;
        RECT 2092.180 300.000 2092.460 304.000 ;
        RECT 2092.240 288.310 2092.380 300.000 ;
        RECT 2092.180 287.990 2092.440 288.310 ;
        RECT 2097.240 287.990 2097.500 288.310 ;
        RECT 2097.300 16.990 2097.440 287.990 ;
        RECT 2097.240 16.670 2097.500 16.990 ;
        RECT 2179.120 16.670 2179.380 16.990 ;
        RECT 2179.180 2.400 2179.320 16.670 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2106.870 288.220 2107.190 288.280 ;
        RECT 2111.010 288.220 2111.330 288.280 ;
        RECT 2106.870 288.080 2111.330 288.220 ;
        RECT 2106.870 288.020 2107.190 288.080 ;
        RECT 2111.010 288.020 2111.330 288.080 ;
        RECT 2111.010 15.200 2111.330 15.260 ;
        RECT 2197.030 15.200 2197.350 15.260 ;
        RECT 2111.010 15.060 2197.350 15.200 ;
        RECT 2111.010 15.000 2111.330 15.060 ;
        RECT 2197.030 15.000 2197.350 15.060 ;
      LAYER via ;
        RECT 2106.900 288.020 2107.160 288.280 ;
        RECT 2111.040 288.020 2111.300 288.280 ;
        RECT 2111.040 15.000 2111.300 15.260 ;
        RECT 2197.060 15.000 2197.320 15.260 ;
      LAYER met2 ;
        RECT 2106.900 300.000 2107.180 304.000 ;
        RECT 2106.960 288.310 2107.100 300.000 ;
        RECT 2106.900 287.990 2107.160 288.310 ;
        RECT 2111.040 287.990 2111.300 288.310 ;
        RECT 2111.100 15.290 2111.240 287.990 ;
        RECT 2111.040 14.970 2111.300 15.290 ;
        RECT 2197.060 14.970 2197.320 15.290 ;
        RECT 2197.120 2.400 2197.260 14.970 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2124.810 16.220 2125.130 16.280 ;
        RECT 2214.970 16.220 2215.290 16.280 ;
        RECT 2124.810 16.080 2215.290 16.220 ;
        RECT 2124.810 16.020 2125.130 16.080 ;
        RECT 2214.970 16.020 2215.290 16.080 ;
      LAYER via ;
        RECT 2124.840 16.020 2125.100 16.280 ;
        RECT 2215.000 16.020 2215.260 16.280 ;
      LAYER met2 ;
        RECT 2121.620 300.290 2121.900 304.000 ;
        RECT 2121.620 300.150 2125.040 300.290 ;
        RECT 2121.620 300.000 2121.900 300.150 ;
        RECT 2124.900 16.310 2125.040 300.150 ;
        RECT 2124.840 15.990 2125.100 16.310 ;
        RECT 2215.000 15.990 2215.260 16.310 ;
        RECT 2215.060 2.400 2215.200 15.990 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2138.610 15.880 2138.930 15.940 ;
        RECT 2232.910 15.880 2233.230 15.940 ;
        RECT 2138.610 15.740 2233.230 15.880 ;
        RECT 2138.610 15.680 2138.930 15.740 ;
        RECT 2232.910 15.680 2233.230 15.740 ;
      LAYER via ;
        RECT 2138.640 15.680 2138.900 15.940 ;
        RECT 2232.940 15.680 2233.200 15.940 ;
      LAYER met2 ;
        RECT 2136.340 300.290 2136.620 304.000 ;
        RECT 2136.340 300.150 2138.840 300.290 ;
        RECT 2136.340 300.000 2136.620 300.150 ;
        RECT 2138.700 15.970 2138.840 300.150 ;
        RECT 2138.640 15.650 2138.900 15.970 ;
        RECT 2232.940 15.650 2233.200 15.970 ;
        RECT 2233.000 2.400 2233.140 15.650 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.110 289.580 793.430 289.640 ;
        RECT 946.290 289.580 946.610 289.640 ;
        RECT 793.110 289.440 946.610 289.580 ;
        RECT 793.110 289.380 793.430 289.440 ;
        RECT 946.290 289.380 946.610 289.440 ;
        RECT 787.590 17.240 787.910 17.300 ;
        RECT 793.110 17.240 793.430 17.300 ;
        RECT 787.590 17.100 793.430 17.240 ;
        RECT 787.590 17.040 787.910 17.100 ;
        RECT 793.110 17.040 793.430 17.100 ;
      LAYER via ;
        RECT 793.140 289.380 793.400 289.640 ;
        RECT 946.320 289.380 946.580 289.640 ;
        RECT 787.620 17.040 787.880 17.300 ;
        RECT 793.140 17.040 793.400 17.300 ;
      LAYER met2 ;
        RECT 946.320 300.000 946.600 304.000 ;
        RECT 946.380 289.670 946.520 300.000 ;
        RECT 793.140 289.350 793.400 289.670 ;
        RECT 946.320 289.350 946.580 289.670 ;
        RECT 793.200 17.330 793.340 289.350 ;
        RECT 787.620 17.010 787.880 17.330 ;
        RECT 793.140 17.010 793.400 17.330 ;
        RECT 787.680 2.400 787.820 17.010 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2156.165 18.785 2156.335 20.655 ;
        RECT 2165.825 14.025 2165.995 18.955 ;
        RECT 2227.465 14.025 2227.635 17.935 ;
      LAYER mcon ;
        RECT 2156.165 20.485 2156.335 20.655 ;
        RECT 2165.825 18.785 2165.995 18.955 ;
        RECT 2227.465 17.765 2227.635 17.935 ;
      LAYER met1 ;
        RECT 2151.950 20.640 2152.270 20.700 ;
        RECT 2156.105 20.640 2156.395 20.685 ;
        RECT 2151.950 20.500 2156.395 20.640 ;
        RECT 2151.950 20.440 2152.270 20.500 ;
        RECT 2156.105 20.455 2156.395 20.500 ;
        RECT 2156.105 18.940 2156.395 18.985 ;
        RECT 2165.765 18.940 2166.055 18.985 ;
        RECT 2156.105 18.800 2166.055 18.940 ;
        RECT 2156.105 18.755 2156.395 18.800 ;
        RECT 2165.765 18.755 2166.055 18.800 ;
        RECT 2227.405 17.920 2227.695 17.965 ;
        RECT 2250.850 17.920 2251.170 17.980 ;
        RECT 2227.405 17.780 2251.170 17.920 ;
        RECT 2227.405 17.735 2227.695 17.780 ;
        RECT 2250.850 17.720 2251.170 17.780 ;
        RECT 2165.765 14.180 2166.055 14.225 ;
        RECT 2227.405 14.180 2227.695 14.225 ;
        RECT 2165.765 14.040 2227.695 14.180 ;
        RECT 2165.765 13.995 2166.055 14.040 ;
        RECT 2227.405 13.995 2227.695 14.040 ;
      LAYER via ;
        RECT 2151.980 20.440 2152.240 20.700 ;
        RECT 2250.880 17.720 2251.140 17.980 ;
      LAYER met2 ;
        RECT 2151.060 300.290 2151.340 304.000 ;
        RECT 2151.060 300.150 2152.180 300.290 ;
        RECT 2151.060 300.000 2151.340 300.150 ;
        RECT 2152.040 20.730 2152.180 300.150 ;
        RECT 2151.980 20.410 2152.240 20.730 ;
        RECT 2250.880 17.690 2251.140 18.010 ;
        RECT 2250.940 2.400 2251.080 17.690 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2233.445 15.725 2233.615 18.615 ;
      LAYER mcon ;
        RECT 2233.445 18.445 2233.615 18.615 ;
      LAYER met1 ;
        RECT 2166.210 18.940 2166.530 19.000 ;
        RECT 2166.210 18.800 2211.520 18.940 ;
        RECT 2166.210 18.740 2166.530 18.800 ;
        RECT 2211.380 18.600 2211.520 18.800 ;
        RECT 2233.385 18.600 2233.675 18.645 ;
        RECT 2211.380 18.460 2233.675 18.600 ;
        RECT 2233.385 18.415 2233.675 18.460 ;
        RECT 2233.385 15.880 2233.675 15.925 ;
        RECT 2262.810 15.880 2263.130 15.940 ;
        RECT 2233.385 15.740 2263.130 15.880 ;
        RECT 2233.385 15.695 2233.675 15.740 ;
        RECT 2262.810 15.680 2263.130 15.740 ;
        RECT 2263.270 14.180 2263.590 14.240 ;
        RECT 2268.330 14.180 2268.650 14.240 ;
        RECT 2263.270 14.040 2268.650 14.180 ;
        RECT 2263.270 13.980 2263.590 14.040 ;
        RECT 2268.330 13.980 2268.650 14.040 ;
      LAYER via ;
        RECT 2166.240 18.740 2166.500 19.000 ;
        RECT 2262.840 15.680 2263.100 15.940 ;
        RECT 2263.300 13.980 2263.560 14.240 ;
        RECT 2268.360 13.980 2268.620 14.240 ;
      LAYER met2 ;
        RECT 2165.780 300.290 2166.060 304.000 ;
        RECT 2165.780 300.150 2166.440 300.290 ;
        RECT 2165.780 300.000 2166.060 300.150 ;
        RECT 2166.300 19.030 2166.440 300.150 ;
        RECT 2166.240 18.710 2166.500 19.030 ;
        RECT 2262.900 15.970 2263.500 16.050 ;
        RECT 2262.840 15.910 2263.500 15.970 ;
        RECT 2262.840 15.650 2263.100 15.910 ;
        RECT 2263.360 14.270 2263.500 15.910 ;
        RECT 2263.300 13.950 2263.560 14.270 ;
        RECT 2268.360 13.950 2268.620 14.270 ;
        RECT 2268.420 2.400 2268.560 13.950 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.470 285.500 2180.790 285.560 ;
        RECT 2186.910 285.500 2187.230 285.560 ;
        RECT 2180.470 285.360 2187.230 285.500 ;
        RECT 2180.470 285.300 2180.790 285.360 ;
        RECT 2186.910 285.300 2187.230 285.360 ;
        RECT 2186.910 16.900 2187.230 16.960 ;
        RECT 2286.270 16.900 2286.590 16.960 ;
        RECT 2186.910 16.760 2286.590 16.900 ;
        RECT 2186.910 16.700 2187.230 16.760 ;
        RECT 2286.270 16.700 2286.590 16.760 ;
      LAYER via ;
        RECT 2180.500 285.300 2180.760 285.560 ;
        RECT 2186.940 285.300 2187.200 285.560 ;
        RECT 2186.940 16.700 2187.200 16.960 ;
        RECT 2286.300 16.700 2286.560 16.960 ;
      LAYER met2 ;
        RECT 2180.500 300.000 2180.780 304.000 ;
        RECT 2180.560 285.590 2180.700 300.000 ;
        RECT 2180.500 285.270 2180.760 285.590 ;
        RECT 2186.940 285.270 2187.200 285.590 ;
        RECT 2187.000 16.990 2187.140 285.270 ;
        RECT 2186.940 16.670 2187.200 16.990 ;
        RECT 2286.300 16.670 2286.560 16.990 ;
        RECT 2286.360 2.400 2286.500 16.670 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2227.925 14.025 2228.095 15.215 ;
      LAYER mcon ;
        RECT 2227.925 15.045 2228.095 15.215 ;
      LAYER met1 ;
        RECT 2195.190 288.220 2195.510 288.280 ;
        RECT 2200.710 288.220 2201.030 288.280 ;
        RECT 2195.190 288.080 2201.030 288.220 ;
        RECT 2195.190 288.020 2195.510 288.080 ;
        RECT 2200.710 288.020 2201.030 288.080 ;
        RECT 2200.710 15.200 2201.030 15.260 ;
        RECT 2227.865 15.200 2228.155 15.245 ;
        RECT 2200.710 15.060 2228.155 15.200 ;
        RECT 2200.710 15.000 2201.030 15.060 ;
        RECT 2227.865 15.015 2228.155 15.060 ;
        RECT 2227.865 14.180 2228.155 14.225 ;
        RECT 2303.750 14.180 2304.070 14.240 ;
        RECT 2227.865 14.040 2263.040 14.180 ;
        RECT 2227.865 13.995 2228.155 14.040 ;
        RECT 2262.900 13.840 2263.040 14.040 ;
        RECT 2268.880 14.040 2304.070 14.180 ;
        RECT 2268.880 13.840 2269.020 14.040 ;
        RECT 2303.750 13.980 2304.070 14.040 ;
        RECT 2262.900 13.700 2269.020 13.840 ;
      LAYER via ;
        RECT 2195.220 288.020 2195.480 288.280 ;
        RECT 2200.740 288.020 2201.000 288.280 ;
        RECT 2200.740 15.000 2201.000 15.260 ;
        RECT 2303.780 13.980 2304.040 14.240 ;
      LAYER met2 ;
        RECT 2195.220 300.000 2195.500 304.000 ;
        RECT 2195.280 288.310 2195.420 300.000 ;
        RECT 2195.220 287.990 2195.480 288.310 ;
        RECT 2200.740 287.990 2201.000 288.310 ;
        RECT 2200.800 15.290 2200.940 287.990 ;
        RECT 2200.740 14.970 2201.000 15.290 ;
        RECT 2303.780 14.010 2304.040 14.270 ;
        RECT 2303.780 13.950 2304.440 14.010 ;
        RECT 2303.840 13.870 2304.440 13.950 ;
        RECT 2304.300 2.400 2304.440 13.870 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2209.910 288.220 2210.230 288.280 ;
        RECT 2214.510 288.220 2214.830 288.280 ;
        RECT 2209.910 288.080 2214.830 288.220 ;
        RECT 2209.910 288.020 2210.230 288.080 ;
        RECT 2214.510 288.020 2214.830 288.080 ;
        RECT 2214.510 14.860 2214.830 14.920 ;
        RECT 2322.150 14.860 2322.470 14.920 ;
        RECT 2214.510 14.720 2322.470 14.860 ;
        RECT 2214.510 14.660 2214.830 14.720 ;
        RECT 2322.150 14.660 2322.470 14.720 ;
      LAYER via ;
        RECT 2209.940 288.020 2210.200 288.280 ;
        RECT 2214.540 288.020 2214.800 288.280 ;
        RECT 2214.540 14.660 2214.800 14.920 ;
        RECT 2322.180 14.660 2322.440 14.920 ;
      LAYER met2 ;
        RECT 2209.940 300.000 2210.220 304.000 ;
        RECT 2210.000 288.310 2210.140 300.000 ;
        RECT 2209.940 287.990 2210.200 288.310 ;
        RECT 2214.540 287.990 2214.800 288.310 ;
        RECT 2214.600 14.950 2214.740 287.990 ;
        RECT 2214.540 14.630 2214.800 14.950 ;
        RECT 2322.180 14.630 2322.440 14.950 ;
        RECT 2322.240 2.400 2322.380 14.630 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2268.865 15.385 2269.035 18.955 ;
      LAYER mcon ;
        RECT 2268.865 18.785 2269.035 18.955 ;
      LAYER met1 ;
        RECT 2224.630 286.860 2224.950 286.920 ;
        RECT 2228.310 286.860 2228.630 286.920 ;
        RECT 2224.630 286.720 2228.630 286.860 ;
        RECT 2224.630 286.660 2224.950 286.720 ;
        RECT 2228.310 286.660 2228.630 286.720 ;
        RECT 2228.310 18.940 2228.630 19.000 ;
        RECT 2268.805 18.940 2269.095 18.985 ;
        RECT 2228.310 18.800 2269.095 18.940 ;
        RECT 2228.310 18.740 2228.630 18.800 ;
        RECT 2268.805 18.755 2269.095 18.800 ;
        RECT 2268.805 15.540 2269.095 15.585 ;
        RECT 2339.630 15.540 2339.950 15.600 ;
        RECT 2268.805 15.400 2339.950 15.540 ;
        RECT 2268.805 15.355 2269.095 15.400 ;
        RECT 2339.630 15.340 2339.950 15.400 ;
      LAYER via ;
        RECT 2224.660 286.660 2224.920 286.920 ;
        RECT 2228.340 286.660 2228.600 286.920 ;
        RECT 2228.340 18.740 2228.600 19.000 ;
        RECT 2339.660 15.340 2339.920 15.600 ;
      LAYER met2 ;
        RECT 2224.660 300.000 2224.940 304.000 ;
        RECT 2224.720 286.950 2224.860 300.000 ;
        RECT 2224.660 286.630 2224.920 286.950 ;
        RECT 2228.340 286.630 2228.600 286.950 ;
        RECT 2228.400 19.030 2228.540 286.630 ;
        RECT 2228.340 18.710 2228.600 19.030 ;
        RECT 2339.660 15.310 2339.920 15.630 ;
        RECT 2339.720 2.400 2339.860 15.310 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2328.665 17.425 2329.755 17.595 ;
        RECT 2328.665 15.725 2328.835 17.425 ;
      LAYER mcon ;
        RECT 2329.585 17.425 2329.755 17.595 ;
      LAYER met1 ;
        RECT 2329.525 17.580 2329.815 17.625 ;
        RECT 2357.570 17.580 2357.890 17.640 ;
        RECT 2329.525 17.440 2357.890 17.580 ;
        RECT 2329.525 17.395 2329.815 17.440 ;
        RECT 2357.570 17.380 2357.890 17.440 ;
        RECT 2328.605 15.880 2328.895 15.925 ;
        RECT 2263.360 15.740 2328.895 15.880 ;
        RECT 2242.110 15.540 2242.430 15.600 ;
        RECT 2263.360 15.540 2263.500 15.740 ;
        RECT 2328.605 15.695 2328.895 15.740 ;
        RECT 2242.110 15.400 2263.500 15.540 ;
        RECT 2242.110 15.340 2242.430 15.400 ;
      LAYER via ;
        RECT 2357.600 17.380 2357.860 17.640 ;
        RECT 2242.140 15.340 2242.400 15.600 ;
      LAYER met2 ;
        RECT 2239.380 300.290 2239.660 304.000 ;
        RECT 2239.380 300.150 2242.340 300.290 ;
        RECT 2239.380 300.000 2239.660 300.150 ;
        RECT 2242.200 15.630 2242.340 300.150 ;
        RECT 2357.600 17.350 2357.860 17.670 ;
        RECT 2242.140 15.310 2242.400 15.630 ;
        RECT 2357.660 2.400 2357.800 17.350 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2279.905 16.405 2280.075 17.935 ;
      LAYER mcon ;
        RECT 2279.905 17.765 2280.075 17.935 ;
      LAYER met1 ;
        RECT 2255.910 17.920 2256.230 17.980 ;
        RECT 2279.845 17.920 2280.135 17.965 ;
        RECT 2255.910 17.780 2280.135 17.920 ;
        RECT 2255.910 17.720 2256.230 17.780 ;
        RECT 2279.845 17.735 2280.135 17.780 ;
        RECT 2279.845 16.560 2280.135 16.605 ;
        RECT 2375.510 16.560 2375.830 16.620 ;
        RECT 2279.845 16.420 2375.830 16.560 ;
        RECT 2279.845 16.375 2280.135 16.420 ;
        RECT 2375.510 16.360 2375.830 16.420 ;
      LAYER via ;
        RECT 2255.940 17.720 2256.200 17.980 ;
        RECT 2375.540 16.360 2375.800 16.620 ;
      LAYER met2 ;
        RECT 2254.100 300.290 2254.380 304.000 ;
        RECT 2254.100 300.150 2256.140 300.290 ;
        RECT 2254.100 300.000 2254.380 300.150 ;
        RECT 2256.000 18.010 2256.140 300.150 ;
        RECT 2255.940 17.690 2256.200 18.010 ;
        RECT 2375.540 16.330 2375.800 16.650 ;
        RECT 2375.600 2.400 2375.740 16.330 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2359.025 16.065 2359.195 18.955 ;
      LAYER mcon ;
        RECT 2359.025 18.785 2359.195 18.955 ;
      LAYER met1 ;
        RECT 2269.250 18.940 2269.570 19.000 ;
        RECT 2358.965 18.940 2359.255 18.985 ;
        RECT 2269.250 18.800 2359.255 18.940 ;
        RECT 2269.250 18.740 2269.570 18.800 ;
        RECT 2358.965 18.755 2359.255 18.800 ;
        RECT 2393.450 16.560 2393.770 16.620 ;
        RECT 2376.060 16.420 2393.770 16.560 ;
        RECT 2358.965 16.220 2359.255 16.265 ;
        RECT 2376.060 16.220 2376.200 16.420 ;
        RECT 2393.450 16.360 2393.770 16.420 ;
        RECT 2358.965 16.080 2376.200 16.220 ;
        RECT 2358.965 16.035 2359.255 16.080 ;
      LAYER via ;
        RECT 2269.280 18.740 2269.540 19.000 ;
        RECT 2393.480 16.360 2393.740 16.620 ;
      LAYER met2 ;
        RECT 2268.820 300.290 2269.100 304.000 ;
        RECT 2268.820 300.150 2269.480 300.290 ;
        RECT 2268.820 300.000 2269.100 300.150 ;
        RECT 2269.340 19.030 2269.480 300.150 ;
        RECT 2269.280 18.710 2269.540 19.030 ;
        RECT 2393.480 16.330 2393.740 16.650 ;
        RECT 2393.540 2.400 2393.680 16.330 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2283.540 300.290 2283.820 304.000 ;
        RECT 2283.140 300.150 2283.820 300.290 ;
        RECT 2283.140 16.845 2283.280 300.150 ;
        RECT 2283.540 300.000 2283.820 300.150 ;
        RECT 2283.070 16.475 2283.350 16.845 ;
        RECT 2411.410 16.475 2411.690 16.845 ;
        RECT 2411.480 2.400 2411.620 16.475 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
      LAYER via2 ;
        RECT 2283.070 16.520 2283.350 16.800 ;
        RECT 2411.410 16.520 2411.690 16.800 ;
      LAYER met3 ;
        RECT 2283.045 16.810 2283.375 16.825 ;
        RECT 2411.385 16.810 2411.715 16.825 ;
        RECT 2283.045 16.510 2411.715 16.810 ;
        RECT 2283.045 16.495 2283.375 16.510 ;
        RECT 2411.385 16.495 2411.715 16.510 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 807.445 17.765 807.615 19.975 ;
        RECT 845.625 17.765 845.795 19.635 ;
      LAYER mcon ;
        RECT 807.445 19.805 807.615 19.975 ;
        RECT 845.625 19.465 845.795 19.635 ;
      LAYER met1 ;
        RECT 865.790 283.120 866.110 283.180 ;
        RECT 961.010 283.120 961.330 283.180 ;
        RECT 865.790 282.980 961.330 283.120 ;
        RECT 865.790 282.920 866.110 282.980 ;
        RECT 961.010 282.920 961.330 282.980 ;
        RECT 805.530 19.960 805.850 20.020 ;
        RECT 807.385 19.960 807.675 20.005 ;
        RECT 805.530 19.820 807.675 19.960 ;
        RECT 805.530 19.760 805.850 19.820 ;
        RECT 807.385 19.775 807.675 19.820 ;
        RECT 845.565 19.620 845.855 19.665 ;
        RECT 865.790 19.620 866.110 19.680 ;
        RECT 845.565 19.480 866.110 19.620 ;
        RECT 845.565 19.435 845.855 19.480 ;
        RECT 865.790 19.420 866.110 19.480 ;
        RECT 807.385 17.920 807.675 17.965 ;
        RECT 845.565 17.920 845.855 17.965 ;
        RECT 807.385 17.780 845.855 17.920 ;
        RECT 807.385 17.735 807.675 17.780 ;
        RECT 845.565 17.735 845.855 17.780 ;
      LAYER via ;
        RECT 865.820 282.920 866.080 283.180 ;
        RECT 961.040 282.920 961.300 283.180 ;
        RECT 805.560 19.760 805.820 20.020 ;
        RECT 865.820 19.420 866.080 19.680 ;
      LAYER met2 ;
        RECT 961.040 300.000 961.320 304.000 ;
        RECT 961.100 283.210 961.240 300.000 ;
        RECT 865.820 282.890 866.080 283.210 ;
        RECT 961.040 282.890 961.300 283.210 ;
        RECT 805.560 19.730 805.820 20.050 ;
        RECT 805.620 2.400 805.760 19.730 ;
        RECT 865.880 19.710 866.020 282.890 ;
        RECT 865.820 19.390 866.080 19.710 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 24.380 3.150 24.440 ;
        RECT 296.770 24.380 297.090 24.440 ;
        RECT 2.830 24.240 297.090 24.380 ;
        RECT 2.830 24.180 3.150 24.240 ;
        RECT 296.770 24.180 297.090 24.240 ;
      LAYER via ;
        RECT 2.860 24.180 3.120 24.440 ;
        RECT 296.800 24.180 297.060 24.440 ;
      LAYER met2 ;
        RECT 300.020 300.290 300.300 304.000 ;
        RECT 296.860 300.150 300.300 300.290 ;
        RECT 296.860 24.470 297.000 300.150 ;
        RECT 300.020 300.000 300.300 300.150 ;
        RECT 2.860 24.150 3.120 24.470 ;
        RECT 296.800 24.150 297.060 24.470 ;
        RECT 2.920 2.400 3.060 24.150 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 24.040 8.670 24.100 ;
        RECT 304.130 24.040 304.450 24.100 ;
        RECT 8.350 23.900 304.450 24.040 ;
        RECT 8.350 23.840 8.670 23.900 ;
        RECT 304.130 23.840 304.450 23.900 ;
      LAYER via ;
        RECT 8.380 23.840 8.640 24.100 ;
        RECT 304.160 23.840 304.420 24.100 ;
      LAYER met2 ;
        RECT 304.620 300.290 304.900 304.000 ;
        RECT 304.220 300.150 304.900 300.290 ;
        RECT 304.220 24.130 304.360 300.150 ;
        RECT 304.620 300.000 304.900 300.150 ;
        RECT 8.380 23.810 8.640 24.130 ;
        RECT 304.160 23.810 304.420 24.130 ;
        RECT 8.440 2.400 8.580 23.810 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 303.670 289.920 303.990 289.980 ;
        RECT 308.270 289.920 308.590 289.980 ;
        RECT 303.670 289.780 308.590 289.920 ;
        RECT 303.670 289.720 303.990 289.780 ;
        RECT 308.270 289.720 308.590 289.780 ;
        RECT 14.330 25.060 14.650 25.120 ;
        RECT 303.670 25.060 303.990 25.120 ;
        RECT 14.330 24.920 303.990 25.060 ;
        RECT 14.330 24.860 14.650 24.920 ;
        RECT 303.670 24.860 303.990 24.920 ;
      LAYER via ;
        RECT 303.700 289.720 303.960 289.980 ;
        RECT 308.300 289.720 308.560 289.980 ;
        RECT 14.360 24.860 14.620 25.120 ;
        RECT 303.700 24.860 303.960 25.120 ;
      LAYER met2 ;
        RECT 309.680 300.290 309.960 304.000 ;
        RECT 308.360 300.150 309.960 300.290 ;
        RECT 308.360 290.010 308.500 300.150 ;
        RECT 309.680 300.000 309.960 300.150 ;
        RECT 303.700 289.690 303.960 290.010 ;
        RECT 308.300 289.690 308.560 290.010 ;
        RECT 303.760 25.150 303.900 289.690 ;
        RECT 14.360 24.830 14.620 25.150 ;
        RECT 303.700 24.830 303.960 25.150 ;
        RECT 14.420 2.400 14.560 24.830 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 324.830 286.860 325.150 286.920 ;
        RECT 327.590 286.860 327.910 286.920 ;
        RECT 324.830 286.720 327.910 286.860 ;
        RECT 324.830 286.660 325.150 286.720 ;
        RECT 327.590 286.660 327.910 286.720 ;
        RECT 38.250 24.720 38.570 24.780 ;
        RECT 324.830 24.720 325.150 24.780 ;
        RECT 38.250 24.580 325.150 24.720 ;
        RECT 38.250 24.520 38.570 24.580 ;
        RECT 324.830 24.520 325.150 24.580 ;
      LAYER via ;
        RECT 324.860 286.660 325.120 286.920 ;
        RECT 327.620 286.660 327.880 286.920 ;
        RECT 38.280 24.520 38.540 24.780 ;
        RECT 324.860 24.520 325.120 24.780 ;
      LAYER met2 ;
        RECT 329.000 300.290 329.280 304.000 ;
        RECT 327.680 300.150 329.280 300.290 ;
        RECT 327.680 286.950 327.820 300.150 ;
        RECT 329.000 300.000 329.280 300.150 ;
        RECT 324.860 286.630 325.120 286.950 ;
        RECT 327.620 286.630 327.880 286.950 ;
        RECT 324.920 24.810 325.060 286.630 ;
        RECT 38.280 24.490 38.540 24.810 ;
        RECT 324.860 24.490 325.120 24.810 ;
        RECT 38.340 2.400 38.480 24.490 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 492.805 234.685 492.975 241.655 ;
      LAYER mcon ;
        RECT 492.805 241.485 492.975 241.655 ;
      LAYER met1 ;
        RECT 492.730 241.640 493.050 241.700 ;
        RECT 492.535 241.500 493.050 241.640 ;
        RECT 492.730 241.440 493.050 241.500 ;
        RECT 492.730 234.840 493.050 234.900 ;
        RECT 492.535 234.700 493.050 234.840 ;
        RECT 492.730 234.640 493.050 234.700 ;
        RECT 491.350 189.960 491.670 190.020 ;
        RECT 492.270 189.960 492.590 190.020 ;
        RECT 491.350 189.820 492.590 189.960 ;
        RECT 491.350 189.760 491.670 189.820 ;
        RECT 492.270 189.760 492.590 189.820 ;
        RECT 489.970 144.740 490.290 144.800 ;
        RECT 492.270 144.740 492.590 144.800 ;
        RECT 489.970 144.600 492.590 144.740 ;
        RECT 489.970 144.540 490.290 144.600 ;
        RECT 492.270 144.540 492.590 144.600 ;
        RECT 240.650 26.760 240.970 26.820 ;
        RECT 490.890 26.760 491.210 26.820 ;
        RECT 240.650 26.620 491.210 26.760 ;
        RECT 240.650 26.560 240.970 26.620 ;
        RECT 490.890 26.560 491.210 26.620 ;
      LAYER via ;
        RECT 492.760 241.440 493.020 241.700 ;
        RECT 492.760 234.640 493.020 234.900 ;
        RECT 491.380 189.760 491.640 190.020 ;
        RECT 492.300 189.760 492.560 190.020 ;
        RECT 490.000 144.540 490.260 144.800 ;
        RECT 492.300 144.540 492.560 144.800 ;
        RECT 240.680 26.560 240.940 26.820 ;
        RECT 490.920 26.560 491.180 26.820 ;
      LAYER met2 ;
        RECT 495.520 300.000 495.800 304.000 ;
        RECT 495.580 290.885 495.720 300.000 ;
        RECT 495.510 290.515 495.790 290.885 ;
        RECT 492.290 290.090 492.570 290.205 ;
        RECT 492.290 289.950 492.960 290.090 ;
        RECT 492.290 289.835 492.570 289.950 ;
        RECT 492.820 241.730 492.960 289.950 ;
        RECT 492.760 241.410 493.020 241.730 ;
        RECT 492.760 234.610 493.020 234.930 ;
        RECT 492.820 234.330 492.960 234.610 ;
        RECT 492.360 234.190 492.960 234.330 ;
        RECT 492.360 190.050 492.500 234.190 ;
        RECT 491.380 189.730 491.640 190.050 ;
        RECT 492.300 189.730 492.560 190.050 ;
        RECT 491.440 145.365 491.580 189.730 ;
        RECT 491.370 144.995 491.650 145.365 ;
        RECT 492.290 144.995 492.570 145.365 ;
        RECT 492.360 144.830 492.500 144.995 ;
        RECT 490.000 144.510 490.260 144.830 ;
        RECT 492.300 144.510 492.560 144.830 ;
        RECT 490.060 62.290 490.200 144.510 ;
        RECT 490.060 62.150 491.120 62.290 ;
        RECT 490.980 26.850 491.120 62.150 ;
        RECT 240.680 26.530 240.940 26.850 ;
        RECT 490.920 26.530 491.180 26.850 ;
        RECT 240.740 2.400 240.880 26.530 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 495.510 290.560 495.790 290.840 ;
        RECT 492.290 289.880 492.570 290.160 ;
        RECT 491.370 145.040 491.650 145.320 ;
        RECT 492.290 145.040 492.570 145.320 ;
      LAYER met3 ;
        RECT 495.485 290.850 495.815 290.865 ;
        RECT 491.590 290.550 495.815 290.850 ;
        RECT 491.590 290.170 491.890 290.550 ;
        RECT 495.485 290.535 495.815 290.550 ;
        RECT 492.265 290.170 492.595 290.185 ;
        RECT 491.590 289.870 492.595 290.170 ;
        RECT 492.265 289.855 492.595 289.870 ;
        RECT 491.345 145.330 491.675 145.345 ;
        RECT 492.265 145.330 492.595 145.345 ;
        RECT 491.345 145.030 492.595 145.330 ;
        RECT 491.345 145.015 491.675 145.030 ;
        RECT 492.265 145.015 492.595 145.030 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 504.305 241.485 504.475 261.715 ;
        RECT 505.225 158.185 505.395 193.035 ;
      LAYER mcon ;
        RECT 504.305 261.545 504.475 261.715 ;
        RECT 505.225 192.865 505.395 193.035 ;
      LAYER met1 ;
        RECT 504.245 261.700 504.535 261.745 ;
        RECT 506.070 261.700 506.390 261.760 ;
        RECT 504.245 261.560 506.390 261.700 ;
        RECT 504.245 261.515 504.535 261.560 ;
        RECT 506.070 261.500 506.390 261.560 ;
        RECT 504.230 241.640 504.550 241.700 ;
        RECT 504.035 241.500 504.550 241.640 ;
        RECT 504.230 241.440 504.550 241.500 ;
        RECT 505.150 193.020 505.470 193.080 ;
        RECT 504.955 192.880 505.470 193.020 ;
        RECT 505.150 192.820 505.470 192.880 ;
        RECT 505.165 158.340 505.455 158.385 ;
        RECT 506.070 158.340 506.390 158.400 ;
        RECT 505.165 158.200 506.390 158.340 ;
        RECT 505.165 158.155 505.455 158.200 ;
        RECT 506.070 158.140 506.390 158.200 ;
        RECT 503.770 144.740 504.090 144.800 ;
        RECT 506.070 144.740 506.390 144.800 ;
        RECT 503.770 144.600 506.390 144.740 ;
        RECT 503.770 144.540 504.090 144.600 ;
        RECT 506.070 144.540 506.390 144.600 ;
        RECT 258.130 27.440 258.450 27.500 ;
        RECT 504.690 27.440 505.010 27.500 ;
        RECT 258.130 27.300 505.010 27.440 ;
        RECT 258.130 27.240 258.450 27.300 ;
        RECT 504.690 27.240 505.010 27.300 ;
      LAYER via ;
        RECT 506.100 261.500 506.360 261.760 ;
        RECT 504.260 241.440 504.520 241.700 ;
        RECT 505.180 192.820 505.440 193.080 ;
        RECT 506.100 158.140 506.360 158.400 ;
        RECT 503.800 144.540 504.060 144.800 ;
        RECT 506.100 144.540 506.360 144.800 ;
        RECT 258.160 27.240 258.420 27.500 ;
        RECT 504.720 27.240 504.980 27.500 ;
      LAYER met2 ;
        RECT 510.240 300.970 510.520 304.000 ;
        RECT 506.160 300.830 510.520 300.970 ;
        RECT 506.160 261.790 506.300 300.830 ;
        RECT 510.240 300.000 510.520 300.830 ;
        RECT 506.100 261.470 506.360 261.790 ;
        RECT 504.260 241.410 504.520 241.730 ;
        RECT 504.320 217.330 504.460 241.410 ;
        RECT 504.320 217.190 505.380 217.330 ;
        RECT 505.240 193.110 505.380 217.190 ;
        RECT 505.180 192.790 505.440 193.110 ;
        RECT 506.100 158.110 506.360 158.430 ;
        RECT 506.160 144.830 506.300 158.110 ;
        RECT 503.800 144.510 504.060 144.830 ;
        RECT 506.100 144.510 506.360 144.830 ;
        RECT 503.860 62.290 504.000 144.510 ;
        RECT 503.860 62.150 504.920 62.290 ;
        RECT 504.780 27.530 504.920 62.150 ;
        RECT 258.160 27.210 258.420 27.530 ;
        RECT 504.720 27.210 504.980 27.530 ;
        RECT 258.220 2.400 258.360 27.210 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 276.070 23.700 276.390 23.760 ;
        RECT 524.930 23.700 525.250 23.760 ;
        RECT 276.070 23.560 525.250 23.700 ;
        RECT 276.070 23.500 276.390 23.560 ;
        RECT 524.930 23.500 525.250 23.560 ;
      LAYER via ;
        RECT 276.100 23.500 276.360 23.760 ;
        RECT 524.960 23.500 525.220 23.760 ;
      LAYER met2 ;
        RECT 524.960 300.000 525.240 304.000 ;
        RECT 525.020 23.790 525.160 300.000 ;
        RECT 276.100 23.470 276.360 23.790 ;
        RECT 524.960 23.470 525.220 23.790 ;
        RECT 276.160 2.400 276.300 23.470 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 27.100 294.330 27.160 ;
        RECT 538.730 27.100 539.050 27.160 ;
        RECT 294.010 26.960 539.050 27.100 ;
        RECT 294.010 26.900 294.330 26.960 ;
        RECT 538.730 26.900 539.050 26.960 ;
      LAYER via ;
        RECT 294.040 26.900 294.300 27.160 ;
        RECT 538.760 26.900 539.020 27.160 ;
      LAYER met2 ;
        RECT 539.680 300.290 539.960 304.000 ;
        RECT 538.820 300.150 539.960 300.290 ;
        RECT 538.820 27.190 538.960 300.150 ;
        RECT 539.680 300.000 539.960 300.150 ;
        RECT 294.040 26.870 294.300 27.190 ;
        RECT 538.760 26.870 539.020 27.190 ;
        RECT 294.100 2.400 294.240 26.870 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 24.040 312.270 24.100 ;
        RECT 552.070 24.040 552.390 24.100 ;
        RECT 311.950 23.900 552.390 24.040 ;
        RECT 311.950 23.840 312.270 23.900 ;
        RECT 552.070 23.840 552.390 23.900 ;
      LAYER via ;
        RECT 311.980 23.840 312.240 24.100 ;
        RECT 552.100 23.840 552.360 24.100 ;
      LAYER met2 ;
        RECT 554.400 300.290 554.680 304.000 ;
        RECT 552.160 300.150 554.680 300.290 ;
        RECT 552.160 24.130 552.300 300.150 ;
        RECT 554.400 300.000 554.680 300.150 ;
        RECT 311.980 23.810 312.240 24.130 ;
        RECT 552.100 23.810 552.360 24.130 ;
        RECT 312.040 2.400 312.180 23.810 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 24.380 330.210 24.440 ;
        RECT 565.870 24.380 566.190 24.440 ;
        RECT 329.890 24.240 566.190 24.380 ;
        RECT 329.890 24.180 330.210 24.240 ;
        RECT 565.870 24.180 566.190 24.240 ;
      LAYER via ;
        RECT 329.920 24.180 330.180 24.440 ;
        RECT 565.900 24.180 566.160 24.440 ;
      LAYER met2 ;
        RECT 569.120 300.290 569.400 304.000 ;
        RECT 565.960 300.150 569.400 300.290 ;
        RECT 565.960 24.470 566.100 300.150 ;
        RECT 569.120 300.000 569.400 300.150 ;
        RECT 329.920 24.150 330.180 24.470 ;
        RECT 565.900 24.150 566.160 24.470 ;
        RECT 329.980 2.400 330.120 24.150 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 25.060 347.690 25.120 ;
        RECT 579.670 25.060 579.990 25.120 ;
        RECT 347.370 24.920 579.990 25.060 ;
        RECT 347.370 24.860 347.690 24.920 ;
        RECT 579.670 24.860 579.990 24.920 ;
      LAYER via ;
        RECT 347.400 24.860 347.660 25.120 ;
        RECT 579.700 24.860 579.960 25.120 ;
      LAYER met2 ;
        RECT 583.840 300.290 584.120 304.000 ;
        RECT 579.760 300.150 584.120 300.290 ;
        RECT 579.760 25.150 579.900 300.150 ;
        RECT 583.840 300.000 584.120 300.150 ;
        RECT 347.400 24.830 347.660 25.150 ;
        RECT 579.700 24.830 579.960 25.150 ;
        RECT 347.460 2.400 347.600 24.830 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 24.720 365.630 24.780 ;
        RECT 593.930 24.720 594.250 24.780 ;
        RECT 365.310 24.580 594.250 24.720 ;
        RECT 365.310 24.520 365.630 24.580 ;
        RECT 593.930 24.520 594.250 24.580 ;
      LAYER via ;
        RECT 365.340 24.520 365.600 24.780 ;
        RECT 593.960 24.520 594.220 24.780 ;
      LAYER met2 ;
        RECT 598.560 300.290 598.840 304.000 ;
        RECT 594.020 300.150 598.840 300.290 ;
        RECT 594.020 24.810 594.160 300.150 ;
        RECT 598.560 300.000 598.840 300.150 ;
        RECT 365.340 24.490 365.600 24.810 ;
        RECT 593.960 24.490 594.220 24.810 ;
        RECT 365.400 2.400 365.540 24.490 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 607.805 241.485 607.975 257.975 ;
        RECT 608.265 89.845 608.435 137.955 ;
      LAYER mcon ;
        RECT 607.805 257.805 607.975 257.975 ;
        RECT 608.265 137.785 608.435 137.955 ;
      LAYER met1 ;
        RECT 607.745 257.960 608.035 258.005 ;
        RECT 608.650 257.960 608.970 258.020 ;
        RECT 607.745 257.820 608.970 257.960 ;
        RECT 607.745 257.775 608.035 257.820 ;
        RECT 608.650 257.760 608.970 257.820 ;
        RECT 607.730 241.640 608.050 241.700 ;
        RECT 607.535 241.500 608.050 241.640 ;
        RECT 607.730 241.440 608.050 241.500 ;
        RECT 607.270 206.960 607.590 207.020 ;
        RECT 608.190 206.960 608.510 207.020 ;
        RECT 607.270 206.820 608.510 206.960 ;
        RECT 607.270 206.760 607.590 206.820 ;
        RECT 608.190 206.760 608.510 206.820 ;
        RECT 608.190 158.820 608.510 159.080 ;
        RECT 608.280 158.340 608.420 158.820 ;
        RECT 608.650 158.340 608.970 158.400 ;
        RECT 608.280 158.200 608.970 158.340 ;
        RECT 608.650 158.140 608.970 158.200 ;
        RECT 608.205 137.940 608.495 137.985 ;
        RECT 608.650 137.940 608.970 138.000 ;
        RECT 608.205 137.800 608.970 137.940 ;
        RECT 608.205 137.755 608.495 137.800 ;
        RECT 608.650 137.740 608.970 137.800 ;
        RECT 608.190 90.000 608.510 90.060 ;
        RECT 607.995 89.860 608.510 90.000 ;
        RECT 608.190 89.800 608.510 89.860 ;
        RECT 608.190 62.460 608.510 62.520 ;
        RECT 607.820 62.320 608.510 62.460 ;
        RECT 607.820 62.180 607.960 62.320 ;
        RECT 608.190 62.260 608.510 62.320 ;
        RECT 607.730 61.920 608.050 62.180 ;
        RECT 383.250 26.080 383.570 26.140 ;
        RECT 607.730 26.080 608.050 26.140 ;
        RECT 383.250 25.940 608.050 26.080 ;
        RECT 383.250 25.880 383.570 25.940 ;
        RECT 607.730 25.880 608.050 25.940 ;
      LAYER via ;
        RECT 608.680 257.760 608.940 258.020 ;
        RECT 607.760 241.440 608.020 241.700 ;
        RECT 607.300 206.760 607.560 207.020 ;
        RECT 608.220 206.760 608.480 207.020 ;
        RECT 608.220 158.820 608.480 159.080 ;
        RECT 608.680 158.140 608.940 158.400 ;
        RECT 608.680 137.740 608.940 138.000 ;
        RECT 608.220 89.800 608.480 90.060 ;
        RECT 608.220 62.260 608.480 62.520 ;
        RECT 607.760 61.920 608.020 62.180 ;
        RECT 383.280 25.880 383.540 26.140 ;
        RECT 607.760 25.880 608.020 26.140 ;
      LAYER met2 ;
        RECT 613.280 300.970 613.560 304.000 ;
        RECT 608.740 300.830 613.560 300.970 ;
        RECT 608.740 258.050 608.880 300.830 ;
        RECT 613.280 300.000 613.560 300.830 ;
        RECT 608.680 257.730 608.940 258.050 ;
        RECT 607.760 241.410 608.020 241.730 ;
        RECT 607.820 207.130 607.960 241.410 ;
        RECT 607.360 207.050 607.960 207.130 ;
        RECT 607.300 206.990 607.960 207.050 ;
        RECT 607.300 206.730 607.560 206.990 ;
        RECT 608.220 206.730 608.480 207.050 ;
        RECT 608.280 159.110 608.420 206.730 ;
        RECT 608.220 158.790 608.480 159.110 ;
        RECT 608.680 158.110 608.940 158.430 ;
        RECT 608.740 138.030 608.880 158.110 ;
        RECT 608.680 137.710 608.940 138.030 ;
        RECT 608.220 89.770 608.480 90.090 ;
        RECT 608.280 62.550 608.420 89.770 ;
        RECT 608.220 62.230 608.480 62.550 ;
        RECT 607.760 61.890 608.020 62.210 ;
        RECT 607.820 26.170 607.960 61.890 ;
        RECT 383.280 25.850 383.540 26.170 ;
        RECT 607.760 25.850 608.020 26.170 ;
        RECT 383.340 2.400 383.480 25.850 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 25.740 401.510 25.800 ;
        RECT 627.970 25.740 628.290 25.800 ;
        RECT 401.190 25.600 628.290 25.740 ;
        RECT 401.190 25.540 401.510 25.600 ;
        RECT 627.970 25.540 628.290 25.600 ;
      LAYER via ;
        RECT 401.220 25.540 401.480 25.800 ;
        RECT 628.000 25.540 628.260 25.800 ;
      LAYER met2 ;
        RECT 628.000 300.000 628.280 304.000 ;
        RECT 628.060 25.830 628.200 300.000 ;
        RECT 401.220 25.510 401.480 25.830 ;
        RECT 628.000 25.510 628.260 25.830 ;
        RECT 401.280 2.400 401.420 25.510 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 62.170 26.080 62.490 26.140 ;
        RECT 345.070 26.080 345.390 26.140 ;
        RECT 62.170 25.940 345.390 26.080 ;
        RECT 62.170 25.880 62.490 25.940 ;
        RECT 345.070 25.880 345.390 25.940 ;
      LAYER via ;
        RECT 62.200 25.880 62.460 26.140 ;
        RECT 345.100 25.880 345.360 26.140 ;
      LAYER met2 ;
        RECT 348.780 300.290 349.060 304.000 ;
        RECT 345.160 300.150 349.060 300.290 ;
        RECT 345.160 26.170 345.300 300.150 ;
        RECT 348.780 300.000 349.060 300.150 ;
        RECT 62.200 25.850 62.460 26.170 ;
        RECT 345.100 25.850 345.360 26.170 ;
        RECT 62.260 2.400 62.400 25.850 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 25.400 419.450 25.460 ;
        RECT 642.230 25.400 642.550 25.460 ;
        RECT 419.130 25.260 642.550 25.400 ;
        RECT 419.130 25.200 419.450 25.260 ;
        RECT 642.230 25.200 642.550 25.260 ;
      LAYER via ;
        RECT 419.160 25.200 419.420 25.460 ;
        RECT 642.260 25.200 642.520 25.460 ;
      LAYER met2 ;
        RECT 642.720 300.290 643.000 304.000 ;
        RECT 642.320 300.150 643.000 300.290 ;
        RECT 642.320 25.490 642.460 300.150 ;
        RECT 642.720 300.000 643.000 300.150 ;
        RECT 419.160 25.170 419.420 25.490 ;
        RECT 642.260 25.170 642.520 25.490 ;
        RECT 419.220 2.400 419.360 25.170 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 30.840 436.930 30.900 ;
        RECT 656.030 30.840 656.350 30.900 ;
        RECT 436.610 30.700 656.350 30.840 ;
        RECT 436.610 30.640 436.930 30.700 ;
        RECT 656.030 30.640 656.350 30.700 ;
      LAYER via ;
        RECT 436.640 30.640 436.900 30.900 ;
        RECT 656.060 30.640 656.320 30.900 ;
      LAYER met2 ;
        RECT 657.440 300.290 657.720 304.000 ;
        RECT 656.120 300.150 657.720 300.290 ;
        RECT 656.120 30.930 656.260 300.150 ;
        RECT 657.440 300.000 657.720 300.150 ;
        RECT 436.640 30.610 436.900 30.930 ;
        RECT 656.060 30.610 656.320 30.930 ;
        RECT 436.700 2.400 436.840 30.610 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 454.550 26.420 454.870 26.480 ;
        RECT 669.370 26.420 669.690 26.480 ;
        RECT 454.550 26.280 669.690 26.420 ;
        RECT 454.550 26.220 454.870 26.280 ;
        RECT 669.370 26.220 669.690 26.280 ;
      LAYER via ;
        RECT 454.580 26.220 454.840 26.480 ;
        RECT 669.400 26.220 669.660 26.480 ;
      LAYER met2 ;
        RECT 672.160 300.290 672.440 304.000 ;
        RECT 669.460 300.150 672.440 300.290 ;
        RECT 669.460 26.510 669.600 300.150 ;
        RECT 672.160 300.000 672.440 300.150 ;
        RECT 454.580 26.190 454.840 26.510 ;
        RECT 669.400 26.190 669.660 26.510 ;
        RECT 454.640 2.400 454.780 26.190 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.490 31.180 472.810 31.240 ;
        RECT 683.170 31.180 683.490 31.240 ;
        RECT 472.490 31.040 683.490 31.180 ;
        RECT 472.490 30.980 472.810 31.040 ;
        RECT 683.170 30.980 683.490 31.040 ;
      LAYER via ;
        RECT 472.520 30.980 472.780 31.240 ;
        RECT 683.200 30.980 683.460 31.240 ;
      LAYER met2 ;
        RECT 686.880 300.290 687.160 304.000 ;
        RECT 683.260 300.150 687.160 300.290 ;
        RECT 683.260 31.270 683.400 300.150 ;
        RECT 686.880 300.000 687.160 300.150 ;
        RECT 472.520 30.950 472.780 31.270 ;
        RECT 683.200 30.950 683.460 31.270 ;
        RECT 472.580 2.400 472.720 30.950 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 490.430 23.360 490.750 23.420 ;
        RECT 696.970 23.360 697.290 23.420 ;
        RECT 490.430 23.220 697.290 23.360 ;
        RECT 490.430 23.160 490.750 23.220 ;
        RECT 696.970 23.160 697.290 23.220 ;
      LAYER via ;
        RECT 490.460 23.160 490.720 23.420 ;
        RECT 697.000 23.160 697.260 23.420 ;
      LAYER met2 ;
        RECT 701.600 300.290 701.880 304.000 ;
        RECT 697.060 300.150 701.880 300.290 ;
        RECT 697.060 23.450 697.200 300.150 ;
        RECT 701.600 300.000 701.880 300.150 ;
        RECT 490.460 23.130 490.720 23.450 ;
        RECT 697.000 23.130 697.260 23.450 ;
        RECT 490.520 2.400 490.660 23.130 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 26.760 508.230 26.820 ;
        RECT 711.690 26.760 712.010 26.820 ;
        RECT 507.910 26.620 712.010 26.760 ;
        RECT 507.910 26.560 508.230 26.620 ;
        RECT 711.690 26.560 712.010 26.620 ;
      LAYER via ;
        RECT 507.940 26.560 508.200 26.820 ;
        RECT 711.720 26.560 711.980 26.820 ;
      LAYER met2 ;
        RECT 715.860 300.290 716.140 304.000 ;
        RECT 711.780 300.150 716.140 300.290 ;
        RECT 711.780 26.850 711.920 300.150 ;
        RECT 715.860 300.000 716.140 300.150 ;
        RECT 507.940 26.530 508.200 26.850 ;
        RECT 711.720 26.530 711.980 26.850 ;
        RECT 508.000 2.400 508.140 26.530 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 725.105 144.925 725.275 178.755 ;
      LAYER mcon ;
        RECT 725.105 178.585 725.275 178.755 ;
      LAYER met1 ;
        RECT 725.950 241.640 726.270 241.700 ;
        RECT 726.410 241.640 726.730 241.700 ;
        RECT 725.950 241.500 726.730 241.640 ;
        RECT 725.950 241.440 726.270 241.500 ;
        RECT 726.410 241.440 726.730 241.500 ;
        RECT 725.030 193.360 725.350 193.420 ;
        RECT 725.490 193.360 725.810 193.420 ;
        RECT 725.030 193.220 725.810 193.360 ;
        RECT 725.030 193.160 725.350 193.220 ;
        RECT 725.490 193.160 725.810 193.220 ;
        RECT 725.030 178.740 725.350 178.800 ;
        RECT 724.835 178.600 725.350 178.740 ;
        RECT 725.030 178.540 725.350 178.600 ;
        RECT 725.045 145.080 725.335 145.125 ;
        RECT 725.950 145.080 726.270 145.140 ;
        RECT 725.045 144.940 726.270 145.080 ;
        RECT 725.045 144.895 725.335 144.940 ;
        RECT 725.950 144.880 726.270 144.940 ;
        RECT 725.030 96.800 725.350 96.860 ;
        RECT 725.490 96.800 725.810 96.860 ;
        RECT 725.030 96.660 725.810 96.800 ;
        RECT 725.030 96.600 725.350 96.660 ;
        RECT 725.490 96.600 725.810 96.660 ;
        RECT 525.850 27.440 526.170 27.500 ;
        RECT 725.490 27.440 725.810 27.500 ;
        RECT 525.850 27.300 725.810 27.440 ;
        RECT 525.850 27.240 526.170 27.300 ;
        RECT 725.490 27.240 725.810 27.300 ;
      LAYER via ;
        RECT 725.980 241.440 726.240 241.700 ;
        RECT 726.440 241.440 726.700 241.700 ;
        RECT 725.060 193.160 725.320 193.420 ;
        RECT 725.520 193.160 725.780 193.420 ;
        RECT 725.060 178.540 725.320 178.800 ;
        RECT 725.980 144.880 726.240 145.140 ;
        RECT 725.060 96.600 725.320 96.860 ;
        RECT 725.520 96.600 725.780 96.860 ;
        RECT 525.880 27.240 526.140 27.500 ;
        RECT 725.520 27.240 725.780 27.500 ;
      LAYER met2 ;
        RECT 730.580 300.970 730.860 304.000 ;
        RECT 726.500 300.830 730.860 300.970 ;
        RECT 726.500 241.730 726.640 300.830 ;
        RECT 730.580 300.000 730.860 300.830 ;
        RECT 725.980 241.410 726.240 241.730 ;
        RECT 726.440 241.410 726.700 241.730 ;
        RECT 726.040 207.810 726.180 241.410 ;
        RECT 725.580 207.670 726.180 207.810 ;
        RECT 725.580 193.450 725.720 207.670 ;
        RECT 725.060 193.130 725.320 193.450 ;
        RECT 725.520 193.130 725.780 193.450 ;
        RECT 725.120 178.830 725.260 193.130 ;
        RECT 725.060 178.510 725.320 178.830 ;
        RECT 725.980 144.850 726.240 145.170 ;
        RECT 726.040 111.250 726.180 144.850 ;
        RECT 725.580 111.110 726.180 111.250 ;
        RECT 725.580 96.890 725.720 111.110 ;
        RECT 725.060 96.570 725.320 96.890 ;
        RECT 725.520 96.570 725.780 96.890 ;
        RECT 725.120 62.290 725.260 96.570 ;
        RECT 725.120 62.150 725.720 62.290 ;
        RECT 725.580 27.530 725.720 62.150 ;
        RECT 525.880 27.210 526.140 27.530 ;
        RECT 725.520 27.210 725.780 27.530 ;
        RECT 525.940 2.400 526.080 27.210 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 544.710 289.580 545.030 289.640 ;
        RECT 544.710 289.440 560.120 289.580 ;
        RECT 544.710 289.380 545.030 289.440 ;
        RECT 559.980 289.240 560.120 289.440 ;
        RECT 745.270 289.240 745.590 289.300 ;
        RECT 559.980 289.100 745.590 289.240 ;
        RECT 745.270 289.040 745.590 289.100 ;
      LAYER via ;
        RECT 544.740 289.380 545.000 289.640 ;
        RECT 745.300 289.040 745.560 289.300 ;
      LAYER met2 ;
        RECT 745.300 300.000 745.580 304.000 ;
        RECT 544.740 289.350 545.000 289.670 ;
        RECT 544.800 3.130 544.940 289.350 ;
        RECT 745.360 289.330 745.500 300.000 ;
        RECT 745.300 289.010 745.560 289.330 ;
        RECT 543.880 2.990 544.940 3.130 ;
        RECT 543.880 2.400 544.020 2.990 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 565.410 289.580 565.730 289.640 ;
        RECT 759.990 289.580 760.310 289.640 ;
        RECT 565.410 289.440 760.310 289.580 ;
        RECT 565.410 289.380 565.730 289.440 ;
        RECT 759.990 289.380 760.310 289.440 ;
        RECT 561.730 20.640 562.050 20.700 ;
        RECT 565.410 20.640 565.730 20.700 ;
        RECT 561.730 20.500 565.730 20.640 ;
        RECT 561.730 20.440 562.050 20.500 ;
        RECT 565.410 20.440 565.730 20.500 ;
      LAYER via ;
        RECT 565.440 289.380 565.700 289.640 ;
        RECT 760.020 289.380 760.280 289.640 ;
        RECT 561.760 20.440 562.020 20.700 ;
        RECT 565.440 20.440 565.700 20.700 ;
      LAYER met2 ;
        RECT 760.020 300.000 760.300 304.000 ;
        RECT 760.080 289.670 760.220 300.000 ;
        RECT 565.440 289.350 565.700 289.670 ;
        RECT 760.020 289.350 760.280 289.670 ;
        RECT 565.500 20.730 565.640 289.350 ;
        RECT 561.760 20.410 562.020 20.730 ;
        RECT 565.440 20.410 565.700 20.730 ;
        RECT 561.820 2.400 561.960 20.410 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 586.110 285.500 586.430 285.560 ;
        RECT 774.710 285.500 775.030 285.560 ;
        RECT 586.110 285.360 775.030 285.500 ;
        RECT 586.110 285.300 586.430 285.360 ;
        RECT 774.710 285.300 775.030 285.360 ;
        RECT 579.670 18.600 579.990 18.660 ;
        RECT 586.110 18.600 586.430 18.660 ;
        RECT 579.670 18.460 586.430 18.600 ;
        RECT 579.670 18.400 579.990 18.460 ;
        RECT 586.110 18.400 586.430 18.460 ;
      LAYER via ;
        RECT 586.140 285.300 586.400 285.560 ;
        RECT 774.740 285.300 775.000 285.560 ;
        RECT 579.700 18.400 579.960 18.660 ;
        RECT 586.140 18.400 586.400 18.660 ;
      LAYER met2 ;
        RECT 774.740 300.000 775.020 304.000 ;
        RECT 774.800 285.590 774.940 300.000 ;
        RECT 586.140 285.270 586.400 285.590 ;
        RECT 774.740 285.270 775.000 285.590 ;
        RECT 586.200 18.690 586.340 285.270 ;
        RECT 579.700 18.370 579.960 18.690 ;
        RECT 586.140 18.370 586.400 18.690 ;
        RECT 579.760 2.400 579.900 18.370 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 25.400 86.410 25.460 ;
        RECT 365.770 25.400 366.090 25.460 ;
        RECT 86.090 25.260 366.090 25.400 ;
        RECT 86.090 25.200 86.410 25.260 ;
        RECT 365.770 25.200 366.090 25.260 ;
      LAYER via ;
        RECT 86.120 25.200 86.380 25.460 ;
        RECT 365.800 25.200 366.060 25.460 ;
      LAYER met2 ;
        RECT 368.560 300.290 368.840 304.000 ;
        RECT 365.860 300.150 368.840 300.290 ;
        RECT 365.860 25.490 366.000 300.150 ;
        RECT 368.560 300.000 368.840 300.150 ;
        RECT 86.120 25.170 86.380 25.490 ;
        RECT 365.800 25.170 366.060 25.490 ;
        RECT 86.180 2.400 86.320 25.170 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 599.910 285.160 600.230 285.220 ;
        RECT 789.430 285.160 789.750 285.220 ;
        RECT 599.910 285.020 789.750 285.160 ;
        RECT 599.910 284.960 600.230 285.020 ;
        RECT 789.430 284.960 789.750 285.020 ;
        RECT 597.150 20.640 597.470 20.700 ;
        RECT 599.910 20.640 600.230 20.700 ;
        RECT 597.150 20.500 600.230 20.640 ;
        RECT 597.150 20.440 597.470 20.500 ;
        RECT 599.910 20.440 600.230 20.500 ;
      LAYER via ;
        RECT 599.940 284.960 600.200 285.220 ;
        RECT 789.460 284.960 789.720 285.220 ;
        RECT 597.180 20.440 597.440 20.700 ;
        RECT 599.940 20.440 600.200 20.700 ;
      LAYER met2 ;
        RECT 789.460 300.000 789.740 304.000 ;
        RECT 789.520 285.250 789.660 300.000 ;
        RECT 599.940 284.930 600.200 285.250 ;
        RECT 789.460 284.930 789.720 285.250 ;
        RECT 600.000 20.730 600.140 284.930 ;
        RECT 597.180 20.410 597.440 20.730 ;
        RECT 599.940 20.410 600.200 20.730 ;
        RECT 597.240 2.400 597.380 20.410 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 661.165 286.025 661.335 287.215 ;
      LAYER mcon ;
        RECT 661.165 287.045 661.335 287.215 ;
      LAYER met1 ;
        RECT 620.610 287.200 620.930 287.260 ;
        RECT 661.105 287.200 661.395 287.245 ;
        RECT 620.610 287.060 661.395 287.200 ;
        RECT 620.610 287.000 620.930 287.060 ;
        RECT 661.105 287.015 661.395 287.060 ;
        RECT 661.105 286.180 661.395 286.225 ;
        RECT 804.150 286.180 804.470 286.240 ;
        RECT 661.105 286.040 804.470 286.180 ;
        RECT 661.105 285.995 661.395 286.040 ;
        RECT 804.150 285.980 804.470 286.040 ;
        RECT 615.090 20.640 615.410 20.700 ;
        RECT 620.610 20.640 620.930 20.700 ;
        RECT 615.090 20.500 620.930 20.640 ;
        RECT 615.090 20.440 615.410 20.500 ;
        RECT 620.610 20.440 620.930 20.500 ;
      LAYER via ;
        RECT 620.640 287.000 620.900 287.260 ;
        RECT 804.180 285.980 804.440 286.240 ;
        RECT 615.120 20.440 615.380 20.700 ;
        RECT 620.640 20.440 620.900 20.700 ;
      LAYER met2 ;
        RECT 804.180 300.000 804.460 304.000 ;
        RECT 620.640 286.970 620.900 287.290 ;
        RECT 620.700 20.730 620.840 286.970 ;
        RECT 804.240 286.270 804.380 300.000 ;
        RECT 804.180 285.950 804.440 286.270 ;
        RECT 615.120 20.410 615.380 20.730 ;
        RECT 620.640 20.410 620.900 20.730 ;
        RECT 615.180 2.400 615.320 20.410 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 110.010 25.740 110.330 25.800 ;
        RECT 386.930 25.740 387.250 25.800 ;
        RECT 110.010 25.600 387.250 25.740 ;
        RECT 110.010 25.540 110.330 25.600 ;
        RECT 386.930 25.540 387.250 25.600 ;
      LAYER via ;
        RECT 110.040 25.540 110.300 25.800 ;
        RECT 386.960 25.540 387.220 25.800 ;
      LAYER met2 ;
        RECT 387.880 300.290 388.160 304.000 ;
        RECT 387.020 300.150 388.160 300.290 ;
        RECT 387.020 25.830 387.160 300.150 ;
        RECT 387.880 300.000 388.160 300.150 ;
        RECT 110.040 25.510 110.300 25.830 ;
        RECT 386.960 25.510 387.220 25.830 ;
        RECT 110.100 13.330 110.240 25.510 ;
        RECT 109.640 13.190 110.240 13.330 ;
        RECT 109.640 2.400 109.780 13.190 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 390.150 288.220 390.470 288.280 ;
        RECT 407.630 288.220 407.950 288.280 ;
        RECT 390.150 288.080 407.950 288.220 ;
        RECT 390.150 288.020 390.470 288.080 ;
        RECT 407.630 288.020 407.950 288.080 ;
        RECT 388.770 16.900 389.090 16.960 ;
        RECT 151.960 16.760 389.090 16.900 ;
        RECT 133.470 16.220 133.790 16.280 ;
        RECT 151.960 16.220 152.100 16.760 ;
        RECT 388.770 16.700 389.090 16.760 ;
        RECT 133.470 16.080 152.100 16.220 ;
        RECT 133.470 16.020 133.790 16.080 ;
      LAYER via ;
        RECT 390.180 288.020 390.440 288.280 ;
        RECT 407.660 288.020 407.920 288.280 ;
        RECT 133.500 16.020 133.760 16.280 ;
        RECT 388.800 16.700 389.060 16.960 ;
      LAYER met2 ;
        RECT 407.660 300.000 407.940 304.000 ;
        RECT 407.720 288.310 407.860 300.000 ;
        RECT 390.180 287.990 390.440 288.310 ;
        RECT 407.660 287.990 407.920 288.310 ;
        RECT 390.240 17.410 390.380 287.990 ;
        RECT 388.860 17.270 390.380 17.410 ;
        RECT 388.860 16.990 389.000 17.270 ;
        RECT 388.800 16.670 389.060 16.990 ;
        RECT 133.500 15.990 133.760 16.310 ;
        RECT 133.560 2.400 133.700 15.990 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 26.420 151.730 26.480 ;
        RECT 421.430 26.420 421.750 26.480 ;
        RECT 151.410 26.280 421.750 26.420 ;
        RECT 151.410 26.220 151.730 26.280 ;
        RECT 421.430 26.220 421.750 26.280 ;
      LAYER via ;
        RECT 151.440 26.220 151.700 26.480 ;
        RECT 421.460 26.220 421.720 26.480 ;
      LAYER met2 ;
        RECT 422.380 300.290 422.660 304.000 ;
        RECT 421.520 300.150 422.660 300.290 ;
        RECT 421.520 26.510 421.660 300.150 ;
        RECT 422.380 300.000 422.660 300.150 ;
        RECT 151.440 26.190 151.700 26.510 ;
        RECT 421.460 26.190 421.720 26.510 ;
        RECT 151.500 2.400 151.640 26.190 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 169.350 19.620 169.670 19.680 ;
        RECT 434.770 19.620 435.090 19.680 ;
        RECT 169.350 19.480 435.090 19.620 ;
        RECT 169.350 19.420 169.670 19.480 ;
        RECT 434.770 19.420 435.090 19.480 ;
      LAYER via ;
        RECT 169.380 19.420 169.640 19.680 ;
        RECT 434.800 19.420 435.060 19.680 ;
      LAYER met2 ;
        RECT 437.100 300.290 437.380 304.000 ;
        RECT 434.860 300.150 437.380 300.290 ;
        RECT 434.860 19.710 435.000 300.150 ;
        RECT 437.100 300.000 437.380 300.150 ;
        RECT 169.380 19.390 169.640 19.710 ;
        RECT 434.800 19.390 435.060 19.710 ;
        RECT 169.440 2.400 169.580 19.390 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.350 288.900 192.670 288.960 ;
        RECT 451.790 288.900 452.110 288.960 ;
        RECT 192.350 288.760 452.110 288.900 ;
        RECT 192.350 288.700 192.670 288.760 ;
        RECT 451.790 288.700 452.110 288.760 ;
        RECT 186.830 16.560 187.150 16.620 ;
        RECT 192.350 16.560 192.670 16.620 ;
        RECT 186.830 16.420 192.670 16.560 ;
        RECT 186.830 16.360 187.150 16.420 ;
        RECT 192.350 16.360 192.670 16.420 ;
      LAYER via ;
        RECT 192.380 288.700 192.640 288.960 ;
        RECT 451.820 288.700 452.080 288.960 ;
        RECT 186.860 16.360 187.120 16.620 ;
        RECT 192.380 16.360 192.640 16.620 ;
      LAYER met2 ;
        RECT 451.820 300.000 452.100 304.000 ;
        RECT 451.880 288.990 452.020 300.000 ;
        RECT 192.380 288.670 192.640 288.990 ;
        RECT 451.820 288.670 452.080 288.990 ;
        RECT 192.440 16.650 192.580 288.670 ;
        RECT 186.860 16.330 187.120 16.650 ;
        RECT 192.380 16.330 192.640 16.650 ;
        RECT 186.920 2.400 187.060 16.330 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 206.610 289.240 206.930 289.300 ;
        RECT 466.050 289.240 466.370 289.300 ;
        RECT 206.610 289.100 466.370 289.240 ;
        RECT 206.610 289.040 206.930 289.100 ;
        RECT 466.050 289.040 466.370 289.100 ;
      LAYER via ;
        RECT 206.640 289.040 206.900 289.300 ;
        RECT 466.080 289.040 466.340 289.300 ;
      LAYER met2 ;
        RECT 466.080 300.000 466.360 304.000 ;
        RECT 466.140 289.330 466.280 300.000 ;
        RECT 206.640 289.010 206.900 289.330 ;
        RECT 466.080 289.010 466.340 289.330 ;
        RECT 206.700 17.410 206.840 289.010 ;
        RECT 204.860 17.270 206.840 17.410 ;
        RECT 204.860 2.400 205.000 17.270 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 227.310 285.500 227.630 285.560 ;
        RECT 480.770 285.500 481.090 285.560 ;
        RECT 227.310 285.360 481.090 285.500 ;
        RECT 227.310 285.300 227.630 285.360 ;
        RECT 480.770 285.300 481.090 285.360 ;
        RECT 222.710 16.220 223.030 16.280 ;
        RECT 227.310 16.220 227.630 16.280 ;
        RECT 222.710 16.080 227.630 16.220 ;
        RECT 222.710 16.020 223.030 16.080 ;
        RECT 227.310 16.020 227.630 16.080 ;
      LAYER via ;
        RECT 227.340 285.300 227.600 285.560 ;
        RECT 480.800 285.300 481.060 285.560 ;
        RECT 222.740 16.020 223.000 16.280 ;
        RECT 227.340 16.020 227.600 16.280 ;
      LAYER met2 ;
        RECT 480.800 300.000 481.080 304.000 ;
        RECT 480.860 285.590 481.000 300.000 ;
        RECT 227.340 285.270 227.600 285.590 ;
        RECT 480.800 285.270 481.060 285.590 ;
        RECT 227.400 16.310 227.540 285.270 ;
        RECT 222.740 15.990 223.000 16.310 ;
        RECT 227.340 15.990 227.600 16.310 ;
        RECT 222.800 2.400 222.940 15.990 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 299.605 17.425 299.775 20.995 ;
      LAYER mcon ;
        RECT 299.605 20.825 299.775 20.995 ;
      LAYER met1 ;
        RECT 306.890 284.480 307.210 284.540 ;
        RECT 314.250 284.480 314.570 284.540 ;
        RECT 306.890 284.340 314.570 284.480 ;
        RECT 306.890 284.280 307.210 284.340 ;
        RECT 314.250 284.280 314.570 284.340 ;
        RECT 299.545 20.980 299.835 21.025 ;
        RECT 306.890 20.980 307.210 21.040 ;
        RECT 299.545 20.840 307.210 20.980 ;
        RECT 299.545 20.795 299.835 20.840 ;
        RECT 306.890 20.780 307.210 20.840 ;
        RECT 20.310 17.580 20.630 17.640 ;
        RECT 299.545 17.580 299.835 17.625 ;
        RECT 20.310 17.440 299.835 17.580 ;
        RECT 20.310 17.380 20.630 17.440 ;
        RECT 299.545 17.395 299.835 17.440 ;
      LAYER via ;
        RECT 306.920 284.280 307.180 284.540 ;
        RECT 314.280 284.280 314.540 284.540 ;
        RECT 306.920 20.780 307.180 21.040 ;
        RECT 20.340 17.380 20.600 17.640 ;
      LAYER met2 ;
        RECT 314.280 300.000 314.560 304.000 ;
        RECT 314.340 284.570 314.480 300.000 ;
        RECT 306.920 284.250 307.180 284.570 ;
        RECT 314.280 284.250 314.540 284.570 ;
        RECT 306.980 21.070 307.120 284.250 ;
        RECT 306.920 20.750 307.180 21.070 ;
        RECT 20.340 17.350 20.600 17.670 ;
        RECT 20.400 2.400 20.540 17.350 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 307.350 283.460 307.670 283.520 ;
        RECT 334.030 283.460 334.350 283.520 ;
        RECT 307.350 283.320 334.350 283.460 ;
        RECT 307.350 283.260 307.670 283.320 ;
        RECT 334.030 283.260 334.350 283.320 ;
        RECT 44.230 19.960 44.550 20.020 ;
        RECT 307.350 19.960 307.670 20.020 ;
        RECT 44.230 19.820 307.670 19.960 ;
        RECT 44.230 19.760 44.550 19.820 ;
        RECT 307.350 19.760 307.670 19.820 ;
      LAYER via ;
        RECT 307.380 283.260 307.640 283.520 ;
        RECT 334.060 283.260 334.320 283.520 ;
        RECT 44.260 19.760 44.520 20.020 ;
        RECT 307.380 19.760 307.640 20.020 ;
      LAYER met2 ;
        RECT 334.060 300.000 334.340 304.000 ;
        RECT 334.120 283.550 334.260 300.000 ;
        RECT 307.380 283.230 307.640 283.550 ;
        RECT 334.060 283.230 334.320 283.550 ;
        RECT 307.440 20.050 307.580 283.230 ;
        RECT 44.260 19.730 44.520 20.050 ;
        RECT 307.380 19.730 307.640 20.050 ;
        RECT 44.320 2.400 44.460 19.730 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 493.190 241.300 493.510 241.360 ;
        RECT 500.550 241.300 500.870 241.360 ;
        RECT 493.190 241.160 500.870 241.300 ;
        RECT 493.190 241.100 493.510 241.160 ;
        RECT 500.550 241.100 500.870 241.160 ;
        RECT 493.190 16.560 493.510 16.620 ;
        RECT 269.260 16.420 493.510 16.560 ;
        RECT 246.630 16.220 246.950 16.280 ;
        RECT 269.260 16.220 269.400 16.420 ;
        RECT 493.190 16.360 493.510 16.420 ;
        RECT 246.630 16.080 269.400 16.220 ;
        RECT 246.630 16.020 246.950 16.080 ;
      LAYER via ;
        RECT 493.220 241.100 493.480 241.360 ;
        RECT 500.580 241.100 500.840 241.360 ;
        RECT 246.660 16.020 246.920 16.280 ;
        RECT 493.220 16.360 493.480 16.620 ;
      LAYER met2 ;
        RECT 500.580 300.000 500.860 304.000 ;
        RECT 500.640 241.390 500.780 300.000 ;
        RECT 493.220 241.070 493.480 241.390 ;
        RECT 500.580 241.070 500.840 241.390 ;
        RECT 493.280 16.650 493.420 241.070 ;
        RECT 493.220 16.330 493.480 16.650 ;
        RECT 246.660 15.990 246.920 16.310 ;
        RECT 246.720 2.400 246.860 15.990 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 268.710 284.140 269.030 284.200 ;
        RECT 515.270 284.140 515.590 284.200 ;
        RECT 268.710 284.000 515.590 284.140 ;
        RECT 268.710 283.940 269.030 284.000 ;
        RECT 515.270 283.940 515.590 284.000 ;
        RECT 264.110 16.560 264.430 16.620 ;
        RECT 268.710 16.560 269.030 16.620 ;
        RECT 264.110 16.420 269.030 16.560 ;
        RECT 264.110 16.360 264.430 16.420 ;
        RECT 268.710 16.360 269.030 16.420 ;
      LAYER via ;
        RECT 268.740 283.940 269.000 284.200 ;
        RECT 515.300 283.940 515.560 284.200 ;
        RECT 264.140 16.360 264.400 16.620 ;
        RECT 268.740 16.360 269.000 16.620 ;
      LAYER met2 ;
        RECT 515.300 300.000 515.580 304.000 ;
        RECT 515.360 284.230 515.500 300.000 ;
        RECT 268.740 283.910 269.000 284.230 ;
        RECT 515.300 283.910 515.560 284.230 ;
        RECT 268.800 16.650 268.940 283.910 ;
        RECT 264.140 16.330 264.400 16.650 ;
        RECT 268.740 16.330 269.000 16.650 ;
        RECT 264.200 2.400 264.340 16.330 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 514.350 285.840 514.670 285.900 ;
        RECT 529.990 285.840 530.310 285.900 ;
        RECT 514.350 285.700 530.310 285.840 ;
        RECT 514.350 285.640 514.670 285.700 ;
        RECT 529.990 285.640 530.310 285.700 ;
        RECT 282.050 15.880 282.370 15.940 ;
        RECT 514.350 15.880 514.670 15.940 ;
        RECT 282.050 15.740 514.670 15.880 ;
        RECT 282.050 15.680 282.370 15.740 ;
        RECT 514.350 15.680 514.670 15.740 ;
      LAYER via ;
        RECT 514.380 285.640 514.640 285.900 ;
        RECT 530.020 285.640 530.280 285.900 ;
        RECT 282.080 15.680 282.340 15.940 ;
        RECT 514.380 15.680 514.640 15.940 ;
      LAYER met2 ;
        RECT 530.020 300.000 530.300 304.000 ;
        RECT 530.080 285.930 530.220 300.000 ;
        RECT 514.380 285.610 514.640 285.930 ;
        RECT 530.020 285.610 530.280 285.930 ;
        RECT 514.440 15.970 514.580 285.610 ;
        RECT 282.080 15.650 282.340 15.970 ;
        RECT 514.380 15.650 514.640 15.970 ;
        RECT 282.140 2.400 282.280 15.650 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 513.505 283.305 513.675 284.835 ;
      LAYER mcon ;
        RECT 513.505 284.665 513.675 284.835 ;
      LAYER met1 ;
        RECT 513.445 284.820 513.735 284.865 ;
        RECT 542.870 284.820 543.190 284.880 ;
        RECT 513.445 284.680 543.190 284.820 ;
        RECT 513.445 284.635 513.735 284.680 ;
        RECT 542.870 284.620 543.190 284.680 ;
        RECT 513.445 283.460 513.735 283.505 ;
        RECT 348.380 283.320 513.735 283.460 ;
        RECT 303.210 283.120 303.530 283.180 ;
        RECT 348.380 283.120 348.520 283.320 ;
        RECT 513.445 283.275 513.735 283.320 ;
        RECT 303.210 282.980 348.520 283.120 ;
        RECT 303.210 282.920 303.530 282.980 ;
        RECT 299.990 17.580 300.310 17.640 ;
        RECT 303.210 17.580 303.530 17.640 ;
        RECT 299.990 17.440 303.530 17.580 ;
        RECT 299.990 17.380 300.310 17.440 ;
        RECT 303.210 17.380 303.530 17.440 ;
      LAYER via ;
        RECT 542.900 284.620 543.160 284.880 ;
        RECT 303.240 282.920 303.500 283.180 ;
        RECT 300.020 17.380 300.280 17.640 ;
        RECT 303.240 17.380 303.500 17.640 ;
      LAYER met2 ;
        RECT 544.740 300.290 545.020 304.000 ;
        RECT 542.960 300.150 545.020 300.290 ;
        RECT 542.960 284.910 543.100 300.150 ;
        RECT 544.740 300.000 545.020 300.150 ;
        RECT 542.900 284.590 543.160 284.910 ;
        RECT 303.240 282.890 303.500 283.210 ;
        RECT 303.300 17.670 303.440 282.890 ;
        RECT 300.020 17.350 300.280 17.670 ;
        RECT 303.240 17.350 303.500 17.670 ;
        RECT 300.080 2.400 300.220 17.350 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 520.790 289.240 521.110 289.300 ;
        RECT 559.430 289.240 559.750 289.300 ;
        RECT 520.790 289.100 559.750 289.240 ;
        RECT 520.790 289.040 521.110 289.100 ;
        RECT 559.430 289.040 559.750 289.100 ;
        RECT 317.930 19.960 318.250 20.020 ;
        RECT 520.790 19.960 521.110 20.020 ;
        RECT 317.930 19.820 521.110 19.960 ;
        RECT 317.930 19.760 318.250 19.820 ;
        RECT 520.790 19.760 521.110 19.820 ;
      LAYER via ;
        RECT 520.820 289.040 521.080 289.300 ;
        RECT 559.460 289.040 559.720 289.300 ;
        RECT 317.960 19.760 318.220 20.020 ;
        RECT 520.820 19.760 521.080 20.020 ;
      LAYER met2 ;
        RECT 559.460 300.000 559.740 304.000 ;
        RECT 559.520 289.330 559.660 300.000 ;
        RECT 520.820 289.010 521.080 289.330 ;
        RECT 559.460 289.010 559.720 289.330 ;
        RECT 520.880 20.050 521.020 289.010 ;
        RECT 317.960 19.730 318.220 20.050 ;
        RECT 520.820 19.730 521.080 20.050 ;
        RECT 318.020 2.400 318.160 19.730 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 347.905 283.135 348.075 283.475 ;
        RECT 347.905 282.965 348.995 283.135 ;
        RECT 496.945 282.965 497.115 284.835 ;
        RECT 513.045 283.645 513.215 284.835 ;
      LAYER mcon ;
        RECT 496.945 284.665 497.115 284.835 ;
        RECT 347.905 283.305 348.075 283.475 ;
        RECT 513.045 284.665 513.215 284.835 ;
        RECT 348.825 282.965 348.995 283.135 ;
      LAYER met1 ;
        RECT 496.885 284.820 497.175 284.865 ;
        RECT 512.985 284.820 513.275 284.865 ;
        RECT 496.885 284.680 513.275 284.820 ;
        RECT 496.885 284.635 497.175 284.680 ;
        RECT 512.985 284.635 513.275 284.680 ;
        RECT 512.985 283.800 513.275 283.845 ;
        RECT 512.985 283.660 521.020 283.800 ;
        RECT 512.985 283.615 513.275 283.660 ;
        RECT 337.710 283.460 338.030 283.520 ;
        RECT 347.845 283.460 348.135 283.505 ;
        RECT 337.710 283.320 348.135 283.460 ;
        RECT 520.880 283.460 521.020 283.660 ;
        RECT 574.150 283.460 574.470 283.520 ;
        RECT 520.880 283.320 574.470 283.460 ;
        RECT 337.710 283.260 338.030 283.320 ;
        RECT 347.845 283.275 348.135 283.320 ;
        RECT 574.150 283.260 574.470 283.320 ;
        RECT 348.765 283.120 349.055 283.165 ;
        RECT 496.885 283.120 497.175 283.165 ;
        RECT 348.765 282.980 497.175 283.120 ;
        RECT 348.765 282.935 349.055 282.980 ;
        RECT 496.885 282.935 497.175 282.980 ;
      LAYER via ;
        RECT 337.740 283.260 338.000 283.520 ;
        RECT 574.180 283.260 574.440 283.520 ;
      LAYER met2 ;
        RECT 574.180 300.000 574.460 304.000 ;
        RECT 574.240 283.550 574.380 300.000 ;
        RECT 337.740 283.230 338.000 283.550 ;
        RECT 574.180 283.230 574.440 283.550 ;
        RECT 337.800 3.130 337.940 283.230 ;
        RECT 335.960 2.990 337.940 3.130 ;
        RECT 335.960 2.400 336.100 2.990 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.690 285.160 528.010 285.220 ;
        RECT 588.870 285.160 589.190 285.220 ;
        RECT 527.690 285.020 589.190 285.160 ;
        RECT 527.690 284.960 528.010 285.020 ;
        RECT 588.870 284.960 589.190 285.020 ;
        RECT 353.350 14.860 353.670 14.920 ;
        RECT 527.690 14.860 528.010 14.920 ;
        RECT 353.350 14.720 528.010 14.860 ;
        RECT 353.350 14.660 353.670 14.720 ;
        RECT 527.690 14.660 528.010 14.720 ;
      LAYER via ;
        RECT 527.720 284.960 527.980 285.220 ;
        RECT 588.900 284.960 589.160 285.220 ;
        RECT 353.380 14.660 353.640 14.920 ;
        RECT 527.720 14.660 527.980 14.920 ;
      LAYER met2 ;
        RECT 588.900 300.000 589.180 304.000 ;
        RECT 588.960 285.250 589.100 300.000 ;
        RECT 527.720 284.930 527.980 285.250 ;
        RECT 588.900 284.930 589.160 285.250 ;
        RECT 527.780 14.950 527.920 284.930 ;
        RECT 353.380 14.630 353.640 14.950 ;
        RECT 527.720 14.630 527.980 14.950 ;
        RECT 353.440 2.400 353.580 14.630 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 575.145 283.305 575.315 284.835 ;
        RECT 483.145 20.825 483.775 20.995 ;
        RECT 376.425 18.445 376.595 20.655 ;
        RECT 420.585 18.785 420.755 20.655 ;
        RECT 483.605 20.485 483.775 20.825 ;
        RECT 531.445 20.485 531.615 31.875 ;
      LAYER mcon ;
        RECT 575.145 284.665 575.315 284.835 ;
        RECT 531.445 31.705 531.615 31.875 ;
        RECT 376.425 20.485 376.595 20.655 ;
        RECT 420.585 20.485 420.755 20.655 ;
      LAYER met1 ;
        RECT 555.290 284.820 555.610 284.880 ;
        RECT 575.085 284.820 575.375 284.865 ;
        RECT 555.290 284.680 575.375 284.820 ;
        RECT 555.290 284.620 555.610 284.680 ;
        RECT 575.085 284.635 575.375 284.680 ;
        RECT 575.085 283.460 575.375 283.505 ;
        RECT 603.590 283.460 603.910 283.520 ;
        RECT 575.085 283.320 603.910 283.460 ;
        RECT 575.085 283.275 575.375 283.320 ;
        RECT 603.590 283.260 603.910 283.320 ;
        RECT 531.385 31.860 531.675 31.905 ;
        RECT 555.290 31.860 555.610 31.920 ;
        RECT 531.385 31.720 555.610 31.860 ;
        RECT 531.385 31.675 531.675 31.720 ;
        RECT 555.290 31.660 555.610 31.720 ;
        RECT 483.085 20.980 483.375 21.025 ;
        RECT 372.300 20.840 376.580 20.980 ;
        RECT 371.290 20.640 371.610 20.700 ;
        RECT 372.300 20.640 372.440 20.840 ;
        RECT 376.440 20.685 376.580 20.840 ;
        RECT 466.140 20.840 469.500 20.980 ;
        RECT 371.290 20.500 372.440 20.640 ;
        RECT 371.290 20.440 371.610 20.500 ;
        RECT 376.365 20.455 376.655 20.685 ;
        RECT 420.525 20.640 420.815 20.685 ;
        RECT 466.140 20.640 466.280 20.840 ;
        RECT 420.525 20.500 466.280 20.640 ;
        RECT 469.360 20.640 469.500 20.840 ;
        RECT 478.100 20.840 483.375 20.980 ;
        RECT 478.100 20.640 478.240 20.840 ;
        RECT 483.085 20.795 483.375 20.840 ;
        RECT 469.360 20.500 478.240 20.640 ;
        RECT 483.545 20.640 483.835 20.685 ;
        RECT 531.385 20.640 531.675 20.685 ;
        RECT 483.545 20.500 531.675 20.640 ;
        RECT 420.525 20.455 420.815 20.500 ;
        RECT 483.545 20.455 483.835 20.500 ;
        RECT 531.385 20.455 531.675 20.500 ;
        RECT 420.525 18.940 420.815 18.985 ;
        RECT 400.820 18.800 420.815 18.940 ;
        RECT 376.365 18.600 376.655 18.645 ;
        RECT 400.820 18.600 400.960 18.800 ;
        RECT 420.525 18.755 420.815 18.800 ;
        RECT 376.365 18.460 400.960 18.600 ;
        RECT 376.365 18.415 376.655 18.460 ;
      LAYER via ;
        RECT 555.320 284.620 555.580 284.880 ;
        RECT 603.620 283.260 603.880 283.520 ;
        RECT 555.320 31.660 555.580 31.920 ;
        RECT 371.320 20.440 371.580 20.700 ;
      LAYER met2 ;
        RECT 603.620 300.000 603.900 304.000 ;
        RECT 555.320 284.590 555.580 284.910 ;
        RECT 555.380 31.950 555.520 284.590 ;
        RECT 603.680 283.550 603.820 300.000 ;
        RECT 603.620 283.230 603.880 283.550 ;
        RECT 555.320 31.630 555.580 31.950 ;
        RECT 371.320 20.410 371.580 20.730 ;
        RECT 371.380 2.400 371.520 20.410 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 600.445 285.855 600.615 287.895 ;
        RECT 599.525 285.685 600.615 285.855 ;
        RECT 599.525 285.005 599.695 285.685 ;
        RECT 414.145 16.745 414.315 17.935 ;
      LAYER mcon ;
        RECT 600.445 287.725 600.615 287.895 ;
        RECT 414.145 17.765 414.315 17.935 ;
      LAYER met1 ;
        RECT 600.385 287.880 600.675 287.925 ;
        RECT 612.330 287.880 612.650 287.940 ;
        RECT 600.385 287.740 612.650 287.880 ;
        RECT 600.385 287.695 600.675 287.740 ;
        RECT 612.330 287.680 612.650 287.740 ;
        RECT 589.790 285.160 590.110 285.220 ;
        RECT 599.465 285.160 599.755 285.205 ;
        RECT 589.790 285.020 599.755 285.160 ;
        RECT 589.790 284.960 590.110 285.020 ;
        RECT 599.465 284.975 599.755 285.020 ;
        RECT 414.085 17.920 414.375 17.965 ;
        RECT 589.790 17.920 590.110 17.980 ;
        RECT 414.085 17.780 590.110 17.920 ;
        RECT 414.085 17.735 414.375 17.780 ;
        RECT 589.790 17.720 590.110 17.780 ;
        RECT 389.230 16.900 389.550 16.960 ;
        RECT 414.085 16.900 414.375 16.945 ;
        RECT 389.230 16.760 414.375 16.900 ;
        RECT 389.230 16.700 389.550 16.760 ;
        RECT 414.085 16.715 414.375 16.760 ;
      LAYER via ;
        RECT 612.360 287.680 612.620 287.940 ;
        RECT 589.820 284.960 590.080 285.220 ;
        RECT 589.820 17.720 590.080 17.980 ;
        RECT 389.260 16.700 389.520 16.960 ;
      LAYER met2 ;
        RECT 618.340 300.290 618.620 304.000 ;
        RECT 614.260 300.150 618.620 300.290 ;
        RECT 614.260 288.050 614.400 300.150 ;
        RECT 618.340 300.000 618.620 300.150 ;
        RECT 612.420 287.970 614.400 288.050 ;
        RECT 612.360 287.910 614.400 287.970 ;
        RECT 612.360 287.650 612.620 287.910 ;
        RECT 589.820 284.930 590.080 285.250 ;
        RECT 589.880 18.010 590.020 284.930 ;
        RECT 589.820 17.690 590.080 18.010 ;
        RECT 389.260 16.670 389.520 16.990 ;
        RECT 389.320 2.400 389.460 16.670 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 599.065 286.025 599.235 286.875 ;
      LAYER mcon ;
        RECT 599.065 286.705 599.235 286.875 ;
      LAYER met1 ;
        RECT 413.610 286.860 413.930 286.920 ;
        RECT 599.005 286.860 599.295 286.905 ;
        RECT 630.730 286.860 631.050 286.920 ;
        RECT 413.610 286.720 599.295 286.860 ;
        RECT 413.610 286.660 413.930 286.720 ;
        RECT 599.005 286.675 599.295 286.720 ;
        RECT 623.460 286.720 631.050 286.860 ;
        RECT 599.005 286.180 599.295 286.225 ;
        RECT 623.460 286.180 623.600 286.720 ;
        RECT 630.730 286.660 631.050 286.720 ;
        RECT 599.005 286.040 623.600 286.180 ;
        RECT 599.005 285.995 599.295 286.040 ;
        RECT 407.170 17.920 407.490 17.980 ;
        RECT 413.610 17.920 413.930 17.980 ;
        RECT 407.170 17.780 413.930 17.920 ;
        RECT 407.170 17.720 407.490 17.780 ;
        RECT 413.610 17.720 413.930 17.780 ;
      LAYER via ;
        RECT 413.640 286.660 413.900 286.920 ;
        RECT 630.760 286.660 631.020 286.920 ;
        RECT 407.200 17.720 407.460 17.980 ;
        RECT 413.640 17.720 413.900 17.980 ;
      LAYER met2 ;
        RECT 632.600 300.290 632.880 304.000 ;
        RECT 630.820 300.150 632.880 300.290 ;
        RECT 630.820 286.950 630.960 300.150 ;
        RECT 632.600 300.000 632.880 300.150 ;
        RECT 413.640 286.630 413.900 286.950 ;
        RECT 630.760 286.630 631.020 286.950 ;
        RECT 413.700 18.010 413.840 286.630 ;
        RECT 407.200 17.690 407.460 18.010 ;
        RECT 413.640 17.690 413.900 18.010 ;
        RECT 407.260 2.400 407.400 17.690 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 325.825 286.705 328.295 286.875 ;
        RECT 324.445 285.855 324.615 286.195 ;
        RECT 325.825 285.855 325.995 286.705 ;
        RECT 324.445 285.685 325.995 285.855 ;
      LAYER mcon ;
        RECT 328.125 286.705 328.295 286.875 ;
        RECT 324.445 286.025 324.615 286.195 ;
      LAYER met1 ;
        RECT 328.065 286.860 328.355 286.905 ;
        RECT 353.810 286.860 354.130 286.920 ;
        RECT 328.065 286.720 354.130 286.860 ;
        RECT 328.065 286.675 328.355 286.720 ;
        RECT 353.810 286.660 354.130 286.720 ;
        RECT 68.150 286.180 68.470 286.240 ;
        RECT 324.385 286.180 324.675 286.225 ;
        RECT 68.150 286.040 324.675 286.180 ;
        RECT 68.150 285.980 68.470 286.040 ;
        RECT 324.385 285.995 324.675 286.040 ;
      LAYER via ;
        RECT 353.840 286.660 354.100 286.920 ;
        RECT 68.180 285.980 68.440 286.240 ;
      LAYER met2 ;
        RECT 353.840 300.000 354.120 304.000 ;
        RECT 353.900 286.950 354.040 300.000 ;
        RECT 353.840 286.630 354.100 286.950 ;
        RECT 68.180 285.950 68.440 286.270 ;
        RECT 68.240 2.400 68.380 285.950 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 473.025 287.385 473.195 288.235 ;
      LAYER mcon ;
        RECT 473.025 288.065 473.195 288.235 ;
      LAYER met1 ;
        RECT 427.410 288.220 427.730 288.280 ;
        RECT 472.965 288.220 473.255 288.265 ;
        RECT 427.410 288.080 473.255 288.220 ;
        RECT 427.410 288.020 427.730 288.080 ;
        RECT 472.965 288.035 473.255 288.080 ;
        RECT 472.965 287.540 473.255 287.585 ;
        RECT 647.290 287.540 647.610 287.600 ;
        RECT 472.965 287.400 647.610 287.540 ;
        RECT 472.965 287.355 473.255 287.400 ;
        RECT 647.290 287.340 647.610 287.400 ;
        RECT 424.650 16.900 424.970 16.960 ;
        RECT 427.410 16.900 427.730 16.960 ;
        RECT 424.650 16.760 427.730 16.900 ;
        RECT 424.650 16.700 424.970 16.760 ;
        RECT 427.410 16.700 427.730 16.760 ;
      LAYER via ;
        RECT 427.440 288.020 427.700 288.280 ;
        RECT 647.320 287.340 647.580 287.600 ;
        RECT 424.680 16.700 424.940 16.960 ;
        RECT 427.440 16.700 427.700 16.960 ;
      LAYER met2 ;
        RECT 647.320 300.000 647.600 304.000 ;
        RECT 427.440 287.990 427.700 288.310 ;
        RECT 427.500 16.990 427.640 287.990 ;
        RECT 647.380 287.630 647.520 300.000 ;
        RECT 647.320 287.310 647.580 287.630 ;
        RECT 424.680 16.670 424.940 16.990 ;
        RECT 427.440 16.670 427.700 16.990 ;
        RECT 424.740 2.400 424.880 16.670 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 599.985 286.365 600.155 287.895 ;
        RECT 622.525 286.365 624.075 286.535 ;
        RECT 648.285 286.365 648.455 287.555 ;
      LAYER mcon ;
        RECT 599.985 287.725 600.155 287.895 ;
        RECT 648.285 287.385 648.455 287.555 ;
        RECT 623.905 286.365 624.075 286.535 ;
      LAYER met1 ;
        RECT 448.110 287.880 448.430 287.940 ;
        RECT 599.925 287.880 600.215 287.925 ;
        RECT 448.110 287.740 600.215 287.880 ;
        RECT 448.110 287.680 448.430 287.740 ;
        RECT 599.925 287.695 600.215 287.740 ;
        RECT 648.225 287.540 648.515 287.585 ;
        RECT 662.010 287.540 662.330 287.600 ;
        RECT 648.225 287.400 662.330 287.540 ;
        RECT 648.225 287.355 648.515 287.400 ;
        RECT 662.010 287.340 662.330 287.400 ;
        RECT 599.925 286.520 600.215 286.565 ;
        RECT 622.465 286.520 622.755 286.565 ;
        RECT 599.925 286.380 622.755 286.520 ;
        RECT 599.925 286.335 600.215 286.380 ;
        RECT 622.465 286.335 622.755 286.380 ;
        RECT 623.845 286.520 624.135 286.565 ;
        RECT 648.225 286.520 648.515 286.565 ;
        RECT 623.845 286.380 648.515 286.520 ;
        RECT 623.845 286.335 624.135 286.380 ;
        RECT 648.225 286.335 648.515 286.380 ;
        RECT 442.590 16.900 442.910 16.960 ;
        RECT 448.110 16.900 448.430 16.960 ;
        RECT 442.590 16.760 448.430 16.900 ;
        RECT 442.590 16.700 442.910 16.760 ;
        RECT 448.110 16.700 448.430 16.760 ;
      LAYER via ;
        RECT 448.140 287.680 448.400 287.940 ;
        RECT 662.040 287.340 662.300 287.600 ;
        RECT 442.620 16.700 442.880 16.960 ;
        RECT 448.140 16.700 448.400 16.960 ;
      LAYER met2 ;
        RECT 662.040 300.000 662.320 304.000 ;
        RECT 448.140 287.650 448.400 287.970 ;
        RECT 448.200 16.990 448.340 287.650 ;
        RECT 662.100 287.630 662.240 300.000 ;
        RECT 662.040 287.310 662.300 287.630 ;
        RECT 442.620 16.670 442.880 16.990 ;
        RECT 448.140 16.670 448.400 16.990 ;
        RECT 442.680 2.400 442.820 16.670 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 644.145 282.965 644.315 284.155 ;
      LAYER mcon ;
        RECT 644.145 283.985 644.315 284.155 ;
      LAYER met1 ;
        RECT 562.190 284.140 562.510 284.200 ;
        RECT 644.085 284.140 644.375 284.185 ;
        RECT 562.190 284.000 644.375 284.140 ;
        RECT 562.190 283.940 562.510 284.000 ;
        RECT 644.085 283.955 644.375 284.000 ;
        RECT 644.085 283.120 644.375 283.165 ;
        RECT 676.730 283.120 677.050 283.180 ;
        RECT 644.085 282.980 677.050 283.120 ;
        RECT 644.085 282.935 644.375 282.980 ;
        RECT 676.730 282.920 677.050 282.980 ;
        RECT 460.530 19.620 460.850 19.680 ;
        RECT 562.190 19.620 562.510 19.680 ;
        RECT 460.530 19.480 562.510 19.620 ;
        RECT 460.530 19.420 460.850 19.480 ;
        RECT 562.190 19.420 562.510 19.480 ;
      LAYER via ;
        RECT 562.220 283.940 562.480 284.200 ;
        RECT 676.760 282.920 677.020 283.180 ;
        RECT 460.560 19.420 460.820 19.680 ;
        RECT 562.220 19.420 562.480 19.680 ;
      LAYER met2 ;
        RECT 676.760 300.000 677.040 304.000 ;
        RECT 562.220 283.910 562.480 284.230 ;
        RECT 562.280 19.710 562.420 283.910 ;
        RECT 676.820 283.210 676.960 300.000 ;
        RECT 676.760 282.890 677.020 283.210 ;
        RECT 460.560 19.390 460.820 19.710 ;
        RECT 562.220 19.390 562.480 19.710 ;
        RECT 460.620 2.400 460.760 19.390 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 288.900 482.930 288.960 ;
        RECT 482.610 288.760 515.500 288.900 ;
        RECT 482.610 288.700 482.930 288.760 ;
        RECT 515.360 288.560 515.500 288.760 ;
        RECT 691.450 288.560 691.770 288.620 ;
        RECT 515.360 288.420 691.770 288.560 ;
        RECT 691.450 288.360 691.770 288.420 ;
        RECT 478.470 20.640 478.790 20.700 ;
        RECT 482.610 20.640 482.930 20.700 ;
        RECT 478.470 20.500 482.930 20.640 ;
        RECT 478.470 20.440 478.790 20.500 ;
        RECT 482.610 20.440 482.930 20.500 ;
      LAYER via ;
        RECT 482.640 288.700 482.900 288.960 ;
        RECT 691.480 288.360 691.740 288.620 ;
        RECT 478.500 20.440 478.760 20.700 ;
        RECT 482.640 20.440 482.900 20.700 ;
      LAYER met2 ;
        RECT 691.480 300.000 691.760 304.000 ;
        RECT 482.640 288.670 482.900 288.990 ;
        RECT 482.700 20.730 482.840 288.670 ;
        RECT 691.540 288.650 691.680 300.000 ;
        RECT 691.480 288.330 691.740 288.650 ;
        RECT 478.500 20.410 478.760 20.730 ;
        RECT 482.640 20.410 482.900 20.730 ;
        RECT 478.560 2.400 478.700 20.410 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 596.690 283.800 597.010 283.860 ;
        RECT 706.170 283.800 706.490 283.860 ;
        RECT 596.690 283.660 706.490 283.800 ;
        RECT 596.690 283.600 597.010 283.660 ;
        RECT 706.170 283.600 706.490 283.660 ;
        RECT 496.410 15.540 496.730 15.600 ;
        RECT 596.690 15.540 597.010 15.600 ;
        RECT 496.410 15.400 597.010 15.540 ;
        RECT 496.410 15.340 496.730 15.400 ;
        RECT 596.690 15.340 597.010 15.400 ;
      LAYER via ;
        RECT 596.720 283.600 596.980 283.860 ;
        RECT 706.200 283.600 706.460 283.860 ;
        RECT 496.440 15.340 496.700 15.600 ;
        RECT 596.720 15.340 596.980 15.600 ;
      LAYER met2 ;
        RECT 706.200 300.000 706.480 304.000 ;
        RECT 706.260 283.890 706.400 300.000 ;
        RECT 596.720 283.570 596.980 283.890 ;
        RECT 706.200 283.570 706.460 283.890 ;
        RECT 596.780 15.630 596.920 283.570 ;
        RECT 496.440 15.310 496.700 15.630 ;
        RECT 596.720 15.310 596.980 15.630 ;
        RECT 496.500 2.400 496.640 15.310 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 713.145 283.305 714.235 283.475 ;
      LAYER mcon ;
        RECT 714.065 283.305 714.235 283.475 ;
      LAYER met1 ;
        RECT 610.490 283.460 610.810 283.520 ;
        RECT 713.085 283.460 713.375 283.505 ;
        RECT 610.490 283.320 713.375 283.460 ;
        RECT 610.490 283.260 610.810 283.320 ;
        RECT 713.085 283.275 713.375 283.320 ;
        RECT 714.005 283.460 714.295 283.505 ;
        RECT 720.890 283.460 721.210 283.520 ;
        RECT 714.005 283.320 721.210 283.460 ;
        RECT 714.005 283.275 714.295 283.320 ;
        RECT 720.890 283.260 721.210 283.320 ;
        RECT 513.890 14.520 514.210 14.580 ;
        RECT 610.490 14.520 610.810 14.580 ;
        RECT 513.890 14.380 610.810 14.520 ;
        RECT 513.890 14.320 514.210 14.380 ;
        RECT 610.490 14.320 610.810 14.380 ;
      LAYER via ;
        RECT 610.520 283.260 610.780 283.520 ;
        RECT 720.920 283.260 721.180 283.520 ;
        RECT 513.920 14.320 514.180 14.580 ;
        RECT 610.520 14.320 610.780 14.580 ;
      LAYER met2 ;
        RECT 720.920 300.000 721.200 304.000 ;
        RECT 720.980 283.550 721.120 300.000 ;
        RECT 610.520 283.230 610.780 283.550 ;
        RECT 720.920 283.230 721.180 283.550 ;
        RECT 610.580 14.610 610.720 283.230 ;
        RECT 513.920 14.290 514.180 14.610 ;
        RECT 610.520 14.290 610.780 14.610 ;
        RECT 513.980 2.400 514.120 14.290 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 709.925 285.685 710.095 287.895 ;
      LAYER mcon ;
        RECT 709.925 287.725 710.095 287.895 ;
      LAYER met1 ;
        RECT 709.865 287.880 710.155 287.925 ;
        RECT 735.610 287.880 735.930 287.940 ;
        RECT 709.865 287.740 735.930 287.880 ;
        RECT 709.865 287.695 710.155 287.740 ;
        RECT 735.610 287.680 735.930 287.740 ;
        RECT 537.810 285.840 538.130 285.900 ;
        RECT 709.865 285.840 710.155 285.885 ;
        RECT 537.810 285.700 710.155 285.840 ;
        RECT 537.810 285.640 538.130 285.700 ;
        RECT 709.865 285.655 710.155 285.700 ;
        RECT 531.830 16.220 532.150 16.280 ;
        RECT 537.810 16.220 538.130 16.280 ;
        RECT 531.830 16.080 538.130 16.220 ;
        RECT 531.830 16.020 532.150 16.080 ;
        RECT 537.810 16.020 538.130 16.080 ;
      LAYER via ;
        RECT 735.640 287.680 735.900 287.940 ;
        RECT 537.840 285.640 538.100 285.900 ;
        RECT 531.860 16.020 532.120 16.280 ;
        RECT 537.840 16.020 538.100 16.280 ;
      LAYER met2 ;
        RECT 735.640 300.000 735.920 304.000 ;
        RECT 735.700 287.970 735.840 300.000 ;
        RECT 735.640 287.650 735.900 287.970 ;
        RECT 537.840 285.610 538.100 285.930 ;
        RECT 537.900 16.310 538.040 285.610 ;
        RECT 531.860 15.990 532.120 16.310 ;
        RECT 537.840 15.990 538.100 16.310 ;
        RECT 531.920 2.400 532.060 15.990 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 549.770 18.260 550.090 18.320 ;
        RECT 745.730 18.260 746.050 18.320 ;
        RECT 549.770 18.120 746.050 18.260 ;
        RECT 549.770 18.060 550.090 18.120 ;
        RECT 745.730 18.060 746.050 18.120 ;
      LAYER via ;
        RECT 549.800 18.060 550.060 18.320 ;
        RECT 745.760 18.060 746.020 18.320 ;
      LAYER met2 ;
        RECT 750.360 300.290 750.640 304.000 ;
        RECT 745.820 300.150 750.640 300.290 ;
        RECT 745.820 18.350 745.960 300.150 ;
        RECT 750.360 300.000 750.640 300.150 ;
        RECT 549.800 18.030 550.060 18.350 ;
        RECT 745.760 18.030 746.020 18.350 ;
        RECT 549.860 2.400 550.000 18.030 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 572.310 284.480 572.630 284.540 ;
        RECT 765.050 284.480 765.370 284.540 ;
        RECT 572.310 284.340 765.370 284.480 ;
        RECT 572.310 284.280 572.630 284.340 ;
        RECT 765.050 284.280 765.370 284.340 ;
        RECT 567.710 20.640 568.030 20.700 ;
        RECT 572.310 20.640 572.630 20.700 ;
        RECT 567.710 20.500 572.630 20.640 ;
        RECT 567.710 20.440 568.030 20.500 ;
        RECT 572.310 20.440 572.630 20.500 ;
      LAYER via ;
        RECT 572.340 284.280 572.600 284.540 ;
        RECT 765.080 284.280 765.340 284.540 ;
        RECT 567.740 20.440 568.000 20.700 ;
        RECT 572.340 20.440 572.600 20.700 ;
      LAYER met2 ;
        RECT 765.080 300.000 765.360 304.000 ;
        RECT 765.140 284.570 765.280 300.000 ;
        RECT 572.340 284.250 572.600 284.570 ;
        RECT 765.080 284.250 765.340 284.570 ;
        RECT 572.400 20.730 572.540 284.250 ;
        RECT 567.740 20.410 568.000 20.730 ;
        RECT 572.340 20.410 572.600 20.730 ;
        RECT 567.800 2.400 567.940 20.410 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 769.190 288.900 769.510 288.960 ;
        RECT 779.770 288.900 780.090 288.960 ;
        RECT 769.190 288.760 780.090 288.900 ;
        RECT 769.190 288.700 769.510 288.760 ;
        RECT 779.770 288.700 780.090 288.760 ;
        RECT 585.650 17.240 585.970 17.300 ;
        RECT 585.650 17.100 743.200 17.240 ;
        RECT 585.650 17.040 585.970 17.100 ;
        RECT 743.060 16.560 743.200 17.100 ;
        RECT 769.190 16.560 769.510 16.620 ;
        RECT 743.060 16.420 769.510 16.560 ;
        RECT 769.190 16.360 769.510 16.420 ;
      LAYER via ;
        RECT 769.220 288.700 769.480 288.960 ;
        RECT 779.800 288.700 780.060 288.960 ;
        RECT 585.680 17.040 585.940 17.300 ;
        RECT 769.220 16.360 769.480 16.620 ;
      LAYER met2 ;
        RECT 779.800 300.000 780.080 304.000 ;
        RECT 779.860 288.990 780.000 300.000 ;
        RECT 769.220 288.670 769.480 288.990 ;
        RECT 779.800 288.670 780.060 288.990 ;
        RECT 585.680 17.010 585.940 17.330 ;
        RECT 585.740 2.400 585.880 17.010 ;
        RECT 769.280 16.650 769.420 288.670 ;
        RECT 769.220 16.330 769.480 16.650 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 179.545 18.445 179.715 20.315 ;
        RECT 227.385 18.445 227.555 20.315 ;
        RECT 276.145 18.445 276.315 21.335 ;
        RECT 323.985 18.445 324.155 21.335 ;
        RECT 324.445 17.255 324.615 18.615 ;
        RECT 359.405 17.255 359.575 17.935 ;
        RECT 324.445 17.085 325.995 17.255 ;
        RECT 358.945 17.085 359.575 17.255 ;
      LAYER mcon ;
        RECT 276.145 21.165 276.315 21.335 ;
        RECT 179.545 20.145 179.715 20.315 ;
        RECT 227.385 20.145 227.555 20.315 ;
        RECT 323.985 21.165 324.155 21.335 ;
        RECT 324.445 18.445 324.615 18.615 ;
        RECT 359.405 17.765 359.575 17.935 ;
        RECT 325.825 17.085 325.995 17.255 ;
      LAYER met1 ;
        RECT 368.990 286.180 369.310 286.240 ;
        RECT 373.130 286.180 373.450 286.240 ;
        RECT 368.990 286.040 373.450 286.180 ;
        RECT 368.990 285.980 369.310 286.040 ;
        RECT 373.130 285.980 373.450 286.040 ;
        RECT 276.085 21.320 276.375 21.365 ;
        RECT 323.925 21.320 324.215 21.365 ;
        RECT 276.085 21.180 324.215 21.320 ;
        RECT 276.085 21.135 276.375 21.180 ;
        RECT 323.925 21.135 324.215 21.180 ;
        RECT 179.485 20.300 179.775 20.345 ;
        RECT 227.325 20.300 227.615 20.345 ;
        RECT 179.485 20.160 227.615 20.300 ;
        RECT 179.485 20.115 179.775 20.160 ;
        RECT 227.325 20.115 227.615 20.160 ;
        RECT 91.610 18.600 91.930 18.660 ;
        RECT 179.485 18.600 179.775 18.645 ;
        RECT 91.610 18.460 179.775 18.600 ;
        RECT 91.610 18.400 91.930 18.460 ;
        RECT 179.485 18.415 179.775 18.460 ;
        RECT 227.325 18.600 227.615 18.645 ;
        RECT 276.085 18.600 276.375 18.645 ;
        RECT 227.325 18.460 276.375 18.600 ;
        RECT 227.325 18.415 227.615 18.460 ;
        RECT 276.085 18.415 276.375 18.460 ;
        RECT 323.925 18.600 324.215 18.645 ;
        RECT 324.385 18.600 324.675 18.645 ;
        RECT 323.925 18.460 324.675 18.600 ;
        RECT 323.925 18.415 324.215 18.460 ;
        RECT 324.385 18.415 324.675 18.460 ;
        RECT 359.345 17.920 359.635 17.965 ;
        RECT 368.990 17.920 369.310 17.980 ;
        RECT 359.345 17.780 369.310 17.920 ;
        RECT 359.345 17.735 359.635 17.780 ;
        RECT 368.990 17.720 369.310 17.780 ;
        RECT 325.765 17.240 326.055 17.285 ;
        RECT 358.885 17.240 359.175 17.285 ;
        RECT 325.765 17.100 359.175 17.240 ;
        RECT 325.765 17.055 326.055 17.100 ;
        RECT 358.885 17.055 359.175 17.100 ;
      LAYER via ;
        RECT 369.020 285.980 369.280 286.240 ;
        RECT 373.160 285.980 373.420 286.240 ;
        RECT 91.640 18.400 91.900 18.660 ;
        RECT 369.020 17.720 369.280 17.980 ;
      LAYER met2 ;
        RECT 373.160 300.000 373.440 304.000 ;
        RECT 373.220 286.270 373.360 300.000 ;
        RECT 369.020 285.950 369.280 286.270 ;
        RECT 373.160 285.950 373.420 286.270 ;
        RECT 91.640 18.370 91.900 18.690 ;
        RECT 91.700 2.400 91.840 18.370 ;
        RECT 369.080 18.010 369.220 285.950 ;
        RECT 369.020 17.690 369.280 18.010 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 284.820 607.130 284.880 ;
        RECT 794.490 284.820 794.810 284.880 ;
        RECT 606.810 284.680 794.810 284.820 ;
        RECT 606.810 284.620 607.130 284.680 ;
        RECT 794.490 284.620 794.810 284.680 ;
        RECT 603.130 20.640 603.450 20.700 ;
        RECT 606.810 20.640 607.130 20.700 ;
        RECT 603.130 20.500 607.130 20.640 ;
        RECT 603.130 20.440 603.450 20.500 ;
        RECT 606.810 20.440 607.130 20.500 ;
      LAYER via ;
        RECT 606.840 284.620 607.100 284.880 ;
        RECT 794.520 284.620 794.780 284.880 ;
        RECT 603.160 20.440 603.420 20.700 ;
        RECT 606.840 20.440 607.100 20.700 ;
      LAYER met2 ;
        RECT 794.520 300.000 794.800 304.000 ;
        RECT 794.580 284.910 794.720 300.000 ;
        RECT 606.840 284.590 607.100 284.910 ;
        RECT 794.520 284.590 794.780 284.910 ;
        RECT 606.900 20.730 607.040 284.590 ;
        RECT 603.160 20.410 603.420 20.730 ;
        RECT 606.840 20.410 607.100 20.730 ;
        RECT 603.220 2.400 603.360 20.410 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 809.210 286.520 809.530 286.580 ;
        RECT 648.760 286.380 809.530 286.520 ;
        RECT 627.510 286.180 627.830 286.240 ;
        RECT 648.760 286.180 648.900 286.380 ;
        RECT 809.210 286.320 809.530 286.380 ;
        RECT 627.510 286.040 648.900 286.180 ;
        RECT 627.510 285.980 627.830 286.040 ;
        RECT 621.070 18.600 621.390 18.660 ;
        RECT 627.510 18.600 627.830 18.660 ;
        RECT 621.070 18.460 627.830 18.600 ;
        RECT 621.070 18.400 621.390 18.460 ;
        RECT 627.510 18.400 627.830 18.460 ;
      LAYER via ;
        RECT 627.540 285.980 627.800 286.240 ;
        RECT 809.240 286.320 809.500 286.580 ;
        RECT 621.100 18.400 621.360 18.660 ;
        RECT 627.540 18.400 627.800 18.660 ;
      LAYER met2 ;
        RECT 809.240 300.000 809.520 304.000 ;
        RECT 809.300 286.610 809.440 300.000 ;
        RECT 809.240 286.290 809.500 286.610 ;
        RECT 627.540 285.950 627.800 286.270 ;
        RECT 627.600 18.690 627.740 285.950 ;
        RECT 621.100 18.370 621.360 18.690 ;
        RECT 627.540 18.370 627.800 18.690 ;
        RECT 621.160 2.400 621.300 18.370 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 116.910 287.540 117.230 287.600 ;
        RECT 392.910 287.540 393.230 287.600 ;
        RECT 116.910 287.400 393.230 287.540 ;
        RECT 116.910 287.340 117.230 287.400 ;
        RECT 392.910 287.340 393.230 287.400 ;
      LAYER via ;
        RECT 116.940 287.340 117.200 287.600 ;
        RECT 392.940 287.340 393.200 287.600 ;
      LAYER met2 ;
        RECT 392.940 300.000 393.220 304.000 ;
        RECT 393.000 287.630 393.140 300.000 ;
        RECT 116.940 287.310 117.200 287.630 ;
        RECT 392.940 287.310 393.200 287.630 ;
        RECT 117.000 17.410 117.140 287.310 ;
        RECT 115.620 17.270 117.140 17.410 ;
        RECT 115.620 2.400 115.760 17.270 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 348.365 15.385 348.535 18.615 ;
      LAYER mcon ;
        RECT 348.365 18.445 348.535 18.615 ;
      LAYER met1 ;
        RECT 375.890 286.180 376.210 286.240 ;
        RECT 412.230 286.180 412.550 286.240 ;
        RECT 375.890 286.040 412.550 286.180 ;
        RECT 375.890 285.980 376.210 286.040 ;
        RECT 412.230 285.980 412.550 286.040 ;
        RECT 348.305 18.600 348.595 18.645 ;
        RECT 375.890 18.600 376.210 18.660 ;
        RECT 348.305 18.460 376.210 18.600 ;
        RECT 348.305 18.415 348.595 18.460 ;
        RECT 375.890 18.400 376.210 18.460 ;
        RECT 139.450 15.540 139.770 15.600 ;
        RECT 348.305 15.540 348.595 15.585 ;
        RECT 139.450 15.400 348.595 15.540 ;
        RECT 139.450 15.340 139.770 15.400 ;
        RECT 348.305 15.355 348.595 15.400 ;
      LAYER via ;
        RECT 375.920 285.980 376.180 286.240 ;
        RECT 412.260 285.980 412.520 286.240 ;
        RECT 375.920 18.400 376.180 18.660 ;
        RECT 139.480 15.340 139.740 15.600 ;
      LAYER met2 ;
        RECT 412.260 300.000 412.540 304.000 ;
        RECT 412.320 286.270 412.460 300.000 ;
        RECT 375.920 285.950 376.180 286.270 ;
        RECT 412.260 285.950 412.520 286.270 ;
        RECT 375.980 18.690 376.120 285.950 ;
        RECT 375.920 18.370 376.180 18.690 ;
        RECT 139.480 15.310 139.740 15.630 ;
        RECT 139.540 2.400 139.680 15.310 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 287.880 158.630 287.940 ;
        RECT 426.950 287.880 427.270 287.940 ;
        RECT 158.310 287.740 427.270 287.880 ;
        RECT 158.310 287.680 158.630 287.740 ;
        RECT 426.950 287.680 427.270 287.740 ;
      LAYER via ;
        RECT 158.340 287.680 158.600 287.940 ;
        RECT 426.980 287.680 427.240 287.940 ;
      LAYER met2 ;
        RECT 426.980 300.000 427.260 304.000 ;
        RECT 427.040 287.970 427.180 300.000 ;
        RECT 158.340 287.650 158.600 287.970 ;
        RECT 426.980 287.650 427.240 287.970 ;
        RECT 158.400 17.410 158.540 287.650 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 174.870 19.280 175.190 19.340 ;
        RECT 441.670 19.280 441.990 19.340 ;
        RECT 174.870 19.140 441.990 19.280 ;
        RECT 174.870 19.080 175.190 19.140 ;
        RECT 441.670 19.080 441.990 19.140 ;
      LAYER via ;
        RECT 174.900 19.080 175.160 19.340 ;
        RECT 441.700 19.080 441.960 19.340 ;
      LAYER met2 ;
        RECT 441.700 300.000 441.980 304.000 ;
        RECT 441.760 19.370 441.900 300.000 ;
        RECT 174.900 19.050 175.160 19.370 ;
        RECT 441.700 19.050 441.960 19.370 ;
        RECT 174.960 2.400 175.100 19.050 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.810 288.560 193.130 288.620 ;
        RECT 456.390 288.560 456.710 288.620 ;
        RECT 192.810 288.420 456.710 288.560 ;
        RECT 192.810 288.360 193.130 288.420 ;
        RECT 456.390 288.360 456.710 288.420 ;
      LAYER via ;
        RECT 192.840 288.360 193.100 288.620 ;
        RECT 456.420 288.360 456.680 288.620 ;
      LAYER met2 ;
        RECT 456.420 300.000 456.700 304.000 ;
        RECT 456.480 288.650 456.620 300.000 ;
        RECT 192.840 288.330 193.100 288.650 ;
        RECT 456.420 288.330 456.680 288.650 ;
        RECT 192.900 2.400 193.040 288.330 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 228.305 16.405 228.475 20.315 ;
        RECT 444.965 19.125 445.135 20.315 ;
      LAYER mcon ;
        RECT 228.305 20.145 228.475 20.315 ;
        RECT 444.965 20.145 445.135 20.315 ;
      LAYER met1 ;
        RECT 228.245 20.300 228.535 20.345 ;
        RECT 444.905 20.300 445.195 20.345 ;
        RECT 228.245 20.160 445.195 20.300 ;
        RECT 228.245 20.115 228.535 20.160 ;
        RECT 444.905 20.115 445.195 20.160 ;
        RECT 444.905 19.280 445.195 19.325 ;
        RECT 469.270 19.280 469.590 19.340 ;
        RECT 444.905 19.140 469.590 19.280 ;
        RECT 444.905 19.095 445.195 19.140 ;
        RECT 469.270 19.080 469.590 19.140 ;
        RECT 228.245 16.560 228.535 16.605 ;
        RECT 220.960 16.420 228.535 16.560 ;
        RECT 210.750 16.220 211.070 16.280 ;
        RECT 220.960 16.220 221.100 16.420 ;
        RECT 228.245 16.375 228.535 16.420 ;
        RECT 210.750 16.080 221.100 16.220 ;
        RECT 210.750 16.020 211.070 16.080 ;
      LAYER via ;
        RECT 469.300 19.080 469.560 19.340 ;
        RECT 210.780 16.020 211.040 16.280 ;
      LAYER met2 ;
        RECT 471.140 300.290 471.420 304.000 ;
        RECT 469.360 300.150 471.420 300.290 ;
        RECT 469.360 19.370 469.500 300.150 ;
        RECT 471.140 300.000 471.420 300.150 ;
        RECT 469.300 19.050 469.560 19.370 ;
        RECT 210.780 15.990 211.040 16.310 ;
        RECT 210.840 2.400 210.980 15.990 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 458.305 284.665 458.475 285.855 ;
      LAYER mcon ;
        RECT 458.305 285.685 458.475 285.855 ;
      LAYER met1 ;
        RECT 458.245 285.840 458.535 285.885 ;
        RECT 485.830 285.840 486.150 285.900 ;
        RECT 458.245 285.700 486.150 285.840 ;
        RECT 458.245 285.655 458.535 285.700 ;
        RECT 485.830 285.640 486.150 285.700 ;
        RECT 234.210 284.820 234.530 284.880 ;
        RECT 458.245 284.820 458.535 284.865 ;
        RECT 234.210 284.680 458.535 284.820 ;
        RECT 234.210 284.620 234.530 284.680 ;
        RECT 458.245 284.635 458.535 284.680 ;
        RECT 228.690 16.560 229.010 16.620 ;
        RECT 234.210 16.560 234.530 16.620 ;
        RECT 228.690 16.420 234.530 16.560 ;
        RECT 228.690 16.360 229.010 16.420 ;
        RECT 234.210 16.360 234.530 16.420 ;
      LAYER via ;
        RECT 485.860 285.640 486.120 285.900 ;
        RECT 234.240 284.620 234.500 284.880 ;
        RECT 228.720 16.360 228.980 16.620 ;
        RECT 234.240 16.360 234.500 16.620 ;
      LAYER met2 ;
        RECT 485.860 300.000 486.140 304.000 ;
        RECT 485.920 285.930 486.060 300.000 ;
        RECT 485.860 285.610 486.120 285.930 ;
        RECT 234.240 284.590 234.500 284.910 ;
        RECT 234.300 16.650 234.440 284.590 ;
        RECT 228.720 16.330 228.980 16.650 ;
        RECT 234.240 16.330 234.500 16.650 ;
        RECT 228.780 2.400 228.920 16.330 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 50.210 18.600 50.530 18.660 ;
        RECT 50.210 18.460 82.640 18.600 ;
        RECT 50.210 18.400 50.530 18.460 ;
        RECT 82.500 17.920 82.640 18.460 ;
        RECT 339.090 17.920 339.410 17.980 ;
        RECT 82.500 17.780 339.410 17.920 ;
        RECT 339.090 17.720 339.410 17.780 ;
      LAYER via ;
        RECT 50.240 18.400 50.500 18.660 ;
        RECT 339.120 17.720 339.380 17.980 ;
      LAYER met2 ;
        RECT 339.120 300.000 339.400 304.000 ;
        RECT 50.240 18.370 50.500 18.690 ;
        RECT 50.300 2.400 50.440 18.370 ;
        RECT 339.180 18.010 339.320 300.000 ;
        RECT 339.120 17.690 339.380 18.010 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 285.160 255.230 285.220 ;
        RECT 505.610 285.160 505.930 285.220 ;
        RECT 254.910 285.020 505.930 285.160 ;
        RECT 254.910 284.960 255.230 285.020 ;
        RECT 505.610 284.960 505.930 285.020 ;
        RECT 252.610 16.560 252.930 16.620 ;
        RECT 254.910 16.560 255.230 16.620 ;
        RECT 252.610 16.420 255.230 16.560 ;
        RECT 252.610 16.360 252.930 16.420 ;
        RECT 254.910 16.360 255.230 16.420 ;
      LAYER via ;
        RECT 254.940 284.960 255.200 285.220 ;
        RECT 505.640 284.960 505.900 285.220 ;
        RECT 252.640 16.360 252.900 16.620 ;
        RECT 254.940 16.360 255.200 16.620 ;
      LAYER met2 ;
        RECT 505.640 300.000 505.920 304.000 ;
        RECT 505.700 285.250 505.840 300.000 ;
        RECT 254.940 284.930 255.200 285.250 ;
        RECT 505.640 284.930 505.900 285.250 ;
        RECT 255.000 16.650 255.140 284.930 ;
        RECT 252.640 16.330 252.900 16.650 ;
        RECT 254.940 16.330 255.200 16.650 ;
        RECT 252.700 2.400 252.840 16.330 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 513.890 283.460 514.210 283.520 ;
        RECT 520.330 283.460 520.650 283.520 ;
        RECT 513.890 283.320 520.650 283.460 ;
        RECT 513.890 283.260 514.210 283.320 ;
        RECT 520.330 283.260 520.650 283.320 ;
        RECT 270.090 16.220 270.410 16.280 ;
        RECT 513.890 16.220 514.210 16.280 ;
        RECT 270.090 16.080 514.210 16.220 ;
        RECT 270.090 16.020 270.410 16.080 ;
        RECT 513.890 16.020 514.210 16.080 ;
      LAYER via ;
        RECT 513.920 283.260 514.180 283.520 ;
        RECT 520.360 283.260 520.620 283.520 ;
        RECT 270.120 16.020 270.380 16.280 ;
        RECT 513.920 16.020 514.180 16.280 ;
      LAYER met2 ;
        RECT 520.360 300.000 520.640 304.000 ;
        RECT 520.420 283.550 520.560 300.000 ;
        RECT 513.920 283.230 514.180 283.550 ;
        RECT 520.360 283.230 520.620 283.550 ;
        RECT 513.980 16.310 514.120 283.230 ;
        RECT 270.120 15.990 270.380 16.310 ;
        RECT 513.920 15.990 514.180 16.310 ;
        RECT 270.180 2.400 270.320 15.990 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 314.785 283.645 314.955 284.495 ;
      LAYER mcon ;
        RECT 314.785 284.325 314.955 284.495 ;
      LAYER met1 ;
        RECT 314.725 284.480 315.015 284.525 ;
        RECT 535.050 284.480 535.370 284.540 ;
        RECT 314.725 284.340 535.370 284.480 ;
        RECT 314.725 284.295 315.015 284.340 ;
        RECT 535.050 284.280 535.370 284.340 ;
        RECT 289.410 283.800 289.730 283.860 ;
        RECT 314.725 283.800 315.015 283.845 ;
        RECT 289.410 283.660 315.015 283.800 ;
        RECT 289.410 283.600 289.730 283.660 ;
        RECT 314.725 283.615 315.015 283.660 ;
      LAYER via ;
        RECT 535.080 284.280 535.340 284.540 ;
        RECT 289.440 283.600 289.700 283.860 ;
      LAYER met2 ;
        RECT 535.080 300.000 535.360 304.000 ;
        RECT 535.140 284.570 535.280 300.000 ;
        RECT 535.080 284.250 535.340 284.570 ;
        RECT 289.440 283.570 289.700 283.890 ;
        RECT 289.500 3.130 289.640 283.570 ;
        RECT 288.120 2.990 289.640 3.130 ;
        RECT 288.120 2.400 288.260 2.990 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 341.005 18.105 342.095 18.275 ;
        RECT 341.005 17.425 341.175 18.105 ;
      LAYER mcon ;
        RECT 341.925 18.105 342.095 18.275 ;
      LAYER met1 ;
        RECT 541.490 283.800 541.810 283.860 ;
        RECT 549.310 283.800 549.630 283.860 ;
        RECT 541.490 283.660 549.630 283.800 ;
        RECT 541.490 283.600 541.810 283.660 ;
        RECT 549.310 283.600 549.630 283.660 ;
        RECT 341.865 18.260 342.155 18.305 ;
        RECT 541.490 18.260 541.810 18.320 ;
        RECT 341.865 18.120 541.810 18.260 ;
        RECT 341.865 18.075 342.155 18.120 ;
        RECT 541.490 18.060 541.810 18.120 ;
        RECT 305.970 17.580 306.290 17.640 ;
        RECT 340.945 17.580 341.235 17.625 ;
        RECT 305.970 17.440 341.235 17.580 ;
        RECT 305.970 17.380 306.290 17.440 ;
        RECT 340.945 17.395 341.235 17.440 ;
      LAYER via ;
        RECT 541.520 283.600 541.780 283.860 ;
        RECT 549.340 283.600 549.600 283.860 ;
        RECT 541.520 18.060 541.780 18.320 ;
        RECT 306.000 17.380 306.260 17.640 ;
      LAYER met2 ;
        RECT 549.340 300.000 549.620 304.000 ;
        RECT 549.400 283.890 549.540 300.000 ;
        RECT 541.520 283.570 541.780 283.890 ;
        RECT 549.340 283.570 549.600 283.890 ;
        RECT 541.580 18.350 541.720 283.570 ;
        RECT 541.520 18.030 541.780 18.350 ;
        RECT 306.000 17.350 306.260 17.670 ;
        RECT 306.060 2.400 306.200 17.350 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 510.285 283.645 510.455 285.515 ;
      LAYER mcon ;
        RECT 510.285 285.345 510.455 285.515 ;
      LAYER met1 ;
        RECT 510.225 285.500 510.515 285.545 ;
        RECT 564.030 285.500 564.350 285.560 ;
        RECT 510.225 285.360 564.350 285.500 ;
        RECT 510.225 285.315 510.515 285.360 ;
        RECT 564.030 285.300 564.350 285.360 ;
        RECT 323.910 283.800 324.230 283.860 ;
        RECT 510.225 283.800 510.515 283.845 ;
        RECT 323.910 283.660 510.515 283.800 ;
        RECT 323.910 283.600 324.230 283.660 ;
        RECT 510.225 283.615 510.515 283.660 ;
      LAYER via ;
        RECT 564.060 285.300 564.320 285.560 ;
        RECT 323.940 283.600 324.200 283.860 ;
      LAYER met2 ;
        RECT 564.060 300.000 564.340 304.000 ;
        RECT 564.120 285.590 564.260 300.000 ;
        RECT 564.060 285.270 564.320 285.590 ;
        RECT 323.940 283.570 324.200 283.890 ;
        RECT 324.000 2.400 324.140 283.570 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 520.865 16.745 521.035 17.595 ;
      LAYER mcon ;
        RECT 520.865 17.425 521.035 17.595 ;
      LAYER met1 ;
        RECT 548.390 283.120 548.710 283.180 ;
        RECT 578.750 283.120 579.070 283.180 ;
        RECT 548.390 282.980 579.070 283.120 ;
        RECT 548.390 282.920 548.710 282.980 ;
        RECT 578.750 282.920 579.070 282.980 ;
        RECT 341.390 17.580 341.710 17.640 ;
        RECT 520.805 17.580 521.095 17.625 ;
        RECT 341.390 17.440 521.095 17.580 ;
        RECT 341.390 17.380 341.710 17.440 ;
        RECT 520.805 17.395 521.095 17.440 ;
        RECT 520.805 16.900 521.095 16.945 ;
        RECT 548.390 16.900 548.710 16.960 ;
        RECT 520.805 16.760 548.710 16.900 ;
        RECT 520.805 16.715 521.095 16.760 ;
        RECT 548.390 16.700 548.710 16.760 ;
      LAYER via ;
        RECT 548.420 282.920 548.680 283.180 ;
        RECT 578.780 282.920 579.040 283.180 ;
        RECT 341.420 17.380 341.680 17.640 ;
        RECT 548.420 16.700 548.680 16.960 ;
      LAYER met2 ;
        RECT 578.780 300.000 579.060 304.000 ;
        RECT 578.840 283.210 578.980 300.000 ;
        RECT 548.420 282.890 548.680 283.210 ;
        RECT 578.780 282.890 579.040 283.210 ;
        RECT 341.420 17.350 341.680 17.670 ;
        RECT 341.480 2.400 341.620 17.350 ;
        RECT 548.480 16.990 548.620 282.890 ;
        RECT 548.420 16.670 548.680 16.990 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 575.990 286.180 576.310 286.240 ;
        RECT 593.470 286.180 593.790 286.240 ;
        RECT 575.990 286.040 593.790 286.180 ;
        RECT 575.990 285.980 576.310 286.040 ;
        RECT 593.470 285.980 593.790 286.040 ;
        RECT 359.330 17.240 359.650 17.300 ;
        RECT 575.990 17.240 576.310 17.300 ;
        RECT 359.330 17.100 576.310 17.240 ;
        RECT 359.330 17.040 359.650 17.100 ;
        RECT 575.990 17.040 576.310 17.100 ;
      LAYER via ;
        RECT 576.020 285.980 576.280 286.240 ;
        RECT 593.500 285.980 593.760 286.240 ;
        RECT 359.360 17.040 359.620 17.300 ;
        RECT 576.020 17.040 576.280 17.300 ;
      LAYER met2 ;
        RECT 593.500 300.000 593.780 304.000 ;
        RECT 593.560 286.270 593.700 300.000 ;
        RECT 576.020 285.950 576.280 286.270 ;
        RECT 593.500 285.950 593.760 286.270 ;
        RECT 576.080 17.330 576.220 285.950 ;
        RECT 359.360 17.010 359.620 17.330 ;
        RECT 576.020 17.010 576.280 17.330 ;
        RECT 359.420 2.400 359.560 17.010 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 412.765 286.025 412.935 286.875 ;
        RECT 575.605 284.665 575.775 286.195 ;
      LAYER mcon ;
        RECT 412.765 286.705 412.935 286.875 ;
        RECT 575.605 286.025 575.775 286.195 ;
      LAYER met1 ;
        RECT 412.705 286.860 412.995 286.905 ;
        RECT 398.060 286.720 412.995 286.860 ;
        RECT 379.110 286.520 379.430 286.580 ;
        RECT 398.060 286.520 398.200 286.720 ;
        RECT 412.705 286.675 412.995 286.720 ;
        RECT 379.110 286.380 398.200 286.520 ;
        RECT 379.110 286.320 379.430 286.380 ;
        RECT 412.705 286.180 412.995 286.225 ;
        RECT 575.545 286.180 575.835 286.225 ;
        RECT 412.705 286.040 575.835 286.180 ;
        RECT 412.705 285.995 412.995 286.040 ;
        RECT 575.545 285.995 575.835 286.040 ;
        RECT 575.545 284.820 575.835 284.865 ;
        RECT 606.350 284.820 606.670 284.880 ;
        RECT 575.545 284.680 606.670 284.820 ;
        RECT 575.545 284.635 575.835 284.680 ;
        RECT 606.350 284.620 606.670 284.680 ;
      LAYER via ;
        RECT 379.140 286.320 379.400 286.580 ;
        RECT 606.380 284.620 606.640 284.880 ;
      LAYER met2 ;
        RECT 608.220 300.290 608.500 304.000 ;
        RECT 607.360 300.150 608.500 300.290 ;
        RECT 379.140 286.290 379.400 286.610 ;
        RECT 379.200 3.130 379.340 286.290 ;
        RECT 607.360 285.330 607.500 300.150 ;
        RECT 608.220 300.000 608.500 300.150 ;
        RECT 606.440 285.190 607.500 285.330 ;
        RECT 606.440 284.910 606.580 285.190 ;
        RECT 606.380 284.590 606.640 284.910 ;
        RECT 377.360 2.990 379.340 3.130 ;
        RECT 377.360 2.400 377.500 2.990 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 622.910 286.860 623.230 286.920 ;
        RECT 599.540 286.720 623.230 286.860 ;
        RECT 399.810 286.520 400.130 286.580 ;
        RECT 599.540 286.520 599.680 286.720 ;
        RECT 622.910 286.660 623.230 286.720 ;
        RECT 399.810 286.380 599.680 286.520 ;
        RECT 399.810 286.320 400.130 286.380 ;
        RECT 395.210 17.920 395.530 17.980 ;
        RECT 399.810 17.920 400.130 17.980 ;
        RECT 395.210 17.780 400.130 17.920 ;
        RECT 395.210 17.720 395.530 17.780 ;
        RECT 399.810 17.720 400.130 17.780 ;
      LAYER via ;
        RECT 399.840 286.320 400.100 286.580 ;
        RECT 622.940 286.660 623.200 286.920 ;
        RECT 395.240 17.720 395.500 17.980 ;
        RECT 399.840 17.720 400.100 17.980 ;
      LAYER met2 ;
        RECT 622.940 300.000 623.220 304.000 ;
        RECT 623.000 286.950 623.140 300.000 ;
        RECT 622.940 286.630 623.200 286.950 ;
        RECT 399.840 286.290 400.100 286.610 ;
        RECT 399.900 18.010 400.040 286.290 ;
        RECT 395.240 17.690 395.500 18.010 ;
        RECT 399.840 17.690 400.100 18.010 ;
        RECT 395.300 2.400 395.440 17.690 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 413.150 18.600 413.470 18.660 ;
        RECT 576.450 18.600 576.770 18.660 ;
        RECT 413.150 18.460 576.770 18.600 ;
        RECT 413.150 18.400 413.470 18.460 ;
        RECT 576.450 18.400 576.770 18.460 ;
      LAYER via ;
        RECT 413.180 18.400 413.440 18.660 ;
        RECT 576.480 18.400 576.740 18.660 ;
      LAYER met2 ;
        RECT 637.660 300.000 637.940 304.000 ;
        RECT 637.720 286.125 637.860 300.000 ;
        RECT 576.470 285.755 576.750 286.125 ;
        RECT 637.650 285.755 637.930 286.125 ;
        RECT 576.540 18.690 576.680 285.755 ;
        RECT 413.180 18.370 413.440 18.690 ;
        RECT 576.480 18.370 576.740 18.690 ;
        RECT 413.240 2.400 413.380 18.370 ;
        RECT 413.030 -4.800 413.590 2.400 ;
      LAYER via2 ;
        RECT 576.470 285.800 576.750 286.080 ;
        RECT 637.650 285.800 637.930 286.080 ;
      LAYER met3 ;
        RECT 576.445 286.090 576.775 286.105 ;
        RECT 637.625 286.090 637.955 286.105 ;
        RECT 576.445 285.790 637.955 286.090 ;
        RECT 576.445 285.775 576.775 285.790 ;
        RECT 637.625 285.775 637.955 285.790 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 324.445 286.705 325.075 286.875 ;
        RECT 324.905 286.025 325.075 286.705 ;
      LAYER met1 ;
        RECT 75.510 286.860 75.830 286.920 ;
        RECT 324.385 286.860 324.675 286.905 ;
        RECT 75.510 286.720 324.675 286.860 ;
        RECT 75.510 286.660 75.830 286.720 ;
        RECT 324.385 286.675 324.675 286.720 ;
        RECT 324.845 286.180 325.135 286.225 ;
        RECT 358.410 286.180 358.730 286.240 ;
        RECT 324.845 286.040 358.730 286.180 ;
        RECT 324.845 285.995 325.135 286.040 ;
        RECT 358.410 285.980 358.730 286.040 ;
        RECT 74.130 2.960 74.450 3.020 ;
        RECT 75.510 2.960 75.830 3.020 ;
        RECT 74.130 2.820 75.830 2.960 ;
        RECT 74.130 2.760 74.450 2.820 ;
        RECT 75.510 2.760 75.830 2.820 ;
      LAYER via ;
        RECT 75.540 286.660 75.800 286.920 ;
        RECT 358.440 285.980 358.700 286.240 ;
        RECT 74.160 2.760 74.420 3.020 ;
        RECT 75.540 2.760 75.800 3.020 ;
      LAYER met2 ;
        RECT 358.440 300.000 358.720 304.000 ;
        RECT 75.540 286.630 75.800 286.950 ;
        RECT 75.600 3.050 75.740 286.630 ;
        RECT 358.500 286.270 358.640 300.000 ;
        RECT 358.440 285.950 358.700 286.270 ;
        RECT 74.160 2.730 74.420 3.050 ;
        RECT 75.540 2.730 75.800 3.050 ;
        RECT 74.220 2.400 74.360 2.730 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 612.865 287.045 613.035 287.895 ;
      LAYER mcon ;
        RECT 612.865 287.725 613.035 287.895 ;
      LAYER met1 ;
        RECT 612.805 287.880 613.095 287.925 ;
        RECT 652.350 287.880 652.670 287.940 ;
        RECT 612.805 287.740 652.670 287.880 ;
        RECT 612.805 287.695 613.095 287.740 ;
        RECT 652.350 287.680 652.670 287.740 ;
        RECT 434.310 287.540 434.630 287.600 ;
        RECT 434.310 287.400 472.720 287.540 ;
        RECT 434.310 287.340 434.630 287.400 ;
        RECT 472.580 287.200 472.720 287.400 ;
        RECT 612.805 287.200 613.095 287.245 ;
        RECT 472.580 287.060 613.095 287.200 ;
        RECT 612.805 287.015 613.095 287.060 ;
        RECT 430.630 16.900 430.950 16.960 ;
        RECT 434.310 16.900 434.630 16.960 ;
        RECT 430.630 16.760 434.630 16.900 ;
        RECT 430.630 16.700 430.950 16.760 ;
        RECT 434.310 16.700 434.630 16.760 ;
      LAYER via ;
        RECT 652.380 287.680 652.640 287.940 ;
        RECT 434.340 287.340 434.600 287.600 ;
        RECT 430.660 16.700 430.920 16.960 ;
        RECT 434.340 16.700 434.600 16.960 ;
      LAYER met2 ;
        RECT 652.380 300.000 652.660 304.000 ;
        RECT 652.440 287.970 652.580 300.000 ;
        RECT 652.380 287.650 652.640 287.970 ;
        RECT 434.340 287.310 434.600 287.630 ;
        RECT 434.400 16.990 434.540 287.310 ;
        RECT 430.660 16.670 430.920 16.990 ;
        RECT 434.340 16.670 434.600 16.990 ;
        RECT 430.720 2.400 430.860 16.670 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 652.885 282.625 653.055 287.895 ;
      LAYER mcon ;
        RECT 652.885 287.725 653.055 287.895 ;
      LAYER met1 ;
        RECT 652.825 287.880 653.115 287.925 ;
        RECT 667.070 287.880 667.390 287.940 ;
        RECT 652.825 287.740 667.390 287.880 ;
        RECT 652.825 287.695 653.115 287.740 ;
        RECT 667.070 287.680 667.390 287.740 ;
        RECT 610.950 283.120 611.270 283.180 ;
        RECT 610.950 282.980 643.840 283.120 ;
        RECT 610.950 282.920 611.270 282.980 ;
        RECT 643.700 282.780 643.840 282.980 ;
        RECT 652.825 282.780 653.115 282.825 ;
        RECT 643.700 282.640 653.115 282.780 ;
        RECT 652.825 282.595 653.115 282.640 ;
        RECT 448.570 18.940 448.890 19.000 ;
        RECT 610.950 18.940 611.270 19.000 ;
        RECT 448.570 18.800 611.270 18.940 ;
        RECT 448.570 18.740 448.890 18.800 ;
        RECT 610.950 18.740 611.270 18.800 ;
      LAYER via ;
        RECT 667.100 287.680 667.360 287.940 ;
        RECT 610.980 282.920 611.240 283.180 ;
        RECT 448.600 18.740 448.860 19.000 ;
        RECT 610.980 18.740 611.240 19.000 ;
      LAYER met2 ;
        RECT 667.100 300.000 667.380 304.000 ;
        RECT 667.160 287.970 667.300 300.000 ;
        RECT 667.100 287.650 667.360 287.970 ;
        RECT 610.980 282.890 611.240 283.210 ;
        RECT 611.040 19.030 611.180 282.890 ;
        RECT 448.600 18.710 448.860 19.030 ;
        RECT 610.980 18.710 611.240 19.030 ;
        RECT 448.660 2.400 448.800 18.710 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 468.810 288.560 469.130 288.620 ;
        RECT 468.810 288.420 480.540 288.560 ;
        RECT 468.810 288.360 469.130 288.420 ;
        RECT 480.400 288.220 480.540 288.420 ;
        RECT 681.790 288.220 682.110 288.280 ;
        RECT 480.400 288.080 682.110 288.220 ;
        RECT 681.790 288.020 682.110 288.080 ;
        RECT 466.510 20.640 466.830 20.700 ;
        RECT 468.810 20.640 469.130 20.700 ;
        RECT 466.510 20.500 469.130 20.640 ;
        RECT 466.510 20.440 466.830 20.500 ;
        RECT 468.810 20.440 469.130 20.500 ;
      LAYER via ;
        RECT 468.840 288.360 469.100 288.620 ;
        RECT 681.820 288.020 682.080 288.280 ;
        RECT 466.540 20.440 466.800 20.700 ;
        RECT 468.840 20.440 469.100 20.700 ;
      LAYER met2 ;
        RECT 681.820 300.000 682.100 304.000 ;
        RECT 468.840 288.330 469.100 288.650 ;
        RECT 468.900 20.730 469.040 288.330 ;
        RECT 681.880 288.310 682.020 300.000 ;
        RECT 681.820 287.990 682.080 288.310 ;
        RECT 466.540 20.410 466.800 20.730 ;
        RECT 468.840 20.410 469.100 20.730 ;
        RECT 466.600 2.400 466.740 20.410 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 631.190 286.860 631.510 286.920 ;
        RECT 696.510 286.860 696.830 286.920 ;
        RECT 631.190 286.720 696.830 286.860 ;
        RECT 631.190 286.660 631.510 286.720 ;
        RECT 696.510 286.660 696.830 286.720 ;
        RECT 484.450 19.280 484.770 19.340 ;
        RECT 631.190 19.280 631.510 19.340 ;
        RECT 484.450 19.140 631.510 19.280 ;
        RECT 484.450 19.080 484.770 19.140 ;
        RECT 631.190 19.080 631.510 19.140 ;
      LAYER via ;
        RECT 631.220 286.660 631.480 286.920 ;
        RECT 696.540 286.660 696.800 286.920 ;
        RECT 484.480 19.080 484.740 19.340 ;
        RECT 631.220 19.080 631.480 19.340 ;
      LAYER met2 ;
        RECT 696.540 300.000 696.820 304.000 ;
        RECT 696.600 286.950 696.740 300.000 ;
        RECT 631.220 286.630 631.480 286.950 ;
        RECT 696.540 286.630 696.800 286.950 ;
        RECT 631.280 19.370 631.420 286.630 ;
        RECT 484.480 19.050 484.740 19.370 ;
        RECT 631.220 19.050 631.480 19.370 ;
        RECT 484.540 2.400 484.680 19.050 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 503.310 289.240 503.630 289.300 ;
        RECT 503.310 289.100 515.960 289.240 ;
        RECT 503.310 289.040 503.630 289.100 ;
        RECT 515.820 288.900 515.960 289.100 ;
        RECT 711.230 288.900 711.550 288.960 ;
        RECT 515.820 288.760 711.550 288.900 ;
        RECT 711.230 288.700 711.550 288.760 ;
      LAYER via ;
        RECT 503.340 289.040 503.600 289.300 ;
        RECT 711.260 288.700 711.520 288.960 ;
      LAYER met2 ;
        RECT 711.260 300.000 711.540 304.000 ;
        RECT 503.340 289.010 503.600 289.330 ;
        RECT 503.400 3.130 503.540 289.010 ;
        RECT 711.320 288.990 711.460 300.000 ;
        RECT 711.260 288.670 711.520 288.990 ;
        RECT 502.480 2.990 503.540 3.130 ;
        RECT 502.480 2.400 502.620 2.990 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 662.545 241.485 662.715 287.555 ;
        RECT 643.225 138.465 643.395 186.235 ;
        RECT 644.605 95.965 644.775 137.955 ;
      LAYER mcon ;
        RECT 662.545 287.385 662.715 287.555 ;
        RECT 643.225 186.065 643.395 186.235 ;
        RECT 644.605 137.785 644.775 137.955 ;
      LAYER met1 ;
        RECT 662.485 287.540 662.775 287.585 ;
        RECT 725.950 287.540 726.270 287.600 ;
        RECT 662.485 287.400 726.270 287.540 ;
        RECT 662.485 287.355 662.775 287.400 ;
        RECT 725.950 287.340 726.270 287.400 ;
        RECT 644.990 241.640 645.310 241.700 ;
        RECT 662.485 241.640 662.775 241.685 ;
        RECT 644.990 241.500 662.775 241.640 ;
        RECT 644.990 241.440 645.310 241.500 ;
        RECT 662.485 241.455 662.775 241.500 ;
        RECT 643.165 186.220 643.455 186.265 ;
        RECT 644.070 186.220 644.390 186.280 ;
        RECT 643.165 186.080 644.390 186.220 ;
        RECT 643.165 186.035 643.455 186.080 ;
        RECT 644.070 186.020 644.390 186.080 ;
        RECT 643.150 138.620 643.470 138.680 ;
        RECT 642.955 138.480 643.470 138.620 ;
        RECT 643.150 138.420 643.470 138.480 ;
        RECT 643.150 137.940 643.470 138.000 ;
        RECT 644.545 137.940 644.835 137.985 ;
        RECT 643.150 137.800 644.835 137.940 ;
        RECT 643.150 137.740 643.470 137.800 ;
        RECT 644.545 137.755 644.835 137.800 ;
        RECT 644.530 96.120 644.850 96.180 ;
        RECT 644.335 95.980 644.850 96.120 ;
        RECT 644.530 95.920 644.850 95.980 ;
        RECT 644.530 62.260 644.850 62.520 ;
        RECT 644.620 61.840 644.760 62.260 ;
        RECT 644.530 61.580 644.850 61.840 ;
        RECT 644.530 16.220 644.850 16.280 ;
        RECT 538.360 16.080 644.850 16.220 ;
        RECT 519.870 15.880 520.190 15.940 ;
        RECT 538.360 15.880 538.500 16.080 ;
        RECT 644.530 16.020 644.850 16.080 ;
        RECT 519.870 15.740 538.500 15.880 ;
        RECT 519.870 15.680 520.190 15.740 ;
      LAYER via ;
        RECT 725.980 287.340 726.240 287.600 ;
        RECT 645.020 241.440 645.280 241.700 ;
        RECT 644.100 186.020 644.360 186.280 ;
        RECT 643.180 138.420 643.440 138.680 ;
        RECT 643.180 137.740 643.440 138.000 ;
        RECT 644.560 95.920 644.820 96.180 ;
        RECT 644.560 62.260 644.820 62.520 ;
        RECT 644.560 61.580 644.820 61.840 ;
        RECT 519.900 15.680 520.160 15.940 ;
        RECT 644.560 16.020 644.820 16.280 ;
      LAYER met2 ;
        RECT 725.980 300.000 726.260 304.000 ;
        RECT 726.040 287.630 726.180 300.000 ;
        RECT 725.980 287.310 726.240 287.630 ;
        RECT 645.020 241.410 645.280 241.730 ;
        RECT 645.080 207.130 645.220 241.410 ;
        RECT 644.160 206.990 645.220 207.130 ;
        RECT 644.160 186.310 644.300 206.990 ;
        RECT 644.100 185.990 644.360 186.310 ;
        RECT 643.180 138.390 643.440 138.710 ;
        RECT 643.240 138.030 643.380 138.390 ;
        RECT 643.180 137.710 643.440 138.030 ;
        RECT 644.560 95.890 644.820 96.210 ;
        RECT 644.620 62.550 644.760 95.890 ;
        RECT 644.560 62.230 644.820 62.550 ;
        RECT 644.560 61.550 644.820 61.870 ;
        RECT 644.620 16.310 644.760 61.550 ;
        RECT 644.560 15.990 644.820 16.310 ;
        RECT 519.900 15.650 520.160 15.970 ;
        RECT 519.960 2.400 520.100 15.650 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 679.490 284.140 679.810 284.200 ;
        RECT 679.490 284.000 713.760 284.140 ;
        RECT 679.490 283.940 679.810 284.000 ;
        RECT 713.620 283.120 713.760 284.000 ;
        RECT 740.670 283.460 740.990 283.520 ;
        RECT 721.440 283.320 740.990 283.460 ;
        RECT 721.440 283.120 721.580 283.320 ;
        RECT 740.670 283.260 740.990 283.320 ;
        RECT 713.620 282.980 721.580 283.120 ;
        RECT 538.270 16.560 538.590 16.620 ;
        RECT 679.490 16.560 679.810 16.620 ;
        RECT 538.270 16.420 679.810 16.560 ;
        RECT 538.270 16.360 538.590 16.420 ;
        RECT 679.490 16.360 679.810 16.420 ;
      LAYER via ;
        RECT 679.520 283.940 679.780 284.200 ;
        RECT 740.700 283.260 740.960 283.520 ;
        RECT 538.300 16.360 538.560 16.620 ;
        RECT 679.520 16.360 679.780 16.620 ;
      LAYER met2 ;
        RECT 740.700 300.000 740.980 304.000 ;
        RECT 679.520 283.910 679.780 284.230 ;
        RECT 679.580 16.650 679.720 283.910 ;
        RECT 740.760 283.550 740.900 300.000 ;
        RECT 740.700 283.230 740.960 283.550 ;
        RECT 538.300 16.330 538.560 16.650 ;
        RECT 679.520 16.330 679.780 16.650 ;
        RECT 538.360 15.540 538.500 16.330 ;
        RECT 537.900 15.400 538.500 15.540 ;
        RECT 537.900 2.400 538.040 15.400 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 713.990 288.900 714.310 288.960 ;
        RECT 755.390 288.900 755.710 288.960 ;
        RECT 713.990 288.760 755.710 288.900 ;
        RECT 713.990 288.700 714.310 288.760 ;
        RECT 755.390 288.700 755.710 288.760 ;
        RECT 555.750 20.300 556.070 20.360 ;
        RECT 713.990 20.300 714.310 20.360 ;
        RECT 555.750 20.160 714.310 20.300 ;
        RECT 555.750 20.100 556.070 20.160 ;
        RECT 713.990 20.100 714.310 20.160 ;
      LAYER via ;
        RECT 714.020 288.700 714.280 288.960 ;
        RECT 755.420 288.700 755.680 288.960 ;
        RECT 555.780 20.100 556.040 20.360 ;
        RECT 714.020 20.100 714.280 20.360 ;
      LAYER met2 ;
        RECT 755.420 300.000 755.700 304.000 ;
        RECT 755.480 288.990 755.620 300.000 ;
        RECT 714.020 288.670 714.280 288.990 ;
        RECT 755.420 288.670 755.680 288.990 ;
        RECT 714.080 20.390 714.220 288.670 ;
        RECT 555.780 20.070 556.040 20.390 ;
        RECT 714.020 20.070 714.280 20.390 ;
        RECT 555.840 2.400 555.980 20.070 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 727.790 283.120 728.110 283.180 ;
        RECT 770.110 283.120 770.430 283.180 ;
        RECT 727.790 282.980 770.430 283.120 ;
        RECT 727.790 282.920 728.110 282.980 ;
        RECT 770.110 282.920 770.430 282.980 ;
        RECT 573.690 16.900 574.010 16.960 ;
        RECT 727.790 16.900 728.110 16.960 ;
        RECT 573.690 16.760 728.110 16.900 ;
        RECT 573.690 16.700 574.010 16.760 ;
        RECT 727.790 16.700 728.110 16.760 ;
      LAYER via ;
        RECT 727.820 282.920 728.080 283.180 ;
        RECT 770.140 282.920 770.400 283.180 ;
        RECT 573.720 16.700 573.980 16.960 ;
        RECT 727.820 16.700 728.080 16.960 ;
      LAYER met2 ;
        RECT 770.140 300.000 770.420 304.000 ;
        RECT 770.200 283.210 770.340 300.000 ;
        RECT 727.820 282.890 728.080 283.210 ;
        RECT 770.140 282.890 770.400 283.210 ;
        RECT 727.880 16.990 728.020 282.890 ;
        RECT 573.720 16.670 573.980 16.990 ;
        RECT 727.820 16.670 728.080 16.990 ;
        RECT 573.780 2.400 573.920 16.670 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 743.505 17.085 743.675 19.635 ;
      LAYER mcon ;
        RECT 743.505 19.465 743.675 19.635 ;
      LAYER met1 ;
        RECT 762.290 289.580 762.610 289.640 ;
        RECT 784.830 289.580 785.150 289.640 ;
        RECT 762.290 289.440 785.150 289.580 ;
        RECT 762.290 289.380 762.610 289.440 ;
        RECT 784.830 289.380 785.150 289.440 ;
        RECT 591.170 19.620 591.490 19.680 ;
        RECT 743.445 19.620 743.735 19.665 ;
        RECT 591.170 19.480 743.735 19.620 ;
        RECT 591.170 19.420 591.490 19.480 ;
        RECT 743.445 19.435 743.735 19.480 ;
        RECT 743.445 17.240 743.735 17.285 ;
        RECT 762.290 17.240 762.610 17.300 ;
        RECT 743.445 17.100 762.610 17.240 ;
        RECT 743.445 17.055 743.735 17.100 ;
        RECT 762.290 17.040 762.610 17.100 ;
      LAYER via ;
        RECT 762.320 289.380 762.580 289.640 ;
        RECT 784.860 289.380 785.120 289.640 ;
        RECT 591.200 19.420 591.460 19.680 ;
        RECT 762.320 17.040 762.580 17.300 ;
      LAYER met2 ;
        RECT 784.860 300.000 785.140 304.000 ;
        RECT 784.920 289.670 785.060 300.000 ;
        RECT 762.320 289.350 762.580 289.670 ;
        RECT 784.860 289.350 785.120 289.670 ;
        RECT 591.200 19.390 591.460 19.710 ;
        RECT 591.260 2.400 591.400 19.390 ;
        RECT 762.380 17.330 762.520 289.350 ;
        RECT 762.320 17.010 762.580 17.330 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 110.085 19.125 110.255 20.655 ;
      LAYER mcon ;
        RECT 110.085 20.485 110.255 20.655 ;
      LAYER met1 ;
        RECT 355.650 286.520 355.970 286.580 ;
        RECT 378.190 286.520 378.510 286.580 ;
        RECT 355.650 286.380 378.510 286.520 ;
        RECT 355.650 286.320 355.970 286.380 ;
        RECT 378.190 286.320 378.510 286.380 ;
        RECT 110.025 20.640 110.315 20.685 ;
        RECT 355.650 20.640 355.970 20.700 ;
        RECT 110.025 20.500 355.970 20.640 ;
        RECT 110.025 20.455 110.315 20.500 ;
        RECT 355.650 20.440 355.970 20.500 ;
        RECT 97.590 19.280 97.910 19.340 ;
        RECT 110.025 19.280 110.315 19.325 ;
        RECT 97.590 19.140 110.315 19.280 ;
        RECT 97.590 19.080 97.910 19.140 ;
        RECT 110.025 19.095 110.315 19.140 ;
      LAYER via ;
        RECT 355.680 286.320 355.940 286.580 ;
        RECT 378.220 286.320 378.480 286.580 ;
        RECT 355.680 20.440 355.940 20.700 ;
        RECT 97.620 19.080 97.880 19.340 ;
      LAYER met2 ;
        RECT 378.220 300.000 378.500 304.000 ;
        RECT 378.280 286.610 378.420 300.000 ;
        RECT 355.680 286.290 355.940 286.610 ;
        RECT 378.220 286.290 378.480 286.610 ;
        RECT 355.740 20.730 355.880 286.290 ;
        RECT 355.680 20.410 355.940 20.730 ;
        RECT 97.620 19.050 97.880 19.370 ;
        RECT 97.680 2.400 97.820 19.050 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 782.990 285.500 783.310 285.560 ;
        RECT 799.090 285.500 799.410 285.560 ;
        RECT 782.990 285.360 799.410 285.500 ;
        RECT 782.990 285.300 783.310 285.360 ;
        RECT 799.090 285.300 799.410 285.360 ;
        RECT 609.110 19.960 609.430 20.020 ;
        RECT 782.990 19.960 783.310 20.020 ;
        RECT 609.110 19.820 783.310 19.960 ;
        RECT 609.110 19.760 609.430 19.820 ;
        RECT 782.990 19.760 783.310 19.820 ;
      LAYER via ;
        RECT 783.020 285.300 783.280 285.560 ;
        RECT 799.120 285.300 799.380 285.560 ;
        RECT 609.140 19.760 609.400 20.020 ;
        RECT 783.020 19.760 783.280 20.020 ;
      LAYER met2 ;
        RECT 799.120 300.000 799.400 304.000 ;
        RECT 799.180 285.590 799.320 300.000 ;
        RECT 783.020 285.270 783.280 285.590 ;
        RECT 799.120 285.270 799.380 285.590 ;
        RECT 783.080 20.050 783.220 285.270 ;
        RECT 609.140 19.730 609.400 20.050 ;
        RECT 783.020 19.730 783.280 20.050 ;
        RECT 609.200 2.400 609.340 19.730 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 783.525 17.765 783.695 19.975 ;
      LAYER mcon ;
        RECT 783.525 19.805 783.695 19.975 ;
      LAYER met1 ;
        RECT 803.690 283.120 804.010 283.180 ;
        RECT 813.810 283.120 814.130 283.180 ;
        RECT 803.690 282.980 814.130 283.120 ;
        RECT 803.690 282.920 804.010 282.980 ;
        RECT 813.810 282.920 814.130 282.980 ;
        RECT 783.465 19.960 783.755 20.005 ;
        RECT 803.690 19.960 804.010 20.020 ;
        RECT 783.465 19.820 804.010 19.960 ;
        RECT 783.465 19.775 783.755 19.820 ;
        RECT 803.690 19.760 804.010 19.820 ;
        RECT 627.050 17.920 627.370 17.980 ;
        RECT 783.465 17.920 783.755 17.965 ;
        RECT 627.050 17.780 783.755 17.920 ;
        RECT 627.050 17.720 627.370 17.780 ;
        RECT 783.465 17.735 783.755 17.780 ;
      LAYER via ;
        RECT 803.720 282.920 803.980 283.180 ;
        RECT 813.840 282.920 814.100 283.180 ;
        RECT 803.720 19.760 803.980 20.020 ;
        RECT 627.080 17.720 627.340 17.980 ;
      LAYER met2 ;
        RECT 813.840 300.000 814.120 304.000 ;
        RECT 813.900 283.210 814.040 300.000 ;
        RECT 803.720 282.890 803.980 283.210 ;
        RECT 813.840 282.890 814.100 283.210 ;
        RECT 803.780 20.050 803.920 282.890 ;
        RECT 803.720 19.730 803.980 20.050 ;
        RECT 627.080 17.690 627.340 18.010 ;
        RECT 627.140 2.400 627.280 17.690 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 355.190 286.860 355.510 286.920 ;
        RECT 397.510 286.860 397.830 286.920 ;
        RECT 355.190 286.720 397.830 286.860 ;
        RECT 355.190 286.660 355.510 286.720 ;
        RECT 397.510 286.660 397.830 286.720 ;
        RECT 351.970 15.540 352.290 15.600 ;
        RECT 355.190 15.540 355.510 15.600 ;
        RECT 351.970 15.400 355.510 15.540 ;
        RECT 351.970 15.340 352.290 15.400 ;
        RECT 355.190 15.340 355.510 15.400 ;
        RECT 121.510 14.860 121.830 14.920 ;
        RECT 351.970 14.860 352.290 14.920 ;
        RECT 121.510 14.720 352.290 14.860 ;
        RECT 121.510 14.660 121.830 14.720 ;
        RECT 351.970 14.660 352.290 14.720 ;
      LAYER via ;
        RECT 355.220 286.660 355.480 286.920 ;
        RECT 397.540 286.660 397.800 286.920 ;
        RECT 352.000 15.340 352.260 15.600 ;
        RECT 355.220 15.340 355.480 15.600 ;
        RECT 121.540 14.660 121.800 14.920 ;
        RECT 352.000 14.660 352.260 14.920 ;
      LAYER met2 ;
        RECT 397.540 300.000 397.820 304.000 ;
        RECT 397.600 286.950 397.740 300.000 ;
        RECT 355.220 286.630 355.480 286.950 ;
        RECT 397.540 286.630 397.800 286.950 ;
        RECT 355.280 15.630 355.420 286.630 ;
        RECT 352.000 15.310 352.260 15.630 ;
        RECT 355.220 15.310 355.480 15.630 ;
        RECT 352.060 14.950 352.200 15.310 ;
        RECT 121.540 14.630 121.800 14.950 ;
        RECT 352.000 14.630 352.260 14.950 ;
        RECT 121.600 2.400 121.740 14.630 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 389.765 287.045 389.935 288.235 ;
      LAYER mcon ;
        RECT 389.765 288.065 389.935 288.235 ;
      LAYER met1 ;
        RECT 150.950 288.220 151.270 288.280 ;
        RECT 389.705 288.220 389.995 288.265 ;
        RECT 150.950 288.080 389.995 288.220 ;
        RECT 150.950 288.020 151.270 288.080 ;
        RECT 389.705 288.035 389.995 288.080 ;
        RECT 417.290 287.540 417.610 287.600 ;
        RECT 395.300 287.400 417.610 287.540 ;
        RECT 389.705 287.200 389.995 287.245 ;
        RECT 395.300 287.200 395.440 287.400 ;
        RECT 417.290 287.340 417.610 287.400 ;
        RECT 389.705 287.060 395.440 287.200 ;
        RECT 389.705 287.015 389.995 287.060 ;
        RECT 145.430 16.900 145.750 16.960 ;
        RECT 150.950 16.900 151.270 16.960 ;
        RECT 145.430 16.760 151.270 16.900 ;
        RECT 145.430 16.700 145.750 16.760 ;
        RECT 150.950 16.700 151.270 16.760 ;
      LAYER via ;
        RECT 150.980 288.020 151.240 288.280 ;
        RECT 417.320 287.340 417.580 287.600 ;
        RECT 145.460 16.700 145.720 16.960 ;
        RECT 150.980 16.700 151.240 16.960 ;
      LAYER met2 ;
        RECT 417.320 300.000 417.600 304.000 ;
        RECT 150.980 287.990 151.240 288.310 ;
        RECT 151.040 16.990 151.180 287.990 ;
        RECT 417.380 287.630 417.520 300.000 ;
        RECT 417.320 287.310 417.580 287.630 ;
        RECT 145.460 16.670 145.720 16.990 ;
        RECT 150.980 16.670 151.240 16.990 ;
        RECT 145.520 2.400 145.660 16.670 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 395.745 282.625 395.915 287.215 ;
        RECT 408.165 287.045 408.335 288.235 ;
        RECT 417.825 287.385 417.995 288.235 ;
      LAYER mcon ;
        RECT 408.165 288.065 408.335 288.235 ;
        RECT 417.825 288.065 417.995 288.235 ;
        RECT 395.745 287.045 395.915 287.215 ;
      LAYER met1 ;
        RECT 408.105 288.220 408.395 288.265 ;
        RECT 417.765 288.220 418.055 288.265 ;
        RECT 408.105 288.080 418.055 288.220 ;
        RECT 408.105 288.035 408.395 288.080 ;
        RECT 417.765 288.035 418.055 288.080 ;
        RECT 417.765 287.540 418.055 287.585 ;
        RECT 432.010 287.540 432.330 287.600 ;
        RECT 417.765 287.400 432.330 287.540 ;
        RECT 417.765 287.355 418.055 287.400 ;
        RECT 432.010 287.340 432.330 287.400 ;
        RECT 395.685 287.200 395.975 287.245 ;
        RECT 408.105 287.200 408.395 287.245 ;
        RECT 395.685 287.060 408.395 287.200 ;
        RECT 395.685 287.015 395.975 287.060 ;
        RECT 408.105 287.015 408.395 287.060 ;
        RECT 389.690 282.780 390.010 282.840 ;
        RECT 395.685 282.780 395.975 282.825 ;
        RECT 389.690 282.640 395.975 282.780 ;
        RECT 389.690 282.580 390.010 282.640 ;
        RECT 395.685 282.595 395.975 282.640 ;
        RECT 386.470 17.920 386.790 17.980 ;
        RECT 389.690 17.920 390.010 17.980 ;
        RECT 386.470 17.780 390.010 17.920 ;
        RECT 386.470 17.720 386.790 17.780 ;
        RECT 389.690 17.720 390.010 17.780 ;
        RECT 163.370 14.520 163.690 14.580 ;
        RECT 386.470 14.520 386.790 14.580 ;
        RECT 163.370 14.380 386.790 14.520 ;
        RECT 163.370 14.320 163.690 14.380 ;
        RECT 386.470 14.320 386.790 14.380 ;
      LAYER via ;
        RECT 432.040 287.340 432.300 287.600 ;
        RECT 389.720 282.580 389.980 282.840 ;
        RECT 386.500 17.720 386.760 17.980 ;
        RECT 389.720 17.720 389.980 17.980 ;
        RECT 163.400 14.320 163.660 14.580 ;
        RECT 386.500 14.320 386.760 14.580 ;
      LAYER met2 ;
        RECT 432.040 300.000 432.320 304.000 ;
        RECT 432.100 287.630 432.240 300.000 ;
        RECT 432.040 287.310 432.300 287.630 ;
        RECT 389.720 282.550 389.980 282.870 ;
        RECT 389.780 18.010 389.920 282.550 ;
        RECT 386.500 17.690 386.760 18.010 ;
        RECT 389.720 17.690 389.980 18.010 ;
        RECT 386.560 14.610 386.700 17.690 ;
        RECT 163.400 14.290 163.660 14.610 ;
        RECT 386.500 14.290 386.760 14.610 ;
        RECT 163.460 2.400 163.600 14.290 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 185.910 285.840 186.230 285.900 ;
        RECT 446.730 285.840 447.050 285.900 ;
        RECT 185.910 285.700 447.050 285.840 ;
        RECT 185.910 285.640 186.230 285.700 ;
        RECT 446.730 285.640 447.050 285.700 ;
        RECT 180.850 16.560 181.170 16.620 ;
        RECT 185.910 16.560 186.230 16.620 ;
        RECT 180.850 16.420 186.230 16.560 ;
        RECT 180.850 16.360 181.170 16.420 ;
        RECT 185.910 16.360 186.230 16.420 ;
      LAYER via ;
        RECT 185.940 285.640 186.200 285.900 ;
        RECT 446.760 285.640 447.020 285.900 ;
        RECT 180.880 16.360 181.140 16.620 ;
        RECT 185.940 16.360 186.200 16.620 ;
      LAYER met2 ;
        RECT 446.760 300.000 447.040 304.000 ;
        RECT 446.820 285.930 446.960 300.000 ;
        RECT 185.940 285.610 186.200 285.930 ;
        RECT 446.760 285.610 447.020 285.930 ;
        RECT 186.000 16.650 186.140 285.610 ;
        RECT 180.880 16.330 181.140 16.650 ;
        RECT 185.940 16.330 186.200 16.650 ;
        RECT 180.940 2.400 181.080 16.330 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 410.390 287.200 410.710 287.260 ;
        RECT 461.450 287.200 461.770 287.260 ;
        RECT 410.390 287.060 461.770 287.200 ;
        RECT 410.390 287.000 410.710 287.060 ;
        RECT 461.450 287.000 461.770 287.060 ;
        RECT 198.790 15.200 199.110 15.260 ;
        RECT 410.390 15.200 410.710 15.260 ;
        RECT 198.790 15.060 410.710 15.200 ;
        RECT 198.790 15.000 199.110 15.060 ;
        RECT 410.390 15.000 410.710 15.060 ;
      LAYER via ;
        RECT 410.420 287.000 410.680 287.260 ;
        RECT 461.480 287.000 461.740 287.260 ;
        RECT 198.820 15.000 199.080 15.260 ;
        RECT 410.420 15.000 410.680 15.260 ;
      LAYER met2 ;
        RECT 461.480 300.000 461.760 304.000 ;
        RECT 461.540 287.290 461.680 300.000 ;
        RECT 410.420 286.970 410.680 287.290 ;
        RECT 461.480 286.970 461.740 287.290 ;
        RECT 410.480 15.290 410.620 286.970 ;
        RECT 198.820 14.970 199.080 15.290 ;
        RECT 410.420 14.970 410.680 15.290 ;
        RECT 198.880 2.400 199.020 14.970 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 220.410 289.580 220.730 289.640 ;
        RECT 476.170 289.580 476.490 289.640 ;
        RECT 220.410 289.440 476.490 289.580 ;
        RECT 220.410 289.380 220.730 289.440 ;
        RECT 476.170 289.380 476.490 289.440 ;
        RECT 216.730 16.560 217.050 16.620 ;
        RECT 220.410 16.560 220.730 16.620 ;
        RECT 216.730 16.420 220.730 16.560 ;
        RECT 216.730 16.360 217.050 16.420 ;
        RECT 220.410 16.360 220.730 16.420 ;
      LAYER via ;
        RECT 220.440 289.380 220.700 289.640 ;
        RECT 476.200 289.380 476.460 289.640 ;
        RECT 216.760 16.360 217.020 16.620 ;
        RECT 220.440 16.360 220.700 16.620 ;
      LAYER met2 ;
        RECT 476.200 300.000 476.480 304.000 ;
        RECT 476.260 289.670 476.400 300.000 ;
        RECT 220.440 289.350 220.700 289.670 ;
        RECT 476.200 289.350 476.460 289.670 ;
        RECT 220.500 16.650 220.640 289.350 ;
        RECT 216.760 16.330 217.020 16.650 ;
        RECT 220.440 16.330 220.700 16.650 ;
        RECT 216.820 2.400 216.960 16.330 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 458.690 284.820 459.010 284.880 ;
        RECT 490.890 284.820 491.210 284.880 ;
        RECT 458.690 284.680 491.210 284.820 ;
        RECT 458.690 284.620 459.010 284.680 ;
        RECT 490.890 284.620 491.210 284.680 ;
        RECT 234.670 14.180 234.990 14.240 ;
        RECT 458.690 14.180 459.010 14.240 ;
        RECT 234.670 14.040 459.010 14.180 ;
        RECT 234.670 13.980 234.990 14.040 ;
        RECT 458.690 13.980 459.010 14.040 ;
      LAYER via ;
        RECT 458.720 284.620 458.980 284.880 ;
        RECT 490.920 284.620 491.180 284.880 ;
        RECT 234.700 13.980 234.960 14.240 ;
        RECT 458.720 13.980 458.980 14.240 ;
      LAYER met2 ;
        RECT 490.920 300.000 491.200 304.000 ;
        RECT 490.980 284.910 491.120 300.000 ;
        RECT 458.720 284.590 458.980 284.910 ;
        RECT 490.920 284.590 491.180 284.910 ;
        RECT 458.780 14.270 458.920 284.590 ;
        RECT 234.700 13.950 234.960 14.270 ;
        RECT 458.720 13.950 458.980 14.270 ;
        RECT 234.760 2.400 234.900 13.950 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 61.710 286.520 62.030 286.580 ;
        RECT 343.690 286.520 344.010 286.580 ;
        RECT 61.710 286.380 344.010 286.520 ;
        RECT 61.710 286.320 62.030 286.380 ;
        RECT 343.690 286.320 344.010 286.380 ;
        RECT 56.190 17.920 56.510 17.980 ;
        RECT 61.710 17.920 62.030 17.980 ;
        RECT 56.190 17.780 62.030 17.920 ;
        RECT 56.190 17.720 56.510 17.780 ;
        RECT 61.710 17.720 62.030 17.780 ;
      LAYER via ;
        RECT 61.740 286.320 62.000 286.580 ;
        RECT 343.720 286.320 343.980 286.580 ;
        RECT 56.220 17.720 56.480 17.980 ;
        RECT 61.740 17.720 62.000 17.980 ;
      LAYER met2 ;
        RECT 343.720 300.000 344.000 304.000 ;
        RECT 343.780 286.610 343.920 300.000 ;
        RECT 61.740 286.290 62.000 286.610 ;
        RECT 343.720 286.290 343.980 286.610 ;
        RECT 61.800 18.010 61.940 286.290 ;
        RECT 56.220 17.690 56.480 18.010 ;
        RECT 61.740 17.690 62.000 18.010 ;
        RECT 56.280 2.400 56.420 17.690 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 130.785 18.105 130.955 19.635 ;
        RECT 180.005 15.725 180.175 18.275 ;
        RECT 226.925 15.725 227.095 18.275 ;
      LAYER mcon ;
        RECT 130.785 19.465 130.955 19.635 ;
        RECT 180.005 18.105 180.175 18.275 ;
        RECT 226.925 18.105 227.095 18.275 ;
      LAYER met1 ;
        RECT 80.110 19.620 80.430 19.680 ;
        RECT 130.725 19.620 131.015 19.665 ;
        RECT 80.110 19.480 131.015 19.620 ;
        RECT 80.110 19.420 80.430 19.480 ;
        RECT 130.725 19.435 131.015 19.480 ;
        RECT 130.725 18.260 131.015 18.305 ;
        RECT 179.945 18.260 180.235 18.305 ;
        RECT 130.725 18.120 180.235 18.260 ;
        RECT 130.725 18.075 131.015 18.120 ;
        RECT 179.945 18.075 180.235 18.120 ;
        RECT 226.865 18.260 227.155 18.305 ;
        RECT 276.530 18.260 276.850 18.320 ;
        RECT 226.865 18.120 276.850 18.260 ;
        RECT 226.865 18.075 227.155 18.120 ;
        RECT 276.530 18.060 276.850 18.120 ;
        RECT 323.450 18.260 323.770 18.320 ;
        RECT 323.450 18.120 341.620 18.260 ;
        RECT 323.450 18.060 323.770 18.120 ;
        RECT 341.480 17.920 341.620 18.120 ;
        RECT 358.870 17.920 359.190 17.980 ;
        RECT 341.480 17.780 359.190 17.920 ;
        RECT 358.870 17.720 359.190 17.780 ;
        RECT 179.945 15.880 180.235 15.925 ;
        RECT 226.865 15.880 227.155 15.925 ;
        RECT 179.945 15.740 227.155 15.880 ;
        RECT 179.945 15.695 180.235 15.740 ;
        RECT 226.865 15.695 227.155 15.740 ;
      LAYER via ;
        RECT 80.140 19.420 80.400 19.680 ;
        RECT 276.560 18.060 276.820 18.320 ;
        RECT 323.480 18.060 323.740 18.320 ;
        RECT 358.900 17.720 359.160 17.980 ;
      LAYER met2 ;
        RECT 363.500 300.290 363.780 304.000 ;
        RECT 358.960 300.150 363.780 300.290 ;
        RECT 80.140 19.390 80.400 19.710 ;
        RECT 80.200 2.400 80.340 19.390 ;
        RECT 276.560 18.205 276.820 18.350 ;
        RECT 323.480 18.205 323.740 18.350 ;
        RECT 276.550 17.835 276.830 18.205 ;
        RECT 323.470 17.835 323.750 18.205 ;
        RECT 358.960 18.010 359.100 300.150 ;
        RECT 363.500 300.000 363.780 300.150 ;
        RECT 358.900 17.690 359.160 18.010 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 276.550 17.880 276.830 18.160 ;
        RECT 323.470 17.880 323.750 18.160 ;
      LAYER met3 ;
        RECT 276.525 18.170 276.855 18.185 ;
        RECT 323.445 18.170 323.775 18.185 ;
        RECT 276.525 17.870 323.775 18.170 ;
        RECT 276.525 17.855 276.855 17.870 ;
        RECT 323.445 17.855 323.775 17.870 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 287.200 109.870 287.260 ;
        RECT 382.790 287.200 383.110 287.260 ;
        RECT 109.550 287.060 383.110 287.200 ;
        RECT 109.550 287.000 109.870 287.060 ;
        RECT 382.790 287.000 383.110 287.060 ;
        RECT 103.570 20.640 103.890 20.700 ;
        RECT 109.550 20.640 109.870 20.700 ;
        RECT 103.570 20.500 109.870 20.640 ;
        RECT 103.570 20.440 103.890 20.500 ;
        RECT 109.550 20.440 109.870 20.500 ;
      LAYER via ;
        RECT 109.580 287.000 109.840 287.260 ;
        RECT 382.820 287.000 383.080 287.260 ;
        RECT 103.600 20.440 103.860 20.700 ;
        RECT 109.580 20.440 109.840 20.700 ;
      LAYER met2 ;
        RECT 382.820 300.000 383.100 304.000 ;
        RECT 382.880 287.290 383.020 300.000 ;
        RECT 109.580 286.970 109.840 287.290 ;
        RECT 382.820 286.970 383.080 287.290 ;
        RECT 109.640 20.730 109.780 286.970 ;
        RECT 103.600 20.410 103.860 20.730 ;
        RECT 109.580 20.410 109.840 20.730 ;
        RECT 103.660 2.400 103.800 20.410 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 127.490 18.940 127.810 19.000 ;
        RECT 400.270 18.940 400.590 19.000 ;
        RECT 127.490 18.800 400.590 18.940 ;
        RECT 127.490 18.740 127.810 18.800 ;
        RECT 400.270 18.740 400.590 18.800 ;
      LAYER via ;
        RECT 127.520 18.740 127.780 19.000 ;
        RECT 400.300 18.740 400.560 19.000 ;
      LAYER met2 ;
        RECT 402.600 300.290 402.880 304.000 ;
        RECT 400.360 300.150 402.880 300.290 ;
        RECT 400.360 19.030 400.500 300.150 ;
        RECT 402.600 300.000 402.880 300.150 ;
        RECT 127.520 18.710 127.780 19.030 ;
        RECT 400.300 18.710 400.560 19.030 ;
        RECT 127.580 2.400 127.720 18.710 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.290 2.960 26.610 3.020 ;
        RECT 27.210 2.960 27.530 3.020 ;
        RECT 26.290 2.820 27.530 2.960 ;
        RECT 26.290 2.760 26.610 2.820 ;
        RECT 27.210 2.760 27.530 2.820 ;
      LAYER via ;
        RECT 26.320 2.760 26.580 3.020 ;
        RECT 27.240 2.760 27.500 3.020 ;
      LAYER met2 ;
        RECT 319.340 300.000 319.620 304.000 ;
        RECT 319.400 286.125 319.540 300.000 ;
        RECT 27.230 285.755 27.510 286.125 ;
        RECT 319.330 285.755 319.610 286.125 ;
        RECT 27.300 3.050 27.440 285.755 ;
        RECT 26.320 2.730 26.580 3.050 ;
        RECT 27.240 2.730 27.500 3.050 ;
        RECT 26.380 2.400 26.520 2.730 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 27.230 285.800 27.510 286.080 ;
        RECT 319.330 285.800 319.610 286.080 ;
      LAYER met3 ;
        RECT 27.205 286.090 27.535 286.105 ;
        RECT 319.305 286.090 319.635 286.105 ;
        RECT 27.205 285.790 319.635 286.090 ;
        RECT 27.205 285.775 27.535 285.790 ;
        RECT 319.305 285.775 319.635 285.790 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.270 17.240 32.590 17.300 ;
        RECT 325.290 17.240 325.610 17.300 ;
        RECT 32.270 17.100 325.610 17.240 ;
        RECT 32.270 17.040 32.590 17.100 ;
        RECT 325.290 17.040 325.610 17.100 ;
      LAYER via ;
        RECT 32.300 17.040 32.560 17.300 ;
        RECT 325.320 17.040 325.580 17.300 ;
      LAYER met2 ;
        RECT 324.400 300.290 324.680 304.000 ;
        RECT 324.400 300.150 325.520 300.290 ;
        RECT 324.400 300.000 324.680 300.150 ;
        RECT 325.380 17.330 325.520 300.150 ;
        RECT 32.300 17.010 32.560 17.330 ;
        RECT 325.320 17.010 325.580 17.330 ;
        RECT 32.360 2.400 32.500 17.010 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 364.020 -9.320 367.020 3529.000 ;
        RECT 544.020 -9.320 547.020 3529.000 ;
        RECT 724.020 -9.320 727.020 3529.000 ;
        RECT 904.020 -9.320 907.020 3529.000 ;
        RECT 1084.020 -9.320 1087.020 3529.000 ;
        RECT 1264.020 -9.320 1267.020 3529.000 ;
        RECT 1444.020 -9.320 1447.020 3529.000 ;
        RECT 1624.020 -9.320 1627.020 3529.000 ;
        RECT 1804.020 -9.320 1807.020 3529.000 ;
        RECT 1984.020 -9.320 1987.020 3529.000 ;
        RECT 2164.020 -9.320 2167.020 3529.000 ;
        RECT 2344.020 -9.320 2347.020 3529.000 ;
        RECT 2524.020 -9.320 2527.020 3529.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 454.020 -9.320 457.020 3529.000 ;
        RECT 634.020 -9.320 637.020 3529.000 ;
        RECT 814.020 -9.320 817.020 3529.000 ;
        RECT 994.020 -9.320 997.020 3529.000 ;
        RECT 1174.020 -9.320 1177.020 3529.000 ;
        RECT 1354.020 -9.320 1357.020 3529.000 ;
        RECT 1534.020 -9.320 1537.020 3529.000 ;
        RECT 1714.020 -9.320 1717.020 3529.000 ;
        RECT 1894.020 -9.320 1897.020 3529.000 ;
        RECT 2074.020 -9.320 2077.020 3529.000 ;
        RECT 2254.020 -9.320 2257.020 3529.000 ;
        RECT 2434.020 -9.320 2437.020 3529.000 ;
        RECT 2614.020 -9.320 2617.020 3529.000 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 382.020 -18.720 385.020 3538.400 ;
        RECT 562.020 -18.720 565.020 3538.400 ;
        RECT 742.020 -18.720 745.020 3538.400 ;
        RECT 922.020 -18.720 925.020 3538.400 ;
        RECT 1102.020 -18.720 1105.020 3538.400 ;
        RECT 1282.020 -18.720 1285.020 3538.400 ;
        RECT 1462.020 -18.720 1465.020 3538.400 ;
        RECT 1642.020 -18.720 1645.020 3538.400 ;
        RECT 1822.020 -18.720 1825.020 3538.400 ;
        RECT 2002.020 -18.720 2005.020 3538.400 ;
        RECT 2182.020 -18.720 2185.020 3538.400 ;
        RECT 2362.020 -18.720 2365.020 3538.400 ;
        RECT 2542.020 -18.720 2545.020 3538.400 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1282.930 2009.090 1284.110 2010.270 ;
        RECT 1282.930 2007.490 1284.110 2008.670 ;
        RECT 1282.930 1829.090 1284.110 1830.270 ;
        RECT 1282.930 1827.490 1284.110 1828.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 1282.020 2010.380 1285.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 1282.020 2007.370 1285.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 1282.020 1830.380 1285.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 1282.020 1827.370 1285.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 292.020 -18.720 295.020 3538.400 ;
        RECT 472.020 -18.720 475.020 3538.400 ;
        RECT 652.020 -18.720 655.020 3538.400 ;
        RECT 832.020 -18.720 835.020 3538.400 ;
        RECT 1012.020 -18.720 1015.020 3538.400 ;
        RECT 1192.020 -18.720 1195.020 3538.400 ;
        RECT 1372.020 -18.720 1375.020 3538.400 ;
        RECT 1552.020 -18.720 1555.020 3538.400 ;
        RECT 1732.020 -18.720 1735.020 3538.400 ;
        RECT 1912.020 -18.720 1915.020 3538.400 ;
        RECT 2092.020 -18.720 2095.020 3538.400 ;
        RECT 2272.020 -18.720 2275.020 3538.400 ;
        RECT 2452.020 -18.720 2455.020 3538.400 ;
        RECT 2632.020 -18.720 2635.020 3538.400 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 400.020 -28.120 403.020 3547.800 ;
        RECT 580.020 -28.120 583.020 3547.800 ;
        RECT 760.020 -28.120 763.020 3547.800 ;
        RECT 940.020 -28.120 943.020 3547.800 ;
        RECT 1120.020 -28.120 1123.020 3547.800 ;
        RECT 1300.020 -28.120 1303.020 3547.800 ;
        RECT 1480.020 -28.120 1483.020 3547.800 ;
        RECT 1660.020 -28.120 1663.020 3547.800 ;
        RECT 1840.020 -28.120 1843.020 3547.800 ;
        RECT 2020.020 -28.120 2023.020 3547.800 ;
        RECT 2200.020 -28.120 2203.020 3547.800 ;
        RECT 2380.020 -28.120 2383.020 3547.800 ;
        RECT 2560.020 -28.120 2563.020 3547.800 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1300.930 2027.090 1302.110 2028.270 ;
        RECT 1300.930 2025.490 1302.110 2026.670 ;
        RECT 1300.930 1847.090 1302.110 1848.270 ;
        RECT 1300.930 1845.490 1302.110 1846.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 1300.020 2028.380 1303.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 1300.020 2025.370 1303.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 1300.020 1848.380 1303.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 1300.020 1845.370 1303.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 310.020 -28.120 313.020 3547.800 ;
        RECT 490.020 -28.120 493.020 3547.800 ;
        RECT 670.020 -28.120 673.020 3547.800 ;
        RECT 850.020 -28.120 853.020 3547.800 ;
        RECT 1030.020 -28.120 1033.020 3547.800 ;
        RECT 1210.020 -28.120 1213.020 3547.800 ;
        RECT 1390.020 -28.120 1393.020 3547.800 ;
        RECT 1570.020 -28.120 1573.020 3547.800 ;
        RECT 1750.020 -28.120 1753.020 3547.800 ;
        RECT 1930.020 -28.120 1933.020 3547.800 ;
        RECT 2110.020 -28.120 2113.020 3547.800 ;
        RECT 2290.020 -28.120 2293.020 3547.800 ;
        RECT 2470.020 -28.120 2473.020 3547.800 ;
        RECT 2650.020 -28.120 2653.020 3547.800 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 1930.930 1757.090 1932.110 1758.270 ;
        RECT 1930.930 1755.490 1932.110 1756.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 1930.020 1758.380 1933.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 1930.020 1755.370 1933.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 418.020 -37.520 421.020 3557.200 ;
        RECT 598.020 -37.520 601.020 3557.200 ;
        RECT 778.020 -37.520 781.020 3557.200 ;
        RECT 958.020 -37.520 961.020 3557.200 ;
        RECT 1138.020 -37.520 1141.020 3557.200 ;
        RECT 1318.020 -37.520 1321.020 3557.200 ;
        RECT 1498.020 -37.520 1501.020 3557.200 ;
        RECT 1678.020 -37.520 1681.020 3557.200 ;
        RECT 1858.020 -37.520 1861.020 3557.200 ;
        RECT 2038.020 -37.520 2041.020 3557.200 ;
        RECT 2218.020 -37.520 2221.020 3557.200 ;
        RECT 2398.020 -37.520 2401.020 3557.200 ;
        RECT 2578.020 -37.520 2581.020 3557.200 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1318.930 2045.090 1320.110 2046.270 ;
        RECT 1318.930 2043.490 1320.110 2044.670 ;
        RECT 1318.930 1865.090 1320.110 1866.270 ;
        RECT 1318.930 1863.490 1320.110 1864.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 1318.020 2046.380 1321.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 1318.020 2043.370 1321.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 1318.020 1866.380 1321.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 1318.020 1863.370 1321.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 328.020 -37.520 331.020 3557.200 ;
        RECT 508.020 -37.520 511.020 3557.200 ;
        RECT 688.020 -37.520 691.020 3557.200 ;
        RECT 868.020 -37.520 871.020 3557.200 ;
        RECT 1048.020 -37.520 1051.020 3557.200 ;
        RECT 1228.020 -37.520 1231.020 3557.200 ;
        RECT 1408.020 -37.520 1411.020 3557.200 ;
        RECT 1588.020 -37.520 1591.020 3557.200 ;
        RECT 1768.020 -37.520 1771.020 3557.200 ;
        RECT 1948.020 -37.520 1951.020 3557.200 ;
        RECT 2128.020 -37.520 2131.020 3557.200 ;
        RECT 2308.020 -37.520 2311.020 3557.200 ;
        RECT 2488.020 -37.520 2491.020 3557.200 ;
        RECT 2668.020 -37.520 2671.020 3557.200 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 1948.930 1775.090 1950.110 1776.270 ;
        RECT 1948.930 1773.490 1950.110 1774.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 1948.020 1776.380 1951.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 1948.020 1773.370 1951.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 303.150 310.795 2691.930 3286.645 ;
      LAYER met1 ;
        RECT 300.000 304.460 2691.930 3292.300 ;
      LAYER met2 ;
        RECT 300.030 3295.720 307.560 3296.000 ;
        RECT 308.400 3295.720 328.260 3296.000 ;
        RECT 329.100 3295.720 349.420 3296.000 ;
        RECT 350.260 3295.720 370.580 3296.000 ;
        RECT 371.420 3295.720 391.740 3296.000 ;
        RECT 392.580 3295.720 412.440 3296.000 ;
        RECT 413.280 3295.720 433.600 3296.000 ;
        RECT 434.440 3295.720 454.760 3296.000 ;
        RECT 455.600 3295.720 475.920 3296.000 ;
        RECT 476.760 3295.720 496.620 3296.000 ;
        RECT 497.460 3295.720 517.780 3296.000 ;
        RECT 518.620 3295.720 538.940 3296.000 ;
        RECT 539.780 3295.720 560.100 3296.000 ;
        RECT 560.940 3295.720 580.800 3296.000 ;
        RECT 581.640 3295.720 601.960 3296.000 ;
        RECT 602.800 3295.720 623.120 3296.000 ;
        RECT 623.960 3295.720 644.280 3296.000 ;
        RECT 645.120 3295.720 664.980 3296.000 ;
        RECT 665.820 3295.720 686.140 3296.000 ;
        RECT 686.980 3295.720 707.300 3296.000 ;
        RECT 708.140 3295.720 728.460 3296.000 ;
        RECT 729.300 3295.720 749.620 3296.000 ;
        RECT 750.460 3295.720 770.320 3296.000 ;
        RECT 771.160 3295.720 791.480 3296.000 ;
        RECT 792.320 3295.720 812.640 3296.000 ;
        RECT 813.480 3295.720 833.800 3296.000 ;
        RECT 834.640 3295.720 854.500 3296.000 ;
        RECT 855.340 3295.720 875.660 3296.000 ;
        RECT 876.500 3295.720 896.820 3296.000 ;
        RECT 897.660 3295.720 917.980 3296.000 ;
        RECT 918.820 3295.720 938.680 3296.000 ;
        RECT 939.520 3295.720 959.840 3296.000 ;
        RECT 960.680 3295.720 981.000 3296.000 ;
        RECT 981.840 3295.720 1002.160 3296.000 ;
        RECT 1003.000 3295.720 1022.860 3296.000 ;
        RECT 1023.700 3295.720 1044.020 3296.000 ;
        RECT 1044.860 3295.720 1065.180 3296.000 ;
        RECT 1066.020 3295.720 1086.340 3296.000 ;
        RECT 1087.180 3295.720 1107.500 3296.000 ;
        RECT 1108.340 3295.720 1128.200 3296.000 ;
        RECT 1129.040 3295.720 1149.360 3296.000 ;
        RECT 1150.200 3295.720 1170.520 3296.000 ;
        RECT 1171.360 3295.720 1191.680 3296.000 ;
        RECT 1192.520 3295.720 1212.380 3296.000 ;
        RECT 1213.220 3295.720 1233.540 3296.000 ;
        RECT 1234.380 3295.720 1254.700 3296.000 ;
        RECT 1255.540 3295.720 1275.860 3296.000 ;
        RECT 1276.700 3295.720 1296.560 3296.000 ;
        RECT 1297.400 3295.720 1317.720 3296.000 ;
        RECT 1318.560 3295.720 1338.880 3296.000 ;
        RECT 1339.720 3295.720 1360.040 3296.000 ;
        RECT 1360.880 3295.720 1380.740 3296.000 ;
        RECT 1381.580 3295.720 1401.900 3296.000 ;
        RECT 1402.740 3295.720 1423.060 3296.000 ;
        RECT 1423.900 3295.720 1444.220 3296.000 ;
        RECT 1445.060 3295.720 1464.920 3296.000 ;
        RECT 1465.760 3295.720 1486.080 3296.000 ;
        RECT 1486.920 3295.720 1507.240 3296.000 ;
        RECT 1508.080 3295.720 1528.400 3296.000 ;
        RECT 1529.240 3295.720 1549.560 3296.000 ;
        RECT 1550.400 3295.720 1570.260 3296.000 ;
        RECT 1571.100 3295.720 1591.420 3296.000 ;
        RECT 1592.260 3295.720 1612.580 3296.000 ;
        RECT 1613.420 3295.720 1633.740 3296.000 ;
        RECT 1634.580 3295.720 1654.440 3296.000 ;
        RECT 1655.280 3295.720 1675.600 3296.000 ;
        RECT 1676.440 3295.720 1696.760 3296.000 ;
        RECT 1697.600 3295.720 1717.920 3296.000 ;
        RECT 1718.760 3295.720 1738.620 3296.000 ;
        RECT 1739.460 3295.720 1759.780 3296.000 ;
        RECT 1760.620 3295.720 1780.940 3296.000 ;
        RECT 1781.780 3295.720 1802.100 3296.000 ;
        RECT 1802.940 3295.720 1822.800 3296.000 ;
        RECT 1823.640 3295.720 1843.960 3296.000 ;
        RECT 1844.800 3295.720 1865.120 3296.000 ;
        RECT 1865.960 3295.720 1886.280 3296.000 ;
        RECT 1887.120 3295.720 1907.440 3296.000 ;
        RECT 1908.280 3295.720 1928.140 3296.000 ;
        RECT 1928.980 3295.720 1949.300 3296.000 ;
        RECT 1950.140 3295.720 1970.460 3296.000 ;
        RECT 1971.300 3295.720 1991.620 3296.000 ;
        RECT 1992.460 3295.720 2012.320 3296.000 ;
        RECT 2013.160 3295.720 2033.480 3296.000 ;
        RECT 2034.320 3295.720 2054.640 3296.000 ;
        RECT 2055.480 3295.720 2075.800 3296.000 ;
        RECT 2076.640 3295.720 2096.500 3296.000 ;
        RECT 2097.340 3295.720 2117.660 3296.000 ;
        RECT 2118.500 3295.720 2138.820 3296.000 ;
        RECT 2139.660 3295.720 2159.980 3296.000 ;
        RECT 2160.820 3295.720 2180.680 3296.000 ;
        RECT 2181.520 3295.720 2201.840 3296.000 ;
        RECT 2202.680 3295.720 2223.000 3296.000 ;
        RECT 2223.840 3295.720 2244.160 3296.000 ;
        RECT 2245.000 3295.720 2264.860 3296.000 ;
        RECT 2265.700 3295.720 2286.020 3296.000 ;
        RECT 2286.860 3295.720 2307.180 3296.000 ;
        RECT 2308.020 3295.720 2328.340 3296.000 ;
        RECT 2329.180 3295.720 2349.500 3296.000 ;
        RECT 2350.340 3295.720 2370.200 3296.000 ;
        RECT 2371.040 3295.720 2391.360 3296.000 ;
        RECT 2392.200 3295.720 2412.520 3296.000 ;
        RECT 2413.360 3295.720 2433.680 3296.000 ;
        RECT 2434.520 3295.720 2454.380 3296.000 ;
        RECT 2455.220 3295.720 2475.540 3296.000 ;
        RECT 2476.380 3295.720 2496.700 3296.000 ;
        RECT 2497.540 3295.720 2517.860 3296.000 ;
        RECT 2518.700 3295.720 2538.560 3296.000 ;
        RECT 2539.400 3295.720 2559.720 3296.000 ;
        RECT 2560.560 3295.720 2580.880 3296.000 ;
        RECT 2581.720 3295.720 2602.040 3296.000 ;
        RECT 2602.880 3295.720 2622.740 3296.000 ;
        RECT 2623.580 3295.720 2643.900 3296.000 ;
        RECT 2644.740 3295.720 2665.060 3296.000 ;
        RECT 2665.900 3295.720 2686.220 3296.000 ;
        RECT 2687.060 3295.720 2689.990 3296.000 ;
        RECT 300.030 304.280 2689.990 3295.720 ;
        RECT 300.580 304.000 304.340 304.280 ;
        RECT 305.180 304.000 309.400 304.280 ;
        RECT 310.240 304.000 314.000 304.280 ;
        RECT 314.840 304.000 319.060 304.280 ;
        RECT 319.900 304.000 324.120 304.280 ;
        RECT 324.960 304.000 328.720 304.280 ;
        RECT 329.560 304.000 333.780 304.280 ;
        RECT 334.620 304.000 338.840 304.280 ;
        RECT 339.680 304.000 343.440 304.280 ;
        RECT 344.280 304.000 348.500 304.280 ;
        RECT 349.340 304.000 353.560 304.280 ;
        RECT 354.400 304.000 358.160 304.280 ;
        RECT 359.000 304.000 363.220 304.280 ;
        RECT 364.060 304.000 368.280 304.280 ;
        RECT 369.120 304.000 372.880 304.280 ;
        RECT 373.720 304.000 377.940 304.280 ;
        RECT 378.780 304.000 382.540 304.280 ;
        RECT 383.380 304.000 387.600 304.280 ;
        RECT 388.440 304.000 392.660 304.280 ;
        RECT 393.500 304.000 397.260 304.280 ;
        RECT 398.100 304.000 402.320 304.280 ;
        RECT 403.160 304.000 407.380 304.280 ;
        RECT 408.220 304.000 411.980 304.280 ;
        RECT 412.820 304.000 417.040 304.280 ;
        RECT 417.880 304.000 422.100 304.280 ;
        RECT 422.940 304.000 426.700 304.280 ;
        RECT 427.540 304.000 431.760 304.280 ;
        RECT 432.600 304.000 436.820 304.280 ;
        RECT 437.660 304.000 441.420 304.280 ;
        RECT 442.260 304.000 446.480 304.280 ;
        RECT 447.320 304.000 451.540 304.280 ;
        RECT 452.380 304.000 456.140 304.280 ;
        RECT 456.980 304.000 461.200 304.280 ;
        RECT 462.040 304.000 465.800 304.280 ;
        RECT 466.640 304.000 470.860 304.280 ;
        RECT 471.700 304.000 475.920 304.280 ;
        RECT 476.760 304.000 480.520 304.280 ;
        RECT 481.360 304.000 485.580 304.280 ;
        RECT 486.420 304.000 490.640 304.280 ;
        RECT 491.480 304.000 495.240 304.280 ;
        RECT 496.080 304.000 500.300 304.280 ;
        RECT 501.140 304.000 505.360 304.280 ;
        RECT 506.200 304.000 509.960 304.280 ;
        RECT 510.800 304.000 515.020 304.280 ;
        RECT 515.860 304.000 520.080 304.280 ;
        RECT 520.920 304.000 524.680 304.280 ;
        RECT 525.520 304.000 529.740 304.280 ;
        RECT 530.580 304.000 534.800 304.280 ;
        RECT 535.640 304.000 539.400 304.280 ;
        RECT 540.240 304.000 544.460 304.280 ;
        RECT 545.300 304.000 549.060 304.280 ;
        RECT 549.900 304.000 554.120 304.280 ;
        RECT 554.960 304.000 559.180 304.280 ;
        RECT 560.020 304.000 563.780 304.280 ;
        RECT 564.620 304.000 568.840 304.280 ;
        RECT 569.680 304.000 573.900 304.280 ;
        RECT 574.740 304.000 578.500 304.280 ;
        RECT 579.340 304.000 583.560 304.280 ;
        RECT 584.400 304.000 588.620 304.280 ;
        RECT 589.460 304.000 593.220 304.280 ;
        RECT 594.060 304.000 598.280 304.280 ;
        RECT 599.120 304.000 603.340 304.280 ;
        RECT 604.180 304.000 607.940 304.280 ;
        RECT 608.780 304.000 613.000 304.280 ;
        RECT 613.840 304.000 618.060 304.280 ;
        RECT 618.900 304.000 622.660 304.280 ;
        RECT 623.500 304.000 627.720 304.280 ;
        RECT 628.560 304.000 632.320 304.280 ;
        RECT 633.160 304.000 637.380 304.280 ;
        RECT 638.220 304.000 642.440 304.280 ;
        RECT 643.280 304.000 647.040 304.280 ;
        RECT 647.880 304.000 652.100 304.280 ;
        RECT 652.940 304.000 657.160 304.280 ;
        RECT 658.000 304.000 661.760 304.280 ;
        RECT 662.600 304.000 666.820 304.280 ;
        RECT 667.660 304.000 671.880 304.280 ;
        RECT 672.720 304.000 676.480 304.280 ;
        RECT 677.320 304.000 681.540 304.280 ;
        RECT 682.380 304.000 686.600 304.280 ;
        RECT 687.440 304.000 691.200 304.280 ;
        RECT 692.040 304.000 696.260 304.280 ;
        RECT 697.100 304.000 701.320 304.280 ;
        RECT 702.160 304.000 705.920 304.280 ;
        RECT 706.760 304.000 710.980 304.280 ;
        RECT 711.820 304.000 715.580 304.280 ;
        RECT 716.420 304.000 720.640 304.280 ;
        RECT 721.480 304.000 725.700 304.280 ;
        RECT 726.540 304.000 730.300 304.280 ;
        RECT 731.140 304.000 735.360 304.280 ;
        RECT 736.200 304.000 740.420 304.280 ;
        RECT 741.260 304.000 745.020 304.280 ;
        RECT 745.860 304.000 750.080 304.280 ;
        RECT 750.920 304.000 755.140 304.280 ;
        RECT 755.980 304.000 759.740 304.280 ;
        RECT 760.580 304.000 764.800 304.280 ;
        RECT 765.640 304.000 769.860 304.280 ;
        RECT 770.700 304.000 774.460 304.280 ;
        RECT 775.300 304.000 779.520 304.280 ;
        RECT 780.360 304.000 784.580 304.280 ;
        RECT 785.420 304.000 789.180 304.280 ;
        RECT 790.020 304.000 794.240 304.280 ;
        RECT 795.080 304.000 798.840 304.280 ;
        RECT 799.680 304.000 803.900 304.280 ;
        RECT 804.740 304.000 808.960 304.280 ;
        RECT 809.800 304.000 813.560 304.280 ;
        RECT 814.400 304.000 818.620 304.280 ;
        RECT 819.460 304.000 823.680 304.280 ;
        RECT 824.520 304.000 828.280 304.280 ;
        RECT 829.120 304.000 833.340 304.280 ;
        RECT 834.180 304.000 838.400 304.280 ;
        RECT 839.240 304.000 843.000 304.280 ;
        RECT 843.840 304.000 848.060 304.280 ;
        RECT 848.900 304.000 853.120 304.280 ;
        RECT 853.960 304.000 857.720 304.280 ;
        RECT 858.560 304.000 862.780 304.280 ;
        RECT 863.620 304.000 867.840 304.280 ;
        RECT 868.680 304.000 872.440 304.280 ;
        RECT 873.280 304.000 877.500 304.280 ;
        RECT 878.340 304.000 882.100 304.280 ;
        RECT 882.940 304.000 887.160 304.280 ;
        RECT 888.000 304.000 892.220 304.280 ;
        RECT 893.060 304.000 896.820 304.280 ;
        RECT 897.660 304.000 901.880 304.280 ;
        RECT 902.720 304.000 906.940 304.280 ;
        RECT 907.780 304.000 911.540 304.280 ;
        RECT 912.380 304.000 916.600 304.280 ;
        RECT 917.440 304.000 921.660 304.280 ;
        RECT 922.500 304.000 926.260 304.280 ;
        RECT 927.100 304.000 931.320 304.280 ;
        RECT 932.160 304.000 936.380 304.280 ;
        RECT 937.220 304.000 940.980 304.280 ;
        RECT 941.820 304.000 946.040 304.280 ;
        RECT 946.880 304.000 951.100 304.280 ;
        RECT 951.940 304.000 955.700 304.280 ;
        RECT 956.540 304.000 960.760 304.280 ;
        RECT 961.600 304.000 965.360 304.280 ;
        RECT 966.200 304.000 970.420 304.280 ;
        RECT 971.260 304.000 975.480 304.280 ;
        RECT 976.320 304.000 980.080 304.280 ;
        RECT 980.920 304.000 985.140 304.280 ;
        RECT 985.980 304.000 990.200 304.280 ;
        RECT 991.040 304.000 994.800 304.280 ;
        RECT 995.640 304.000 999.860 304.280 ;
        RECT 1000.700 304.000 1004.920 304.280 ;
        RECT 1005.760 304.000 1009.520 304.280 ;
        RECT 1010.360 304.000 1014.580 304.280 ;
        RECT 1015.420 304.000 1019.640 304.280 ;
        RECT 1020.480 304.000 1024.240 304.280 ;
        RECT 1025.080 304.000 1029.300 304.280 ;
        RECT 1030.140 304.000 1034.360 304.280 ;
        RECT 1035.200 304.000 1038.960 304.280 ;
        RECT 1039.800 304.000 1044.020 304.280 ;
        RECT 1044.860 304.000 1048.620 304.280 ;
        RECT 1049.460 304.000 1053.680 304.280 ;
        RECT 1054.520 304.000 1058.740 304.280 ;
        RECT 1059.580 304.000 1063.340 304.280 ;
        RECT 1064.180 304.000 1068.400 304.280 ;
        RECT 1069.240 304.000 1073.460 304.280 ;
        RECT 1074.300 304.000 1078.060 304.280 ;
        RECT 1078.900 304.000 1083.120 304.280 ;
        RECT 1083.960 304.000 1088.180 304.280 ;
        RECT 1089.020 304.000 1092.780 304.280 ;
        RECT 1093.620 304.000 1097.840 304.280 ;
        RECT 1098.680 304.000 1102.900 304.280 ;
        RECT 1103.740 304.000 1107.500 304.280 ;
        RECT 1108.340 304.000 1112.560 304.280 ;
        RECT 1113.400 304.000 1117.620 304.280 ;
        RECT 1118.460 304.000 1122.220 304.280 ;
        RECT 1123.060 304.000 1127.280 304.280 ;
        RECT 1128.120 304.000 1131.880 304.280 ;
        RECT 1132.720 304.000 1136.940 304.280 ;
        RECT 1137.780 304.000 1142.000 304.280 ;
        RECT 1142.840 304.000 1146.600 304.280 ;
        RECT 1147.440 304.000 1151.660 304.280 ;
        RECT 1152.500 304.000 1156.720 304.280 ;
        RECT 1157.560 304.000 1161.320 304.280 ;
        RECT 1162.160 304.000 1166.380 304.280 ;
        RECT 1167.220 304.000 1171.440 304.280 ;
        RECT 1172.280 304.000 1176.040 304.280 ;
        RECT 1176.880 304.000 1181.100 304.280 ;
        RECT 1181.940 304.000 1186.160 304.280 ;
        RECT 1187.000 304.000 1190.760 304.280 ;
        RECT 1191.600 304.000 1195.820 304.280 ;
        RECT 1196.660 304.000 1200.880 304.280 ;
        RECT 1201.720 304.000 1205.480 304.280 ;
        RECT 1206.320 304.000 1210.540 304.280 ;
        RECT 1211.380 304.000 1215.140 304.280 ;
        RECT 1215.980 304.000 1220.200 304.280 ;
        RECT 1221.040 304.000 1225.260 304.280 ;
        RECT 1226.100 304.000 1229.860 304.280 ;
        RECT 1230.700 304.000 1234.920 304.280 ;
        RECT 1235.760 304.000 1239.980 304.280 ;
        RECT 1240.820 304.000 1244.580 304.280 ;
        RECT 1245.420 304.000 1249.640 304.280 ;
        RECT 1250.480 304.000 1254.700 304.280 ;
        RECT 1255.540 304.000 1259.300 304.280 ;
        RECT 1260.140 304.000 1264.360 304.280 ;
        RECT 1265.200 304.000 1269.420 304.280 ;
        RECT 1270.260 304.000 1274.020 304.280 ;
        RECT 1274.860 304.000 1279.080 304.280 ;
        RECT 1279.920 304.000 1284.140 304.280 ;
        RECT 1284.980 304.000 1288.740 304.280 ;
        RECT 1289.580 304.000 1293.800 304.280 ;
        RECT 1294.640 304.000 1298.400 304.280 ;
        RECT 1299.240 304.000 1303.460 304.280 ;
        RECT 1304.300 304.000 1308.520 304.280 ;
        RECT 1309.360 304.000 1313.120 304.280 ;
        RECT 1313.960 304.000 1318.180 304.280 ;
        RECT 1319.020 304.000 1323.240 304.280 ;
        RECT 1324.080 304.000 1327.840 304.280 ;
        RECT 1328.680 304.000 1332.900 304.280 ;
        RECT 1333.740 304.000 1337.960 304.280 ;
        RECT 1338.800 304.000 1342.560 304.280 ;
        RECT 1343.400 304.000 1347.620 304.280 ;
        RECT 1348.460 304.000 1352.680 304.280 ;
        RECT 1353.520 304.000 1357.280 304.280 ;
        RECT 1358.120 304.000 1362.340 304.280 ;
        RECT 1363.180 304.000 1367.400 304.280 ;
        RECT 1368.240 304.000 1372.000 304.280 ;
        RECT 1372.840 304.000 1377.060 304.280 ;
        RECT 1377.900 304.000 1381.660 304.280 ;
        RECT 1382.500 304.000 1386.720 304.280 ;
        RECT 1387.560 304.000 1391.780 304.280 ;
        RECT 1392.620 304.000 1396.380 304.280 ;
        RECT 1397.220 304.000 1401.440 304.280 ;
        RECT 1402.280 304.000 1406.500 304.280 ;
        RECT 1407.340 304.000 1411.100 304.280 ;
        RECT 1411.940 304.000 1416.160 304.280 ;
        RECT 1417.000 304.000 1421.220 304.280 ;
        RECT 1422.060 304.000 1425.820 304.280 ;
        RECT 1426.660 304.000 1430.880 304.280 ;
        RECT 1431.720 304.000 1435.940 304.280 ;
        RECT 1436.780 304.000 1440.540 304.280 ;
        RECT 1441.380 304.000 1445.600 304.280 ;
        RECT 1446.440 304.000 1450.660 304.280 ;
        RECT 1451.500 304.000 1455.260 304.280 ;
        RECT 1456.100 304.000 1460.320 304.280 ;
        RECT 1461.160 304.000 1464.920 304.280 ;
        RECT 1465.760 304.000 1469.980 304.280 ;
        RECT 1470.820 304.000 1475.040 304.280 ;
        RECT 1475.880 304.000 1479.640 304.280 ;
        RECT 1480.480 304.000 1484.700 304.280 ;
        RECT 1485.540 304.000 1489.760 304.280 ;
        RECT 1490.600 304.000 1494.360 304.280 ;
        RECT 1495.200 304.000 1499.420 304.280 ;
        RECT 1500.260 304.000 1504.480 304.280 ;
        RECT 1505.320 304.000 1509.080 304.280 ;
        RECT 1509.920 304.000 1514.140 304.280 ;
        RECT 1514.980 304.000 1519.200 304.280 ;
        RECT 1520.040 304.000 1523.800 304.280 ;
        RECT 1524.640 304.000 1528.860 304.280 ;
        RECT 1529.700 304.000 1533.920 304.280 ;
        RECT 1534.760 304.000 1538.520 304.280 ;
        RECT 1539.360 304.000 1543.580 304.280 ;
        RECT 1544.420 304.000 1548.180 304.280 ;
        RECT 1549.020 304.000 1553.240 304.280 ;
        RECT 1554.080 304.000 1558.300 304.280 ;
        RECT 1559.140 304.000 1562.900 304.280 ;
        RECT 1563.740 304.000 1567.960 304.280 ;
        RECT 1568.800 304.000 1573.020 304.280 ;
        RECT 1573.860 304.000 1577.620 304.280 ;
        RECT 1578.460 304.000 1582.680 304.280 ;
        RECT 1583.520 304.000 1587.740 304.280 ;
        RECT 1588.580 304.000 1592.340 304.280 ;
        RECT 1593.180 304.000 1597.400 304.280 ;
        RECT 1598.240 304.000 1602.460 304.280 ;
        RECT 1603.300 304.000 1607.060 304.280 ;
        RECT 1607.900 304.000 1612.120 304.280 ;
        RECT 1612.960 304.000 1617.180 304.280 ;
        RECT 1618.020 304.000 1621.780 304.280 ;
        RECT 1622.620 304.000 1626.840 304.280 ;
        RECT 1627.680 304.000 1631.440 304.280 ;
        RECT 1632.280 304.000 1636.500 304.280 ;
        RECT 1637.340 304.000 1641.560 304.280 ;
        RECT 1642.400 304.000 1646.160 304.280 ;
        RECT 1647.000 304.000 1651.220 304.280 ;
        RECT 1652.060 304.000 1656.280 304.280 ;
        RECT 1657.120 304.000 1660.880 304.280 ;
        RECT 1661.720 304.000 1665.940 304.280 ;
        RECT 1666.780 304.000 1671.000 304.280 ;
        RECT 1671.840 304.000 1675.600 304.280 ;
        RECT 1676.440 304.000 1680.660 304.280 ;
        RECT 1681.500 304.000 1685.720 304.280 ;
        RECT 1686.560 304.000 1690.320 304.280 ;
        RECT 1691.160 304.000 1695.380 304.280 ;
        RECT 1696.220 304.000 1700.440 304.280 ;
        RECT 1701.280 304.000 1705.040 304.280 ;
        RECT 1705.880 304.000 1710.100 304.280 ;
        RECT 1710.940 304.000 1714.700 304.280 ;
        RECT 1715.540 304.000 1719.760 304.280 ;
        RECT 1720.600 304.000 1724.820 304.280 ;
        RECT 1725.660 304.000 1729.420 304.280 ;
        RECT 1730.260 304.000 1734.480 304.280 ;
        RECT 1735.320 304.000 1739.540 304.280 ;
        RECT 1740.380 304.000 1744.140 304.280 ;
        RECT 1744.980 304.000 1749.200 304.280 ;
        RECT 1750.040 304.000 1754.260 304.280 ;
        RECT 1755.100 304.000 1758.860 304.280 ;
        RECT 1759.700 304.000 1763.920 304.280 ;
        RECT 1764.760 304.000 1768.980 304.280 ;
        RECT 1769.820 304.000 1773.580 304.280 ;
        RECT 1774.420 304.000 1778.640 304.280 ;
        RECT 1779.480 304.000 1783.700 304.280 ;
        RECT 1784.540 304.000 1788.300 304.280 ;
        RECT 1789.140 304.000 1793.360 304.280 ;
        RECT 1794.200 304.000 1797.960 304.280 ;
        RECT 1798.800 304.000 1803.020 304.280 ;
        RECT 1803.860 304.000 1808.080 304.280 ;
        RECT 1808.920 304.000 1812.680 304.280 ;
        RECT 1813.520 304.000 1817.740 304.280 ;
        RECT 1818.580 304.000 1822.800 304.280 ;
        RECT 1823.640 304.000 1827.400 304.280 ;
        RECT 1828.240 304.000 1832.460 304.280 ;
        RECT 1833.300 304.000 1837.520 304.280 ;
        RECT 1838.360 304.000 1842.120 304.280 ;
        RECT 1842.960 304.000 1847.180 304.280 ;
        RECT 1848.020 304.000 1852.240 304.280 ;
        RECT 1853.080 304.000 1856.840 304.280 ;
        RECT 1857.680 304.000 1861.900 304.280 ;
        RECT 1862.740 304.000 1866.960 304.280 ;
        RECT 1867.800 304.000 1871.560 304.280 ;
        RECT 1872.400 304.000 1876.620 304.280 ;
        RECT 1877.460 304.000 1881.220 304.280 ;
        RECT 1882.060 304.000 1886.280 304.280 ;
        RECT 1887.120 304.000 1891.340 304.280 ;
        RECT 1892.180 304.000 1895.940 304.280 ;
        RECT 1896.780 304.000 1901.000 304.280 ;
        RECT 1901.840 304.000 1906.060 304.280 ;
        RECT 1906.900 304.000 1910.660 304.280 ;
        RECT 1911.500 304.000 1915.720 304.280 ;
        RECT 1916.560 304.000 1920.780 304.280 ;
        RECT 1921.620 304.000 1925.380 304.280 ;
        RECT 1926.220 304.000 1930.440 304.280 ;
        RECT 1931.280 304.000 1935.500 304.280 ;
        RECT 1936.340 304.000 1940.100 304.280 ;
        RECT 1940.940 304.000 1945.160 304.280 ;
        RECT 1946.000 304.000 1950.220 304.280 ;
        RECT 1951.060 304.000 1954.820 304.280 ;
        RECT 1955.660 304.000 1959.880 304.280 ;
        RECT 1960.720 304.000 1964.480 304.280 ;
        RECT 1965.320 304.000 1969.540 304.280 ;
        RECT 1970.380 304.000 1974.600 304.280 ;
        RECT 1975.440 304.000 1979.200 304.280 ;
        RECT 1980.040 304.000 1984.260 304.280 ;
        RECT 1985.100 304.000 1989.320 304.280 ;
        RECT 1990.160 304.000 1993.920 304.280 ;
        RECT 1994.760 304.000 1998.980 304.280 ;
        RECT 1999.820 304.000 2004.040 304.280 ;
        RECT 2004.880 304.000 2008.640 304.280 ;
        RECT 2009.480 304.000 2013.700 304.280 ;
        RECT 2014.540 304.000 2018.760 304.280 ;
        RECT 2019.600 304.000 2023.360 304.280 ;
        RECT 2024.200 304.000 2028.420 304.280 ;
        RECT 2029.260 304.000 2033.480 304.280 ;
        RECT 2034.320 304.000 2038.080 304.280 ;
        RECT 2038.920 304.000 2043.140 304.280 ;
        RECT 2043.980 304.000 2047.740 304.280 ;
        RECT 2048.580 304.000 2052.800 304.280 ;
        RECT 2053.640 304.000 2057.860 304.280 ;
        RECT 2058.700 304.000 2062.460 304.280 ;
        RECT 2063.300 304.000 2067.520 304.280 ;
        RECT 2068.360 304.000 2072.580 304.280 ;
        RECT 2073.420 304.000 2077.180 304.280 ;
        RECT 2078.020 304.000 2082.240 304.280 ;
        RECT 2083.080 304.000 2087.300 304.280 ;
        RECT 2088.140 304.000 2091.900 304.280 ;
        RECT 2092.740 304.000 2096.960 304.280 ;
        RECT 2097.800 304.000 2102.020 304.280 ;
        RECT 2102.860 304.000 2106.620 304.280 ;
        RECT 2107.460 304.000 2111.680 304.280 ;
        RECT 2112.520 304.000 2116.740 304.280 ;
        RECT 2117.580 304.000 2121.340 304.280 ;
        RECT 2122.180 304.000 2126.400 304.280 ;
        RECT 2127.240 304.000 2131.000 304.280 ;
        RECT 2131.840 304.000 2136.060 304.280 ;
        RECT 2136.900 304.000 2141.120 304.280 ;
        RECT 2141.960 304.000 2145.720 304.280 ;
        RECT 2146.560 304.000 2150.780 304.280 ;
        RECT 2151.620 304.000 2155.840 304.280 ;
        RECT 2156.680 304.000 2160.440 304.280 ;
        RECT 2161.280 304.000 2165.500 304.280 ;
        RECT 2166.340 304.000 2170.560 304.280 ;
        RECT 2171.400 304.000 2175.160 304.280 ;
        RECT 2176.000 304.000 2180.220 304.280 ;
        RECT 2181.060 304.000 2185.280 304.280 ;
        RECT 2186.120 304.000 2189.880 304.280 ;
        RECT 2190.720 304.000 2194.940 304.280 ;
        RECT 2195.780 304.000 2200.000 304.280 ;
        RECT 2200.840 304.000 2204.600 304.280 ;
        RECT 2205.440 304.000 2209.660 304.280 ;
        RECT 2210.500 304.000 2214.260 304.280 ;
        RECT 2215.100 304.000 2219.320 304.280 ;
        RECT 2220.160 304.000 2224.380 304.280 ;
        RECT 2225.220 304.000 2228.980 304.280 ;
        RECT 2229.820 304.000 2234.040 304.280 ;
        RECT 2234.880 304.000 2239.100 304.280 ;
        RECT 2239.940 304.000 2243.700 304.280 ;
        RECT 2244.540 304.000 2248.760 304.280 ;
        RECT 2249.600 304.000 2253.820 304.280 ;
        RECT 2254.660 304.000 2258.420 304.280 ;
        RECT 2259.260 304.000 2263.480 304.280 ;
        RECT 2264.320 304.000 2268.540 304.280 ;
        RECT 2269.380 304.000 2273.140 304.280 ;
        RECT 2273.980 304.000 2278.200 304.280 ;
        RECT 2279.040 304.000 2283.260 304.280 ;
        RECT 2284.100 304.000 2287.860 304.280 ;
        RECT 2288.700 304.000 2292.920 304.280 ;
        RECT 2293.760 304.000 2297.520 304.280 ;
        RECT 2298.360 304.000 2302.580 304.280 ;
        RECT 2303.420 304.000 2307.640 304.280 ;
        RECT 2308.480 304.000 2312.240 304.280 ;
        RECT 2313.080 304.000 2317.300 304.280 ;
        RECT 2318.140 304.000 2322.360 304.280 ;
        RECT 2323.200 304.000 2326.960 304.280 ;
        RECT 2327.800 304.000 2332.020 304.280 ;
        RECT 2332.860 304.000 2337.080 304.280 ;
        RECT 2337.920 304.000 2341.680 304.280 ;
        RECT 2342.520 304.000 2346.740 304.280 ;
        RECT 2347.580 304.000 2351.800 304.280 ;
        RECT 2352.640 304.000 2356.400 304.280 ;
        RECT 2357.240 304.000 2361.460 304.280 ;
        RECT 2362.300 304.000 2366.520 304.280 ;
        RECT 2367.360 304.000 2371.120 304.280 ;
        RECT 2371.960 304.000 2376.180 304.280 ;
        RECT 2377.020 304.000 2380.780 304.280 ;
        RECT 2381.620 304.000 2385.840 304.280 ;
        RECT 2386.680 304.000 2390.900 304.280 ;
        RECT 2391.740 304.000 2395.500 304.280 ;
        RECT 2396.340 304.000 2400.560 304.280 ;
        RECT 2401.400 304.000 2405.620 304.280 ;
        RECT 2406.460 304.000 2410.220 304.280 ;
        RECT 2411.060 304.000 2415.280 304.280 ;
        RECT 2416.120 304.000 2420.340 304.280 ;
        RECT 2421.180 304.000 2424.940 304.280 ;
        RECT 2425.780 304.000 2430.000 304.280 ;
        RECT 2430.840 304.000 2435.060 304.280 ;
        RECT 2435.900 304.000 2439.660 304.280 ;
        RECT 2440.500 304.000 2444.720 304.280 ;
        RECT 2445.560 304.000 2449.780 304.280 ;
        RECT 2450.620 304.000 2454.380 304.280 ;
        RECT 2455.220 304.000 2459.440 304.280 ;
        RECT 2460.280 304.000 2464.040 304.280 ;
        RECT 2464.880 304.000 2469.100 304.280 ;
        RECT 2469.940 304.000 2474.160 304.280 ;
        RECT 2475.000 304.000 2478.760 304.280 ;
        RECT 2479.600 304.000 2483.820 304.280 ;
        RECT 2484.660 304.000 2488.880 304.280 ;
        RECT 2489.720 304.000 2493.480 304.280 ;
        RECT 2494.320 304.000 2498.540 304.280 ;
        RECT 2499.380 304.000 2503.600 304.280 ;
        RECT 2504.440 304.000 2508.200 304.280 ;
        RECT 2509.040 304.000 2513.260 304.280 ;
        RECT 2514.100 304.000 2518.320 304.280 ;
        RECT 2519.160 304.000 2522.920 304.280 ;
        RECT 2523.760 304.000 2527.980 304.280 ;
        RECT 2528.820 304.000 2533.040 304.280 ;
        RECT 2533.880 304.000 2537.640 304.280 ;
        RECT 2538.480 304.000 2542.700 304.280 ;
        RECT 2543.540 304.000 2547.300 304.280 ;
        RECT 2548.140 304.000 2552.360 304.280 ;
        RECT 2553.200 304.000 2557.420 304.280 ;
        RECT 2558.260 304.000 2562.020 304.280 ;
        RECT 2562.860 304.000 2567.080 304.280 ;
        RECT 2567.920 304.000 2572.140 304.280 ;
        RECT 2572.980 304.000 2576.740 304.280 ;
        RECT 2577.580 304.000 2581.800 304.280 ;
        RECT 2582.640 304.000 2586.860 304.280 ;
        RECT 2587.700 304.000 2591.460 304.280 ;
        RECT 2592.300 304.000 2596.520 304.280 ;
        RECT 2597.360 304.000 2601.580 304.280 ;
        RECT 2602.420 304.000 2606.180 304.280 ;
        RECT 2607.020 304.000 2611.240 304.280 ;
        RECT 2612.080 304.000 2616.300 304.280 ;
        RECT 2617.140 304.000 2620.900 304.280 ;
        RECT 2621.740 304.000 2625.960 304.280 ;
        RECT 2626.800 304.000 2630.560 304.280 ;
        RECT 2631.400 304.000 2635.620 304.280 ;
        RECT 2636.460 304.000 2640.680 304.280 ;
        RECT 2641.520 304.000 2645.280 304.280 ;
        RECT 2646.120 304.000 2650.340 304.280 ;
        RECT 2651.180 304.000 2655.400 304.280 ;
        RECT 2656.240 304.000 2660.000 304.280 ;
        RECT 2660.840 304.000 2665.060 304.280 ;
        RECT 2665.900 304.000 2670.120 304.280 ;
        RECT 2670.960 304.000 2674.720 304.280 ;
        RECT 2675.560 304.000 2679.780 304.280 ;
        RECT 2680.620 304.000 2684.840 304.280 ;
        RECT 2685.680 304.000 2689.440 304.280 ;
      LAYER met3 ;
        RECT 308.735 304.255 2686.805 3287.745 ;
      LAYER met4 ;
        RECT 318.670 310.640 320.270 3286.800 ;
      LAYER met4 ;
        RECT 320.925 310.640 328.020 3287.745 ;
        RECT 331.020 310.640 364.020 3287.745 ;
        RECT 367.020 310.640 382.020 3287.745 ;
        RECT 385.020 3287.200 400.020 3287.745 ;
        RECT 385.020 310.640 395.070 3287.200 ;
      LAYER met4 ;
        RECT 395.470 310.640 397.070 3286.800 ;
      LAYER met4 ;
        RECT 397.470 310.640 400.020 3287.200 ;
        RECT 403.020 310.640 418.020 3287.745 ;
        RECT 421.020 310.640 454.020 3287.745 ;
        RECT 457.020 310.640 472.020 3287.745 ;
        RECT 475.020 310.640 490.020 3287.745 ;
        RECT 493.020 310.640 508.020 3287.745 ;
        RECT 511.020 310.640 544.020 3287.745 ;
        RECT 547.020 310.640 562.020 3287.745 ;
        RECT 565.020 310.640 580.020 3287.745 ;
        RECT 583.020 310.640 598.020 3287.745 ;
        RECT 601.020 310.640 634.020 3287.745 ;
        RECT 637.020 310.640 652.020 3287.745 ;
        RECT 655.020 310.640 670.020 3287.745 ;
        RECT 673.020 310.640 688.020 3287.745 ;
        RECT 691.020 310.640 724.020 3287.745 ;
        RECT 727.020 310.640 742.020 3287.745 ;
        RECT 745.020 310.640 760.020 3287.745 ;
        RECT 763.020 310.640 778.020 3287.745 ;
        RECT 781.020 310.640 814.020 3287.745 ;
        RECT 817.020 310.640 832.020 3287.745 ;
        RECT 835.020 310.640 850.020 3287.745 ;
        RECT 853.020 310.640 868.020 3287.745 ;
        RECT 871.020 310.640 904.020 3287.745 ;
        RECT 907.020 310.640 922.020 3287.745 ;
        RECT 925.020 310.640 940.020 3287.745 ;
        RECT 943.020 310.640 958.020 3287.745 ;
        RECT 961.020 310.640 994.020 3287.745 ;
        RECT 997.020 310.640 1012.020 3287.745 ;
        RECT 1015.020 310.640 1030.020 3287.745 ;
        RECT 1033.020 310.640 1048.020 3287.745 ;
        RECT 1051.020 310.640 1084.020 3287.745 ;
        RECT 1087.020 310.640 1102.020 3287.745 ;
        RECT 1105.020 310.640 1120.020 3287.745 ;
        RECT 1123.020 310.640 1138.020 3287.745 ;
        RECT 1141.020 310.640 1174.020 3287.745 ;
        RECT 1177.020 310.640 1192.020 3287.745 ;
        RECT 1195.020 310.640 1210.020 3287.745 ;
        RECT 1213.020 310.640 1228.020 3287.745 ;
        RECT 1231.020 310.640 1264.020 3287.745 ;
        RECT 1267.020 310.640 1282.020 3287.745 ;
        RECT 1285.020 310.640 1300.020 3287.745 ;
        RECT 1303.020 310.640 1318.020 3287.745 ;
        RECT 1321.020 310.640 1354.020 3287.745 ;
        RECT 1357.020 310.640 1372.020 3287.745 ;
        RECT 1375.020 310.640 1390.020 3287.745 ;
        RECT 1393.020 310.640 1408.020 3287.745 ;
        RECT 1411.020 310.640 1444.020 3287.745 ;
        RECT 1447.020 310.640 1462.020 3287.745 ;
        RECT 1465.020 310.640 1480.020 3287.745 ;
        RECT 1483.020 310.640 1498.020 3287.745 ;
        RECT 1501.020 310.640 1534.020 3287.745 ;
        RECT 1537.020 310.640 1552.020 3287.745 ;
        RECT 1555.020 310.640 1570.020 3287.745 ;
        RECT 1573.020 310.640 1588.020 3287.745 ;
        RECT 1591.020 310.640 1624.020 3287.745 ;
        RECT 1627.020 310.640 1642.020 3287.745 ;
        RECT 1645.020 310.640 1660.020 3287.745 ;
        RECT 1663.020 310.640 1678.020 3287.745 ;
        RECT 1681.020 310.640 1714.020 3287.745 ;
        RECT 1717.020 310.640 1732.020 3287.745 ;
        RECT 1735.020 310.640 1750.020 3287.745 ;
        RECT 1753.020 310.640 1768.020 3287.745 ;
        RECT 1771.020 310.640 1804.020 3287.745 ;
        RECT 1807.020 310.640 1822.020 3287.745 ;
        RECT 1825.020 310.640 1840.020 3287.745 ;
        RECT 1843.020 310.640 1858.020 3287.745 ;
        RECT 1861.020 310.640 1894.020 3287.745 ;
        RECT 1897.020 310.640 1912.020 3287.745 ;
        RECT 1915.020 310.640 1930.020 3287.745 ;
        RECT 1933.020 310.640 1948.020 3287.745 ;
        RECT 1951.020 310.640 1984.020 3287.745 ;
        RECT 1987.020 310.640 2002.020 3287.745 ;
        RECT 2005.020 310.640 2020.020 3287.745 ;
        RECT 2023.020 310.640 2038.020 3287.745 ;
        RECT 2041.020 310.640 2074.020 3287.745 ;
        RECT 2077.020 310.640 2092.020 3287.745 ;
        RECT 2095.020 310.640 2110.020 3287.745 ;
        RECT 2113.020 310.640 2128.020 3287.745 ;
        RECT 2131.020 310.640 2164.020 3287.745 ;
        RECT 2167.020 310.640 2182.020 3287.745 ;
        RECT 2185.020 310.640 2200.020 3287.745 ;
        RECT 2203.020 310.640 2218.020 3287.745 ;
        RECT 2221.020 310.640 2254.020 3287.745 ;
        RECT 2257.020 310.640 2272.020 3287.745 ;
        RECT 2275.020 310.640 2290.020 3287.745 ;
        RECT 2293.020 310.640 2308.020 3287.745 ;
        RECT 2311.020 310.640 2344.020 3287.745 ;
        RECT 2347.020 310.640 2362.020 3287.745 ;
        RECT 2365.020 310.640 2380.020 3287.745 ;
        RECT 2383.020 310.640 2398.020 3287.745 ;
        RECT 2401.020 310.640 2434.020 3287.745 ;
        RECT 2437.020 310.640 2452.020 3287.745 ;
        RECT 2455.020 310.640 2470.020 3287.745 ;
        RECT 2473.020 310.640 2488.020 3287.745 ;
        RECT 2491.020 310.640 2524.020 3287.745 ;
        RECT 2527.020 310.640 2542.020 3287.745 ;
        RECT 2545.020 310.640 2560.020 3287.745 ;
        RECT 2563.020 310.640 2578.020 3287.745 ;
        RECT 2581.020 310.640 2614.020 3287.745 ;
        RECT 2617.020 310.640 2632.020 3287.745 ;
        RECT 2635.020 310.640 2650.020 3287.745 ;
        RECT 2653.020 310.640 2668.020 3287.745 ;
        RECT 2671.020 310.640 2676.455 3287.745 ;
  END
END user_project_wrapper
END LIBRARY

